//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G58), .A2(G232), .ZN(new_n205));
  INV_X1    g0005(.A(G87), .ZN(new_n206));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g0008(.A1(G107), .A2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n208), .B(new_n209), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n217), .B1(new_n216), .B2(new_n215), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(G50), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT64), .B(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n221), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT0), .Z(new_n231));
  NOR4_X1   g0031(.A1(new_n223), .A2(new_n224), .A3(new_n228), .A4(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT67), .B(G264), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G13), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n211), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n227), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G50), .ZN(new_n259));
  INV_X1    g0059(.A(G20), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n260), .B1(new_n201), .B2(new_n211), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n226), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT72), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT72), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n226), .A2(new_n268), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT8), .B(G58), .Z(new_n271));
  AOI211_X1 g0071(.A(new_n261), .B(new_n265), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n256), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n254), .B(new_n259), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT70), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT70), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G223), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G222), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  OAI211_X1 g0090(.A(G1), .B(G13), .C1(new_n277), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n289), .B(new_n292), .C1(G77), .C2(new_n285), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT69), .ZN(new_n294));
  OR2_X1    g0094(.A1(KEYINPUT68), .A2(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT68), .A2(G45), .ZN(new_n296));
  AOI21_X1  g0096(.A(G41), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n297), .B2(G1), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT68), .A2(G45), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT68), .A2(G45), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(KEYINPUT69), .B(new_n257), .C1(new_n303), .C2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n298), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n291), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G226), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n293), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n305), .A4(new_n309), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(G200), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n313), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n275), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT76), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n317), .B(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n253), .A2(new_n271), .ZN(new_n322));
  INV_X1    g0122(.A(new_n258), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n271), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n281), .A2(new_n260), .A3(new_n284), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT81), .B(KEYINPUT7), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(KEYINPUT64), .A2(G20), .ZN(new_n330));
  NOR2_X1   g0130(.A1(KEYINPUT64), .A2(G20), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(KEYINPUT80), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT80), .A2(G33), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n279), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n332), .B1(new_n335), .B2(new_n283), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT7), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G68), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n262), .A2(G159), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT82), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G58), .ZN(new_n343));
  INV_X1    g0143(.A(G68), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n345), .B2(new_n201), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT16), .B1(new_n339), .B2(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n333), .A2(new_n334), .A3(new_n279), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n226), .B1(new_n349), .B2(new_n278), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  OR2_X1    g0151(.A1(KEYINPUT80), .A2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(KEYINPUT80), .A2(G33), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(KEYINPUT3), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n282), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n327), .A2(new_n260), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n350), .A2(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(KEYINPUT16), .B(new_n347), .C1(new_n357), .C2(new_n344), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n256), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n325), .B1(new_n348), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n212), .A2(G1698), .ZN(new_n361));
  OR2_X1    g0161(.A1(G223), .A2(G1698), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n354), .A2(new_n282), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n292), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n308), .A2(G232), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n305), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G169), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n366), .A2(G179), .A3(new_n305), .A4(new_n367), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n342), .A2(new_n346), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n332), .B1(new_n354), .B2(new_n282), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n333), .A2(new_n334), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n278), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n327), .A2(new_n260), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n375), .A2(KEYINPUT7), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n374), .B1(new_n379), .B2(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n273), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n344), .B1(new_n329), .B2(new_n337), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n374), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n324), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n369), .A2(new_n370), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n373), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n372), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n368), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n366), .A2(new_n391), .A3(new_n305), .A4(new_n367), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n390), .A2(KEYINPUT83), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT83), .B1(new_n390), .B2(new_n392), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n385), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n385), .B(KEYINPUT17), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n388), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n274), .B1(new_n315), .B2(G169), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n401), .A2(KEYINPUT73), .ZN(new_n402));
  INV_X1    g0202(.A(G179), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n315), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(KEYINPUT73), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT75), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT70), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT70), .B1(new_n282), .B2(new_n283), .ZN(new_n409));
  OAI211_X1 g0209(.A(G232), .B(new_n287), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT74), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n285), .A2(new_n412), .A3(G232), .A4(new_n287), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n408), .A2(new_n409), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G107), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n411), .A2(new_n413), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n292), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n308), .A2(G244), .ZN(new_n419));
  AND4_X1   g0219(.A1(new_n407), .A2(new_n418), .A3(new_n305), .A4(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n305), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n417), .B2(new_n292), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n407), .B1(new_n422), .B2(new_n419), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n403), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n418), .A2(new_n305), .A3(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT75), .ZN(new_n426));
  INV_X1    g0226(.A(G169), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n422), .A2(new_n407), .A3(new_n419), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n271), .A2(new_n262), .ZN(new_n430));
  XOR2_X1   g0230(.A(KEYINPUT15), .B(G87), .Z(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n430), .B1(new_n213), .B2(new_n226), .C1(new_n432), .C2(new_n266), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n256), .B1(new_n213), .B2(new_n253), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n213), .B2(new_n323), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n424), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n321), .A2(new_n400), .A3(new_n406), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n212), .A2(new_n287), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n439), .B1(G232), .B2(new_n287), .C1(new_n408), .C2(new_n409), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n292), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT77), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n307), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n291), .A2(KEYINPUT77), .A3(new_n306), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(G238), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n305), .A2(new_n447), .A3(KEYINPUT78), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT78), .B1(new_n305), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT13), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT13), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G169), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT14), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n451), .A2(G179), .A3(new_n453), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT14), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n458), .A3(G169), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT79), .B1(new_n253), .B2(new_n344), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT12), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT11), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n263), .A2(new_n211), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n260), .A2(G68), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(new_n270), .C2(G77), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(new_n273), .ZN(new_n467));
  INV_X1    g0267(.A(new_n465), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n267), .A2(new_n269), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n213), .ZN(new_n470));
  OAI211_X1 g0270(.A(KEYINPUT11), .B(new_n256), .C1(new_n470), .C2(new_n464), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n258), .A2(G68), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n462), .A2(new_n467), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n460), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n454), .B2(new_n391), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n389), .B1(new_n451), .B2(new_n453), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(G190), .B1(new_n420), .B2(new_n423), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n426), .A2(G200), .A3(new_n428), .ZN(new_n480));
  INV_X1    g0280(.A(new_n435), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n438), .A2(new_n484), .A3(KEYINPUT84), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT84), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n437), .B2(new_n483), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n251), .A2(G20), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g0290(.A(new_n490), .B(KEYINPUT25), .Z(new_n491));
  NAND2_X1  g0291(.A1(new_n257), .A2(G33), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n273), .A2(new_n252), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(G87), .B1(new_n408), .B2(new_n409), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT23), .B1(new_n260), .B2(G107), .ZN(new_n498));
  XOR2_X1   g0298(.A(new_n498), .B(KEYINPUT90), .Z(new_n499));
  NAND4_X1  g0299(.A1(new_n377), .A2(KEYINPUT22), .A3(G87), .A4(new_n226), .ZN(new_n500));
  INV_X1    g0300(.A(G116), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n376), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n502), .A2(new_n260), .B1(new_n332), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT24), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n332), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n352), .A2(new_n353), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G116), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n507), .B1(new_n509), .B2(G20), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n496), .B2(new_n495), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(new_n499), .A4(new_n500), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n494), .B1(new_n514), .B2(new_n256), .ZN(new_n515));
  INV_X1    g0315(.A(G45), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(G1), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G41), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G264), .A3(new_n291), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT91), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n521), .A2(KEYINPUT91), .A3(G264), .A4(new_n291), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G257), .A2(G1698), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n207), .B2(G1698), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n354), .A2(new_n282), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n508), .A2(G294), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n292), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n526), .A2(new_n532), .A3(KEYINPUT92), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT92), .B1(new_n526), .B2(new_n532), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n517), .A2(G274), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n518), .A3(new_n520), .ZN(new_n538));
  AOI21_X1  g0338(.A(G200), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n526), .A2(new_n532), .A3(new_n538), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(G190), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n515), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n538), .ZN(new_n543));
  NOR4_X1   g0343(.A1(new_n533), .A2(new_n534), .A3(new_n403), .A4(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n540), .A2(G169), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n273), .B1(new_n506), .B2(new_n513), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n494), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT87), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n291), .B(G250), .C1(G1), .C2(new_n516), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G238), .A2(G1698), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n214), .B2(G1698), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n502), .B1(new_n377), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n536), .B(new_n549), .C1(new_n552), .C2(new_n291), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n548), .B1(new_n553), .B2(new_n391), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n354), .A3(new_n282), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n291), .B1(new_n555), .B2(new_n509), .ZN(new_n556));
  INV_X1    g0356(.A(new_n549), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n556), .A2(new_n537), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(KEYINPUT87), .A3(G190), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n431), .A2(new_n252), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n493), .A2(new_n206), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n226), .B1(new_n562), .B2(new_n441), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n218), .A2(KEYINPUT85), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT85), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(new_n206), .A3(new_n489), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n354), .A2(new_n226), .A3(G68), .A4(new_n282), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n562), .B1(new_n567), .B2(new_n277), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n560), .B(new_n561), .C1(new_n572), .C2(new_n256), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n553), .A2(G200), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n554), .A2(new_n559), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n560), .B1(new_n572), .B2(new_n256), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n273), .A2(new_n252), .A3(new_n492), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n431), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n558), .A2(new_n403), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(G169), .C2(new_n558), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n542), .A2(new_n547), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n521), .A2(new_n291), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n538), .B1(new_n584), .B2(new_n219), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n354), .A2(new_n587), .A3(new_n282), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G244), .ZN(new_n589));
  NOR2_X1   g0389(.A1(KEYINPUT4), .A2(G244), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n287), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n207), .A2(G1698), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT4), .B1(new_n414), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n592), .A2(new_n595), .B1(G33), .B2(G283), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n586), .B1(new_n596), .B2(new_n291), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n427), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G283), .ZN(new_n599));
  AOI211_X1 g0399(.A(G1698), .B(new_n590), .C1(new_n588), .C2(G244), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n587), .B1(new_n285), .B2(new_n593), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n585), .B1(new_n602), .B2(new_n292), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n403), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n262), .A2(G77), .ZN(new_n605));
  XOR2_X1   g0405(.A(G97), .B(G107), .Z(new_n606));
  NAND2_X1  g0406(.A1(new_n489), .A2(KEYINPUT6), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n606), .A2(KEYINPUT6), .B1(new_n567), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n332), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n326), .A2(new_n328), .B1(new_n336), .B2(KEYINPUT7), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n605), .B(new_n609), .C1(new_n610), .C2(new_n489), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n256), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n252), .A2(new_n218), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n577), .B2(new_n218), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(KEYINPUT86), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(KEYINPUT86), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n598), .A2(new_n604), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n611), .A2(new_n256), .B1(new_n615), .B2(new_n616), .ZN(new_n620));
  OAI211_X1 g0420(.A(G190), .B(new_n586), .C1(new_n596), .C2(new_n291), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n389), .C2(new_n603), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G270), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n538), .B1(new_n584), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n377), .A2(KEYINPUT88), .A3(G257), .A4(new_n287), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n354), .A2(G257), .A3(new_n287), .A4(new_n282), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n377), .A2(G264), .A3(G1698), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n281), .A2(G303), .A3(new_n284), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n626), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n625), .B1(new_n632), .B2(new_n292), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G190), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n226), .B(new_n599), .C1(new_n567), .C2(G33), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n255), .A2(new_n227), .B1(G20), .B2(new_n501), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT20), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT89), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT89), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n251), .A2(G20), .A3(new_n501), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n577), .A2(G116), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n635), .A2(KEYINPUT89), .A3(new_n638), .A4(new_n636), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n634), .B(new_n646), .C1(new_n389), .C2(new_n633), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n633), .A2(G179), .A3(new_n645), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(G169), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n633), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n632), .A2(new_n292), .ZN(new_n652));
  INV_X1    g0452(.A(new_n625), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(KEYINPUT21), .A3(G169), .A4(new_n645), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n647), .A2(new_n648), .A3(new_n651), .A4(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n583), .A2(new_n623), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n488), .A2(new_n657), .ZN(G372));
  AND3_X1   g0458(.A1(new_n655), .A2(new_n651), .A3(new_n648), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n526), .A2(new_n532), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT92), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n526), .A2(new_n532), .A3(KEYINPUT92), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n538), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n389), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(G190), .B2(new_n540), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n659), .A2(new_n547), .B1(new_n666), .B2(new_n515), .ZN(new_n667));
  INV_X1    g0467(.A(new_n623), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT93), .B1(new_n558), .B2(G169), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT93), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n553), .A2(new_n670), .A3(new_n427), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n669), .A2(new_n579), .A3(new_n671), .A4(new_n580), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n573), .B(new_n574), .C1(new_n391), .C2(new_n553), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT94), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT94), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n667), .A2(new_n668), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n619), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n582), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n683), .A3(new_n680), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n679), .A2(new_n682), .A3(new_n672), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n488), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n406), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n424), .A2(new_n435), .A3(new_n429), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n478), .A2(new_n688), .B1(new_n460), .B2(new_n474), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n397), .A2(new_n398), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n388), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n687), .B1(new_n691), .B2(new_n321), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(G369));
  INV_X1    g0493(.A(new_n659), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n226), .A2(G13), .ZN(new_n695));
  OR3_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .A3(G1), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT27), .B1(new_n695), .B2(G1), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G213), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n646), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n694), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n656), .B2(new_n702), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n542), .A2(new_n547), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n515), .B2(new_n701), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n547), .B2(new_n701), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n659), .A2(new_n700), .ZN(new_n711));
  INV_X1    g0511(.A(new_n547), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n707), .A2(new_n711), .B1(new_n712), .B2(new_n701), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(G399));
  NOR2_X1   g0514(.A1(new_n568), .A2(G116), .ZN(new_n715));
  INV_X1    g0515(.A(new_n229), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n225), .B2(new_n718), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT29), .B1(new_n685), .B2(new_n701), .ZN(new_n722));
  INV_X1    g0522(.A(new_n672), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n678), .A2(new_n680), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT26), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n619), .B2(new_n622), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n667), .B(new_n678), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n680), .A2(new_n683), .A3(new_n582), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n725), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n731), .A2(new_n701), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n722), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n662), .A2(new_n663), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n597), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n633), .A2(G179), .A3(new_n558), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT30), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n558), .A2(G179), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n597), .A2(new_n664), .A3(new_n654), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n734), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n736), .A2(new_n738), .A3(KEYINPUT30), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n603), .A2(new_n535), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n737), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(KEYINPUT95), .A3(new_n741), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n743), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(new_n747), .A3(new_n741), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n700), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n542), .A2(new_n547), .A3(new_n582), .ZN(new_n755));
  INV_X1    g0555(.A(new_n656), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n668), .A3(new_n756), .A4(new_n701), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n750), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G330), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n733), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n721), .B1(new_n761), .B2(G1), .ZN(G364));
  OR3_X1    g0562(.A1(new_n695), .A2(KEYINPUT97), .A3(new_n516), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT97), .B1(new_n695), .B2(new_n516), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(G1), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n717), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n706), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n704), .ZN(new_n768));
  INV_X1    g0568(.A(new_n766), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n226), .A2(new_n403), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n389), .A2(G190), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n770), .A2(G190), .A3(new_n389), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT101), .Z(new_n778));
  NOR2_X1   g0578(.A1(new_n389), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G20), .A3(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G303), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n226), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT100), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G329), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n332), .A2(G179), .A3(new_n391), .A4(new_n389), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n332), .A2(new_n391), .A3(new_n779), .ZN(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n786), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G294), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n391), .A2(G179), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n226), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n414), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n226), .A2(new_n403), .A3(new_n391), .A4(new_n389), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n790), .B(new_n794), .C1(G326), .C2(new_n795), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n778), .A2(new_n782), .A3(new_n785), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n788), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G107), .ZN(new_n799));
  INV_X1    g0599(.A(new_n783), .ZN(new_n800));
  INV_X1    g0600(.A(G159), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT32), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n799), .B1(new_n206), .B2(new_n780), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n793), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G97), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n773), .B2(new_n344), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n414), .B(new_n804), .C1(KEYINPUT99), .C2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n795), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n809), .A2(new_n211), .B1(new_n776), .B2(new_n343), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n803), .B2(new_n802), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n808), .B(new_n811), .C1(KEYINPUT99), .C2(new_n807), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT98), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n786), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n786), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n213), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n797), .B1(new_n812), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n227), .B1(G20), .B2(new_n427), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n819), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n377), .A2(new_n716), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n225), .B2(new_n303), .C1(new_n248), .C2(new_n516), .ZN(new_n825));
  INV_X1    g0625(.A(G355), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n285), .A2(new_n229), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(G116), .B2(new_n229), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n818), .A2(new_n819), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n822), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n704), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n768), .B1(new_n769), .B2(new_n831), .ZN(G396));
  NAND2_X1  g0632(.A1(new_n685), .A2(new_n701), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n688), .A2(new_n701), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n481), .A2(new_n701), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n420), .A2(new_n423), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n435), .B1(new_n836), .B2(G200), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(new_n837), .B2(new_n479), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n834), .B1(new_n838), .B2(new_n688), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n436), .A2(new_n700), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n482), .B1(new_n481), .B2(new_n701), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n436), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n685), .A2(new_n701), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(new_n760), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n769), .ZN(new_n847));
  INV_X1    g0647(.A(new_n776), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G143), .B1(G137), .B2(new_n795), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n849), .B1(new_n264), .B2(new_n773), .C1(new_n801), .C2(new_n816), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n377), .B1(new_n211), .B2(new_n780), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n784), .B2(G132), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n798), .A2(G68), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n805), .A2(G58), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n851), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n414), .B1(new_n489), .B2(new_n780), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n806), .B1(new_n206), .B2(new_n788), .C1(new_n773), .C2(new_n789), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(G294), .C2(new_n848), .ZN(new_n859));
  INV_X1    g0659(.A(new_n816), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n860), .A2(G116), .B1(new_n784), .B2(G311), .ZN(new_n861));
  INV_X1    g0661(.A(G303), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n859), .B(new_n861), .C1(new_n862), .C2(new_n809), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n819), .A2(new_n820), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT102), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n864), .A2(new_n819), .B1(new_n213), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n766), .B(new_n868), .C1(new_n843), .C2(new_n821), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n847), .A2(new_n869), .ZN(G384));
  NAND2_X1  g0670(.A1(new_n474), .A2(new_n700), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n458), .B1(new_n454), .B2(G169), .ZN(new_n872));
  AOI211_X1 g0672(.A(KEYINPUT14), .B(new_n427), .C1(new_n451), .C2(new_n453), .ZN(new_n873));
  INV_X1    g0673(.A(new_n457), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n478), .B(new_n871), .C1(new_n875), .C2(new_n473), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n476), .A2(new_n477), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n474), .B(new_n700), .C1(new_n460), .C2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n844), .B2(new_n834), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT104), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n359), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n324), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n698), .ZN(new_n887));
  INV_X1    g0687(.A(new_n698), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n885), .A2(new_n324), .B1(new_n371), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n395), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n360), .B1(new_n371), .B2(new_n888), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n395), .A3(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n399), .A2(new_n887), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n883), .B1(new_n895), .B2(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n399), .A2(new_n887), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n891), .A2(new_n894), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n883), .A3(new_n900), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n880), .A2(new_n881), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n882), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n388), .A2(new_n888), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n892), .A2(new_n395), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n913), .A3(KEYINPUT37), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n912), .A2(new_n894), .A3(new_n914), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n400), .A2(new_n385), .A3(new_n698), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n900), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n895), .A2(KEYINPUT38), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n475), .A2(new_n700), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n908), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n907), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n488), .A2(new_n733), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n692), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n924), .B(new_n926), .Z(new_n927));
  NAND3_X1  g0727(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n757), .A2(new_n754), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT106), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n757), .A2(new_n754), .A3(new_n931), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n839), .B1(new_n876), .B2(new_n878), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(new_n902), .A3(new_n903), .A4(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n876), .A2(new_n878), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n843), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n932), .B2(new_n930), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n917), .B2(new_n919), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n935), .A2(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n488), .A2(new_n933), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(G330), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n927), .B(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n695), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n257), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n501), .B1(new_n608), .B2(KEYINPUT35), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n226), .A2(new_n227), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(KEYINPUT35), .C2(new_n608), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT36), .ZN(new_n951));
  OAI21_X1  g0751(.A(G77), .B1(new_n343), .B2(new_n344), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n225), .A2(new_n952), .B1(G50), .B2(new_n344), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(G1), .A3(new_n250), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n947), .A2(new_n951), .A3(new_n954), .ZN(G367));
  OAI22_X1  g0755(.A1(new_n726), .A2(new_n728), .B1(new_n620), .B2(new_n701), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n680), .A2(new_n700), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT107), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n956), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n712), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n700), .B1(new_n962), .B2(new_n619), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n707), .A2(new_n711), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT42), .Z(new_n966));
  OR3_X1    g0766(.A1(new_n963), .A2(new_n966), .A3(KEYINPUT108), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT108), .B1(new_n963), .B2(new_n966), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n701), .A2(new_n573), .ZN(new_n970));
  MUX2_X1   g0770(.A(new_n678), .B(new_n723), .S(new_n970), .Z(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n973), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n959), .A2(new_n961), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n710), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n977), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n717), .B(KEYINPUT41), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n958), .A2(new_n713), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT45), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n958), .A2(new_n713), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT44), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(new_n710), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n964), .B1(new_n709), .B2(new_n711), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(new_n706), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n761), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n981), .B1(new_n992), .B2(new_n761), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n978), .B(new_n979), .C1(new_n993), .C2(new_n765), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n772), .A2(G294), .B1(G317), .B2(new_n783), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n816), .B2(new_n789), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n776), .A2(new_n862), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n780), .B2(new_n501), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n355), .A3(new_n1000), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n997), .B(new_n1001), .C1(G311), .C2(new_n795), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n489), .B2(new_n793), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n567), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n996), .B(new_n1003), .C1(new_n1004), .C2(new_n798), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n783), .A2(G137), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n772), .A2(G159), .B1(G77), .B2(new_n798), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n816), .B2(new_n211), .ZN(new_n1008));
  INV_X1    g0808(.A(G143), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n809), .A2(new_n1009), .B1(new_n344), .B2(new_n793), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n285), .B1(new_n343), .B2(new_n780), .C1(new_n776), .C2(new_n264), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1005), .B1(new_n1006), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  AOI21_X1  g0814(.A(new_n769), .B1(new_n1014), .B2(new_n819), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n824), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n823), .B1(new_n229), .B2(new_n432), .C1(new_n241), .C2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(new_n830), .C2(new_n971), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n994), .A2(new_n1018), .ZN(G387));
  OAI211_X1 g0819(.A(new_n715), .B(new_n516), .C1(new_n344), .C2(new_n213), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n271), .A2(new_n211), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n824), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT109), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n303), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1024), .B1(new_n237), .B2(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(G107), .B2(new_n229), .C1(new_n715), .C2(new_n827), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n823), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n709), .B2(new_n830), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n783), .A2(G326), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n772), .A2(G311), .B1(G322), .B2(new_n795), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n848), .A2(G317), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n816), .C2(new_n862), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT48), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n789), .B2(new_n793), .C1(new_n791), .C2(new_n780), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n377), .B(new_n1030), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .C1(new_n501), .C2(new_n788), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n271), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n773), .A2(new_n1039), .B1(new_n344), .B2(new_n786), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G150), .B2(new_n783), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n218), .B2(new_n788), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n432), .A2(new_n793), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n776), .B2(new_n211), .C1(new_n801), .C2(new_n809), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1046), .B(new_n377), .C1(new_n213), .C2(new_n780), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1038), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT110), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1029), .B1(new_n1049), .B2(new_n819), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1050), .A2(new_n766), .B1(new_n765), .B2(new_n989), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n717), .B1(new_n761), .B2(new_n989), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n991), .B2(new_n1052), .ZN(G393));
  OR2_X1    g0853(.A1(new_n987), .A2(new_n991), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n717), .A3(new_n992), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n976), .A2(new_n822), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n823), .B1(new_n229), .B2(new_n567), .C1(new_n1016), .C2(new_n245), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n414), .B1(new_n501), .B2(new_n793), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n799), .B1(new_n791), .B2(new_n786), .C1(new_n773), .C2(new_n862), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G283), .C2(new_n781), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n848), .A2(G311), .B1(G317), .B2(new_n795), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT52), .Z(new_n1062));
  OAI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(new_n775), .C2(new_n800), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n377), .B1(new_n793), .B2(new_n213), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n773), .A2(new_n211), .B1(new_n206), .B2(new_n788), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(G68), .C2(new_n781), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n809), .A2(new_n264), .B1(new_n776), .B2(new_n801), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(new_n1039), .C2(new_n816), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n800), .A2(new_n1009), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1063), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n769), .B1(new_n1071), .B2(new_n819), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1056), .A2(new_n1057), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n987), .B2(new_n765), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1055), .A2(new_n1074), .ZN(G390));
  AOI21_X1  g0875(.A(KEYINPUT31), .B1(new_n751), .B2(new_n700), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n657), .B2(new_n701), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n931), .B1(new_n1077), .B2(new_n928), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n932), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n934), .B(G330), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT111), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n933), .A2(KEYINPUT111), .A3(G330), .A4(new_n934), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n909), .B(new_n920), .C1(new_n880), .C2(new_n922), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n922), .B1(new_n917), .B2(new_n919), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n842), .A2(new_n436), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n731), .A2(new_n701), .A3(new_n1087), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1088), .A2(new_n834), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n1089), .B2(new_n879), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1084), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n758), .A2(new_n937), .A3(G330), .A4(new_n843), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1090), .A2(new_n1085), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n488), .A2(G330), .A3(new_n933), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n692), .A3(new_n925), .ZN(new_n1097));
  INV_X1    g0897(.A(G330), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n930), .B2(new_n932), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n937), .B1(new_n1099), .B2(new_n843), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1092), .A2(new_n834), .A3(new_n1088), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT112), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(G330), .B(new_n843), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n879), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1092), .A2(new_n834), .A3(new_n1088), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT112), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n879), .B1(new_n759), .B2(new_n839), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1082), .A2(new_n1083), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n844), .A2(new_n834), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1102), .A2(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1095), .B1(new_n1097), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1090), .A2(new_n1085), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1090), .A2(new_n1085), .A3(new_n1093), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1097), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1112), .A2(new_n717), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n765), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n909), .A2(new_n920), .A3(new_n820), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n848), .A2(G132), .B1(G128), .B2(new_n795), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n772), .A2(G137), .B1(G50), .B2(new_n798), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n780), .A2(new_n264), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  AND4_X1   g0929(.A1(new_n285), .A2(new_n1126), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(KEYINPUT54), .B(G143), .Z(new_n1131));
  AOI22_X1  g0931(.A1(new_n860), .A2(new_n1131), .B1(new_n784), .B2(G125), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n801), .C2(new_n793), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n776), .A2(new_n501), .B1(new_n213), .B2(new_n793), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT113), .Z(new_n1135));
  AOI22_X1  g0935(.A1(new_n860), .A2(new_n1004), .B1(new_n784), .B2(G294), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n854), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n414), .B1(new_n773), .B2(new_n489), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G283), .B2(new_n795), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n206), .B2(new_n780), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1133), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(new_n819), .B1(new_n1039), .B2(new_n867), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1125), .A2(new_n766), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT114), .B1(new_n1124), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT114), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1146), .B(new_n1143), .C1(new_n1095), .C2(new_n1123), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1122), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G378));
  INV_X1    g0950(.A(KEYINPUT57), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n274), .A2(new_n888), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT56), .Z(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT55), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n321), .A2(new_n1155), .A3(new_n406), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1155), .B1(new_n321), .B2(new_n406), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1154), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n1156), .A3(new_n1153), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT115), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n941), .B2(G330), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n934), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n936), .B1(new_n1165), .B2(new_n904), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n917), .A2(new_n919), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1167), .A2(new_n933), .A3(KEYINPUT40), .A4(new_n934), .ZN(new_n1168));
  AND4_X1   g0968(.A1(G330), .A2(new_n1166), .A3(new_n1168), .A4(new_n1163), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n924), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1166), .A2(G330), .A3(new_n1168), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1163), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1166), .A2(new_n1168), .A3(new_n1163), .A4(G330), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n923), .A3(new_n907), .A4(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1097), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1151), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT117), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1170), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1117), .B1(new_n1095), .B2(new_n1111), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n924), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(KEYINPUT117), .A3(new_n1174), .A4(new_n1173), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(KEYINPUT57), .A4(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1178), .A2(new_n1184), .A3(new_n717), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n765), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT116), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1159), .A2(new_n1161), .A3(new_n820), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n867), .A2(new_n211), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n795), .A2(G125), .ZN(new_n1191));
  INV_X1    g0991(.A(G128), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n776), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n772), .A2(G132), .B1(new_n781), .B2(new_n1131), .ZN(new_n1194));
  INV_X1    g0994(.A(G137), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n786), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(G150), .C2(new_n805), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT59), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G41), .B1(new_n783), .B2(G124), .ZN(new_n1199));
  AOI21_X1  g0999(.A(G33), .B1(new_n798), .B2(G159), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n355), .B1(new_n793), .B2(new_n344), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n290), .B1(new_n213), .B2(new_n780), .C1(new_n809), .C2(new_n501), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G107), .C2(new_n848), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n786), .A2(new_n432), .B1(new_n788), .B2(new_n343), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n784), .B2(G283), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(new_n218), .C2(new_n773), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G41), .B1(new_n333), .B2(KEYINPUT3), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1201), .B(new_n1208), .C1(G50), .C2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n769), .B1(new_n1210), .B2(new_n819), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1189), .A2(new_n1190), .A3(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1187), .A2(new_n1188), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1123), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1212), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT116), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1185), .A2(new_n1217), .ZN(G375));
  INV_X1    g1018(.A(KEYINPUT119), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1111), .B2(new_n1123), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1120), .A2(KEYINPUT119), .A3(new_n765), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n414), .B1(new_n218), .B2(new_n780), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1044), .B1(new_n213), .B2(new_n788), .C1(new_n773), .C2(new_n501), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(G283), .C2(new_n848), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n860), .A2(G107), .B1(new_n784), .B2(G303), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n791), .C2(new_n809), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n377), .B1(new_n793), .B2(new_n211), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n776), .A2(new_n1195), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(G132), .C2(new_n795), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n772), .A2(new_n1131), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n781), .A2(G159), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n786), .A2(new_n264), .B1(new_n788), .B2(new_n343), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n784), .B2(G128), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1226), .A2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1235), .A2(new_n819), .B1(new_n344), .B2(new_n867), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n766), .B(new_n1236), .C1(new_n937), .C2(new_n821), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1220), .A2(new_n1221), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1118), .A2(new_n1119), .A3(new_n1097), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT118), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1118), .A2(new_n1119), .A3(KEYINPUT118), .A4(new_n1097), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1097), .B2(new_n1111), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1238), .B1(new_n1244), .B2(new_n981), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT120), .ZN(G381));
  NOR4_X1   g1046(.A1(G381), .A2(G396), .A3(G387), .A4(G393), .ZN(new_n1247));
  INV_X1    g1047(.A(G384), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(G375), .A2(G378), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(G407));
  NAND2_X1  g1051(.A1(new_n1181), .A2(new_n1186), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n718), .B1(new_n1252), .B2(new_n1151), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1253), .A2(new_n1184), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1149), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n699), .A2(G213), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT121), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G407), .B(G213), .C1(new_n1255), .C2(new_n1258), .ZN(G409));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT123), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(KEYINPUT123), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1120), .B2(new_n1117), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1261), .A2(new_n1263), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n717), .B1(new_n1239), .B2(new_n1260), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G384), .B(new_n1238), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT124), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1238), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1262), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1261), .B(new_n1269), .C1(new_n1111), .C2(new_n1097), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1265), .B1(new_n1243), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1248), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1243), .A2(new_n1270), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1265), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT124), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(G384), .A4(new_n1238), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1267), .A2(new_n1272), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1257), .A2(G2897), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1279), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1267), .A2(new_n1272), .A3(new_n1277), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1180), .A2(KEYINPUT122), .A3(new_n1183), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT122), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n765), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1215), .B1(new_n1287), .B2(new_n980), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1149), .A3(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1289), .B(new_n1258), .C1(new_n1149), .C2(new_n1254), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1283), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(KEYINPUT126), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1257), .B1(G375), .B2(G378), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1280), .A2(new_n1282), .B1(new_n1289), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1296), .B2(KEYINPUT61), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT62), .B1(new_n1290), .B2(new_n1278), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1278), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT62), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(new_n1295), .A3(new_n1300), .A4(new_n1289), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1293), .A2(new_n1297), .A3(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(G396), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n994), .A2(new_n1018), .A3(G390), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G390), .B1(new_n994), .B2(new_n1018), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1304), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G387), .A2(new_n1249), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n994), .A2(new_n1018), .A3(G390), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1304), .A2(KEYINPUT125), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1305), .A2(KEYINPUT125), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1307), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1303), .A2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1290), .A2(new_n1278), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1313), .B1(KEYINPUT63), .B2(new_n1315), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1291), .A2(KEYINPUT63), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1316), .B(new_n1292), .C1(new_n1317), .C2(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1314), .A2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(G375), .A2(G378), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1255), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(KEYINPUT127), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1320), .A2(new_n1255), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1325), .A2(new_n1307), .A3(new_n1312), .A4(new_n1311), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1313), .A2(new_n1322), .A3(new_n1324), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1326), .A2(new_n1299), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1299), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


