//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n212), .B1(new_n214), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G87), .B(G97), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  XOR2_X1   g0042(.A(KEYINPUT8), .B(G58), .Z(new_n243));
  NAND2_X1  g0043(.A1(new_n206), .A2(G20), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n245), .A2(new_n249), .B1(new_n246), .B2(new_n243), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT16), .ZN(new_n251));
  INV_X1    g0051(.A(G58), .ZN(new_n252));
  INV_X1    g0052(.A(G68), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(G20), .B1(new_n254), .B2(new_n201), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G159), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(G20), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n253), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT74), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n259), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI211_X1 g0069(.A(KEYINPUT74), .B(new_n253), .C1(new_n262), .C2(new_n266), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n251), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n248), .A2(new_n247), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(new_n258), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(KEYINPUT16), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n250), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n277), .A2(KEYINPUT66), .A3(new_n247), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT66), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n279), .B1(new_n213), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(G223), .A2(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G1698), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n283), .B(new_n285), .C1(new_n263), .C2(new_n264), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G87), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n286), .A2(KEYINPUT75), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT75), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT76), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT76), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n292), .B(new_n282), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  AOI21_X1  g0095(.A(G1), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(G274), .ZN(new_n298));
  INV_X1    g0098(.A(G232), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G190), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n291), .A2(new_n293), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  INV_X1    g0105(.A(new_n282), .ZN(new_n306));
  INV_X1    g0106(.A(new_n289), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n286), .A2(KEYINPUT75), .A3(new_n287), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n305), .B1(new_n309), .B2(new_n302), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n276), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT17), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n276), .A2(new_n311), .A3(KEYINPUT17), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT18), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n302), .A2(G179), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n291), .A2(new_n293), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n309), .B2(new_n302), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n317), .B1(new_n276), .B2(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n276), .A2(new_n322), .A3(new_n317), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(KEYINPUT77), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n276), .A2(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT77), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n317), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n316), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n207), .A2(G33), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n243), .A2(new_n331), .B1(G150), .B2(new_n256), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n203), .A2(G20), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n273), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n244), .A2(G50), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n249), .A2(new_n335), .B1(G50), .B2(new_n246), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT9), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT9), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n334), .B2(new_n336), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  OR2_X1    g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  AOI21_X1  g0144(.A(G1698), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G222), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n261), .A2(G223), .A3(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G77), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n261), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n282), .ZN(new_n350));
  INV_X1    g0150(.A(new_n301), .ZN(new_n351));
  INV_X1    g0151(.A(G274), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n213), .B2(new_n280), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n351), .A2(G226), .B1(new_n296), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(G190), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n350), .A2(new_n354), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G200), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n341), .A2(new_n342), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n357), .A2(new_n340), .A3(new_n355), .A4(new_n338), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT10), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n337), .B1(new_n356), .B2(new_n320), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G179), .B2(new_n356), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G87), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n365), .A2(KEYINPUT15), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(KEYINPUT15), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n331), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT8), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(G58), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n252), .A2(KEYINPUT8), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n256), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G20), .A2(G77), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n272), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n244), .A2(G77), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n249), .A2(new_n376), .B1(G77), .B2(new_n246), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G1698), .ZN(new_n380));
  OAI211_X1 g0180(.A(G232), .B(new_n380), .C1(new_n263), .C2(new_n264), .ZN(new_n381));
  OAI211_X1 g0181(.A(G238), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n343), .A2(G107), .A3(new_n344), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n282), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n297), .A2(G244), .A3(new_n300), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n298), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n379), .B1(G200), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G190), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n389), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n377), .B1(new_n374), .B2(new_n272), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n389), .B2(new_n320), .ZN(new_n394));
  INV_X1    g0194(.A(G179), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n385), .A2(new_n395), .A3(new_n388), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT67), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n387), .B1(new_n282), .B2(new_n384), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT67), .B1(new_n399), .B2(new_n395), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n394), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n364), .A2(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n329), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n256), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n202), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n330), .A2(new_n348), .B1(new_n207), .B2(G68), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n272), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT11), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n246), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT72), .B1(new_n411), .B2(new_n253), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT12), .ZN(new_n413));
  INV_X1    g0213(.A(new_n249), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(G68), .A3(new_n244), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n408), .A2(new_n409), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n410), .A2(new_n413), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(G232), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT68), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n261), .A2(KEYINPUT68), .A3(G232), .A4(G1698), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G97), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n261), .A2(G226), .A3(new_n380), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n282), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n351), .A2(KEYINPUT70), .ZN(new_n427));
  INV_X1    g0227(.A(G238), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT70), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n301), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G274), .B1(new_n277), .B2(new_n247), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT69), .B1(new_n431), .B2(new_n300), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT69), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n353), .A2(new_n433), .A3(new_n296), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n427), .A2(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n425), .A2(new_n426), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n391), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n425), .A2(new_n435), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT13), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n417), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n425), .A2(new_n435), .A3(new_n426), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n425), .A2(new_n435), .A3(KEYINPUT71), .A4(new_n426), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(G200), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n426), .B1(new_n425), .B2(new_n435), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n436), .A2(new_n448), .A3(KEYINPUT71), .ZN(new_n449));
  INV_X1    g0249(.A(new_n444), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT14), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n451), .A2(KEYINPUT73), .A3(new_n452), .A4(G169), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT73), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(G169), .A3(new_n444), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(KEYINPUT14), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n436), .A2(new_n448), .A3(new_n395), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n455), .B2(KEYINPUT14), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n447), .B1(new_n459), .B2(new_n417), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n404), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n206), .A2(G33), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n246), .A2(new_n463), .A3(new_n247), .A4(new_n248), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G116), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n411), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n248), .A2(new_n247), .B1(G20), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n470), .B(new_n207), .C1(G33), .C2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n469), .A2(KEYINPUT20), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT20), .B1(new_n469), .B2(new_n472), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n466), .B(new_n468), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n295), .A2(G1), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT78), .B1(new_n481), .B2(new_n431), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n206), .A2(G45), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n294), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n478), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT78), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n353), .ZN(new_n488));
  INV_X1    g0288(.A(new_n297), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n482), .A2(new_n488), .B1(new_n490), .B2(G270), .ZN(new_n491));
  OAI211_X1 g0291(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n492));
  OAI211_X1 g0292(.A(G257), .B(new_n380), .C1(new_n263), .C2(new_n264), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n343), .A2(G303), .A3(new_n344), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n282), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(G190), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n482), .A2(new_n488), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n481), .A2(G270), .A3(new_n297), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n476), .B(new_n497), .C1(new_n501), .C2(new_n305), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(G169), .A3(new_n475), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT21), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n475), .A2(new_n491), .A3(G179), .A4(new_n496), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n500), .A2(KEYINPUT21), .A3(new_n475), .A4(G169), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n502), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT80), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n507), .A2(new_n506), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT80), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n505), .A4(new_n502), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT81), .B1(new_n514), .B2(G20), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT81), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(new_n207), .A3(G33), .A4(G116), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT82), .B1(new_n207), .B2(G107), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT23), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT82), .B(KEYINPUT23), .C1(new_n207), .C2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n523));
  AND4_X1   g0323(.A1(new_n518), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n261), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n207), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n526), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n518), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n531), .A2(new_n532), .B1(KEYINPUT83), .B2(KEYINPUT24), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n272), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT25), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n246), .B2(G107), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n246), .A2(new_n536), .A3(G107), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(KEYINPUT84), .B(new_n536), .C1(new_n246), .C2(G107), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n540), .A2(new_n541), .B1(G107), .B2(new_n465), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n544));
  OAI211_X1 g0344(.A(G250), .B(new_n380), .C1(new_n263), .C2(new_n264), .ZN(new_n545));
  INV_X1    g0345(.A(G33), .ZN(new_n546));
  INV_X1    g0346(.A(G294), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n282), .B1(new_n490), .B2(G264), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n498), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n320), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n395), .A3(new_n498), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n543), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G238), .B(new_n380), .C1(new_n263), .C2(new_n264), .ZN(new_n554));
  OAI211_X1 g0354(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n514), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n282), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n297), .A2(G250), .A3(new_n483), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n431), .B2(new_n483), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n560), .A3(G190), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n282), .B2(new_n556), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n305), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n366), .A2(new_n367), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n246), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n464), .A2(new_n365), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n261), .A2(new_n207), .A3(G68), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n330), .B2(new_n471), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n207), .B1(new_n422), .B2(new_n570), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G97), .A2(G107), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n365), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT79), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n567), .B(new_n568), .C1(new_n582), .C2(new_n272), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n564), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n567), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n565), .A2(new_n464), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n572), .B1(new_n580), .B2(new_n578), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n585), .B(new_n587), .C1(new_n588), .C2(new_n273), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n557), .A2(new_n560), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n320), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n562), .A2(new_n395), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n549), .A2(new_n391), .A3(new_n498), .ZN(new_n594));
  AOI21_X1  g0394(.A(G200), .B1(new_n549), .B2(new_n498), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n584), .B(new_n593), .C1(new_n543), .C2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n246), .A2(G97), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n465), .B2(G97), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g0400(.A(G97), .B(G107), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n602), .A2(new_n471), .A3(G107), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n262), .A2(new_n266), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G107), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n600), .B1(new_n610), .B2(new_n272), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n482), .A2(new_n488), .B1(new_n490), .B2(G257), .ZN(new_n612));
  OAI211_X1 g0412(.A(G250), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n613));
  OAI211_X1 g0413(.A(G244), .B(new_n380), .C1(new_n263), .C2(new_n264), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT4), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n470), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT4), .B1(new_n345), .B2(G244), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n282), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n611), .B(new_n620), .C1(new_n391), .C2(new_n619), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n320), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n604), .B1(new_n602), .B2(new_n601), .ZN(new_n623));
  OAI22_X1  g0423(.A1(new_n623), .A2(new_n207), .B1(new_n348), .B2(new_n405), .ZN(new_n624));
  INV_X1    g0424(.A(G107), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n262), .B2(new_n266), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n272), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n599), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n612), .A2(new_n618), .A3(new_n395), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n621), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n597), .A2(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n462), .A2(new_n513), .A3(new_n553), .A4(new_n632), .ZN(G372));
  NAND2_X1  g0433(.A1(new_n459), .A2(new_n417), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n401), .A2(KEYINPUT85), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT85), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n394), .B(new_n636), .C1(new_n398), .C2(new_n400), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n446), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n316), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n276), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(KEYINPUT18), .A3(new_n319), .A4(new_n321), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n323), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n361), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n363), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n567), .B(new_n586), .C1(new_n582), .C2(new_n272), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n591), .A2(new_n592), .ZN(new_n648));
  INV_X1    g0448(.A(new_n568), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n585), .B(new_n649), .C1(new_n588), .C2(new_n273), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n647), .A2(new_n648), .B1(new_n650), .B2(new_n563), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n646), .B1(new_n651), .B2(new_n630), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n584), .A4(new_n593), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n648), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n656), .A2(new_n589), .B1(new_n564), .B2(new_n583), .ZN(new_n657));
  INV_X1    g0457(.A(new_n542), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n272), .B2(new_n534), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n594), .B2(new_n595), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n657), .A2(new_n660), .A3(new_n630), .A4(new_n621), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n551), .A2(new_n552), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n655), .B(new_n593), .C1(new_n661), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n462), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n645), .A2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n476), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n509), .B2(new_n512), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n664), .A2(new_n676), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n677), .A2(KEYINPUT86), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT86), .B1(new_n677), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n543), .A2(new_n674), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n663), .B1(new_n682), .B2(new_n660), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n553), .A2(new_n674), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n681), .A2(G330), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n660), .A2(new_n682), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n553), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n664), .A2(new_n675), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n684), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n686), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(KEYINPUT87), .ZN(new_n693));
  INV_X1    g0493(.A(new_n210), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(G41), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n210), .A2(KEYINPUT87), .A3(new_n294), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n575), .A2(new_n365), .A3(new_n467), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n698), .A2(new_n206), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n216), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n698), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n666), .A2(new_n675), .ZN(new_n704));
  XNOR2_X1  g0504(.A(KEYINPUT89), .B(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n666), .B(new_n675), .C1(KEYINPUT89), .C2(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n513), .A2(new_n632), .A3(new_n553), .A4(new_n675), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n548), .A2(new_n282), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n490), .A2(G264), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n557), .A3(new_n711), .A4(new_n560), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n498), .A2(new_n496), .A3(G179), .A4(new_n499), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n619), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT30), .B1(new_n714), .B2(KEYINPUT88), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT88), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  INV_X1    g0517(.A(new_n712), .ZN(new_n718));
  INV_X1    g0518(.A(new_n713), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n716), .B(new_n717), .C1(new_n720), .C2(new_n619), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n501), .A2(G179), .A3(new_n562), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(new_n550), .A3(new_n619), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n715), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n674), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n709), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n708), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n703), .B1(new_n731), .B2(new_n206), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT90), .ZN(G364));
  NAND2_X1  g0533(.A1(new_n681), .A2(G330), .ZN(new_n734));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n206), .B1(new_n736), .B2(G45), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n697), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT91), .Z(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G330), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n679), .A2(new_n741), .A3(new_n680), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n734), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n677), .A2(new_n678), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n739), .B(KEYINPUT92), .Z(new_n749));
  NAND2_X1  g0549(.A1(new_n391), .A2(G20), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT93), .B(G159), .Z(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n758));
  AOI21_X1  g0558(.A(new_n207), .B1(new_n752), .B2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n757), .A2(new_n758), .B1(G97), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n207), .A2(new_n391), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G179), .A3(new_n305), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n761), .B1(new_n252), .B2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n750), .A2(new_n395), .A3(new_n305), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n750), .A2(new_n395), .A3(G200), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G68), .A2(new_n765), .B1(new_n766), .B2(G77), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n762), .A2(new_n395), .A3(G200), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n261), .C1(new_n365), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n762), .A2(G179), .A3(G200), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n757), .A2(new_n758), .B1(new_n202), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n764), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n751), .A2(new_n395), .A3(G200), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT95), .Z(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT96), .Z(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G107), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(G283), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n261), .B1(new_n754), .B2(G329), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n547), .B2(new_n759), .ZN(new_n779));
  INV_X1    g0579(.A(G317), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(KEYINPUT33), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n765), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  INV_X1    g0585(.A(new_n766), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n783), .B1(new_n784), .B2(new_n768), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  INV_X1    g0588(.A(G326), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n763), .A2(new_n788), .B1(new_n770), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n779), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n772), .A2(new_n776), .B1(new_n777), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n247), .B1(G20), .B2(new_n320), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n746), .A2(new_n793), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n241), .A2(G45), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n694), .A2(new_n261), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G45), .C2(new_n216), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n694), .A2(new_n265), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(G355), .B1(new_n467), .B2(new_n694), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n797), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n748), .A2(new_n749), .A3(new_n795), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n743), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n675), .A2(new_n393), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n635), .B2(new_n637), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(new_n392), .B2(new_n401), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n809), .A2(KEYINPUT98), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT98), .ZN(new_n812));
  INV_X1    g0612(.A(new_n637), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n396), .A2(new_n397), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n399), .A2(KEYINPUT67), .A3(new_n395), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n636), .B1(new_n816), .B2(new_n394), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n807), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n402), .A2(new_n808), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n811), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n704), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT98), .B1(new_n809), .B2(new_n810), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n818), .A2(new_n819), .A3(new_n812), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n666), .A2(new_n825), .A3(new_n675), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n730), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT99), .Z(new_n829));
  AOI21_X1  g0629(.A(new_n739), .B1(new_n827), .B2(new_n730), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n261), .B1(new_n768), .B2(new_n202), .C1(new_n832), .C2(new_n753), .ZN(new_n833));
  INV_X1    g0633(.A(new_n775), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n253), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(G58), .C2(new_n760), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n756), .A2(new_n766), .B1(G150), .B2(new_n765), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(G143), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n838), .B2(new_n770), .C1(new_n839), .C2(new_n763), .ZN(new_n840));
  XOR2_X1   g0640(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n841));
  XNOR2_X1  g0641(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n775), .A2(G87), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n754), .A2(G311), .B1(G283), .B2(new_n765), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n467), .B2(new_n786), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n265), .B1(new_n759), .B2(new_n471), .C1(new_n768), .C2(new_n625), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n763), .A2(new_n547), .B1(new_n770), .B2(new_n784), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n794), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n793), .A2(new_n744), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n749), .B(new_n851), .C1(new_n348), .C2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n745), .B2(new_n825), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n831), .A2(new_n854), .ZN(G384));
  OAI21_X1  g0655(.A(G77), .B1(new_n252), .B2(new_n253), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n216), .A2(new_n856), .B1(G50), .B2(new_n253), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(G1), .A3(new_n735), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT100), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n467), .B(new_n214), .C1(new_n606), .C2(KEYINPUT35), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(KEYINPUT35), .B2(new_n606), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT36), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  INV_X1    g0664(.A(new_n672), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n640), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n326), .A2(new_n866), .A3(new_n867), .A4(new_n312), .ZN(new_n868));
  INV_X1    g0668(.A(new_n312), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n251), .B1(new_n267), .B2(new_n258), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n250), .B1(new_n275), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n322), .B2(new_n672), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n871), .A2(new_n672), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n329), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT38), .B(new_n874), .C1(new_n329), .C2(new_n875), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n417), .A2(new_n674), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n634), .A2(new_n446), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n417), .B(new_n674), .C1(new_n459), .C2(new_n447), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n816), .A2(new_n394), .A3(new_n675), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n882), .A2(new_n883), .B1(new_n826), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n643), .A2(new_n672), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT101), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  INV_X1    g0691(.A(new_n879), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n276), .A2(new_n311), .A3(KEYINPUT17), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT17), .B1(new_n276), .B2(new_n311), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT102), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT102), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n314), .A2(new_n896), .A3(new_n315), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n897), .A3(new_n642), .ZN(new_n898));
  INV_X1    g0698(.A(new_n866), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n326), .A2(new_n866), .A3(new_n312), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n868), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n891), .B1(new_n892), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n634), .A2(new_n674), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n886), .A2(KEYINPUT101), .A3(new_n887), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n890), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n706), .A2(new_n404), .A3(new_n707), .A4(new_n460), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n645), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n882), .A2(new_n883), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT31), .B1(new_n724), .B2(new_n674), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n821), .B1(new_n917), .B2(new_n709), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n914), .B(new_n918), .C1(new_n892), .C2(new_n904), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT40), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT40), .B1(new_n878), .B2(new_n879), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n729), .A2(new_n825), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n882), .B2(new_n883), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n461), .B1(new_n709), .B2(new_n917), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n741), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n925), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n913), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n206), .B2(new_n736), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n913), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n864), .B1(new_n930), .B2(new_n931), .ZN(G367));
  OAI21_X1  g0732(.A(new_n796), .B1(new_n210), .B2(new_n565), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n799), .B2(new_n233), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n749), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n650), .A2(new_n674), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n657), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n593), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n774), .A2(G77), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n759), .A2(new_n253), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n265), .B(new_n941), .C1(G50), .C2(new_n766), .ZN(new_n942));
  INV_X1    g0742(.A(new_n770), .ZN(new_n943));
  INV_X1    g0743(.A(new_n763), .ZN(new_n944));
  AOI22_X1  g0744(.A1(G143), .A2(new_n943), .B1(new_n944), .B2(G150), .ZN(new_n945));
  INV_X1    g0745(.A(new_n765), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n946), .A2(new_n755), .B1(new_n838), .B2(new_n753), .ZN(new_n947));
  INV_X1    g0747(.A(new_n768), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(G58), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n940), .A2(new_n942), .A3(new_n945), .A4(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(G283), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n265), .B1(new_n753), .B2(new_n780), .C1(new_n786), .C2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n774), .B2(G97), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n763), .A2(new_n784), .B1(new_n759), .B2(new_n625), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT105), .B(G311), .Z(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n943), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT106), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n948), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n768), .B2(new_n467), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n960), .C1(new_n547), .C2(new_n946), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n953), .B(new_n956), .C1(new_n957), .C2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n957), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n950), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT107), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT47), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n935), .B1(new_n747), .B2(new_n939), .C1(new_n966), .C2(new_n794), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n621), .B(new_n630), .C1(new_n611), .C2(new_n675), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n653), .A2(new_n674), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n686), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n939), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n685), .A2(new_n690), .A3(new_n970), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n976), .A2(KEYINPUT103), .A3(KEYINPUT42), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT103), .B1(new_n976), .B2(KEYINPUT42), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n968), .A2(new_n553), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n674), .B1(new_n980), .B2(new_n630), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(KEYINPUT42), .B2(new_n976), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n975), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n979), .A2(new_n974), .A3(new_n973), .A4(new_n982), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n972), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n972), .A3(new_n987), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n737), .ZN(new_n992));
  INV_X1    g0792(.A(new_n731), .ZN(new_n993));
  NOR2_X1   g0793(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n691), .B2(new_n970), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n683), .A2(new_n689), .B1(new_n553), .B2(new_n674), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n971), .C1(KEYINPUT104), .C2(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n996), .B2(new_n971), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1004), .A2(G330), .A3(new_n681), .A4(new_n685), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n686), .A2(new_n1003), .A3(new_n999), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n685), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n689), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n685), .A2(new_n690), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n681), .A2(G330), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(new_n681), .B2(G330), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n993), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n697), .B(KEYINPUT41), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n992), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n967), .B1(new_n991), .B2(new_n1018), .ZN(G387));
  OAI21_X1  g0819(.A(new_n265), .B1(new_n753), .B2(new_n789), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n765), .A2(new_n955), .B1(new_n766), .B2(G303), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n780), .B2(new_n763), .C1(new_n788), .C2(new_n770), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n768), .A2(new_n547), .B1(new_n759), .B2(new_n951), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT108), .Z(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT49), .Z(new_n1029));
  AOI211_X1 g0829(.A(new_n1020), .B(new_n1029), .C1(G116), .C2(new_n774), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n834), .A2(new_n471), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n948), .A2(G77), .B1(new_n765), .B2(new_n243), .ZN(new_n1032));
  INV_X1    g0832(.A(G150), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n1033), .B2(new_n753), .ZN(new_n1034));
  INV_X1    g0834(.A(G159), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n261), .B1(new_n770), .B2(new_n1035), .C1(new_n786), .C2(new_n253), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n566), .A2(new_n760), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n202), .B2(new_n763), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1031), .A2(new_n1034), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n793), .B1(new_n1030), .B2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n801), .A2(new_n699), .B1(new_n625), .B2(new_n694), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n230), .A2(G45), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT50), .B1(new_n243), .B2(new_n202), .ZN(new_n1044));
  AND3_X1   g0844(.A1(new_n243), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n799), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1041), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n749), .B1(new_n796), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1040), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1008), .B2(new_n746), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1014), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n992), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1014), .A2(new_n731), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n993), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n1055), .A3(new_n698), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT109), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT109), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1053), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(G393));
  NAND3_X1  g0861(.A1(new_n1005), .A2(new_n992), .A3(new_n1006), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n763), .A2(new_n1035), .B1(new_n770), .B2(new_n1033), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n759), .A2(new_n348), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n243), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n261), .B1(new_n786), .B2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(G50), .C2(new_n765), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n839), .A2(new_n753), .B1(new_n768), .B2(new_n253), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT110), .Z(new_n1070));
  NAND4_X1  g0870(.A1(new_n844), .A2(new_n1064), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n265), .B1(new_n759), .B2(new_n467), .C1(new_n768), .C2(new_n951), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n786), .A2(new_n547), .B1(new_n753), .B2(new_n788), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G303), .C2(new_n765), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n763), .A2(new_n785), .B1(new_n770), .B2(new_n780), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n776), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n794), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n238), .A2(new_n799), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n797), .B1(G97), .B2(new_n694), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n749), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n970), .B2(new_n747), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1062), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n698), .B1(new_n1007), .B2(new_n1055), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1007), .A2(new_n1055), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(G390));
  NAND2_X1  g0888(.A1(new_n826), .A2(new_n884), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n883), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n881), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n447), .B(new_n1091), .C1(new_n459), .C2(new_n417), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1089), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n906), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n905), .A3(new_n907), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n906), .B1(new_n914), .B2(new_n1089), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n892), .A2(new_n904), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(G330), .B(new_n918), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1096), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n404), .A2(G330), .A3(new_n460), .A4(new_n729), .ZN(new_n1104));
  AND4_X1   g0904(.A1(new_n363), .A2(new_n644), .A3(new_n911), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1089), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n729), .A2(G330), .A3(new_n825), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n882), .A3(new_n883), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1100), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1106), .B1(new_n1100), .B2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n697), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n905), .A2(new_n907), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1099), .B1(new_n1114), .B2(new_n1097), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1100), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1096), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n644), .A2(new_n911), .A3(new_n363), .A4(new_n1104), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1110), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1100), .A2(new_n1108), .A3(new_n1106), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1113), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g0924(.A(KEYINPUT112), .B(new_n1111), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1112), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1114), .A2(new_n744), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n946), .A2(new_n838), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n261), .B1(new_n786), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G125), .C2(new_n754), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n768), .A2(new_n1033), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1133));
  OAI22_X1  g0933(.A1(new_n1132), .A2(new_n1133), .B1(new_n832), .B2(new_n763), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n774), .A2(G50), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n943), .A2(G128), .B1(new_n760), .B2(G159), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1131), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1065), .B1(new_n754), .B2(G294), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n467), .B2(new_n763), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G97), .A2(new_n766), .B1(new_n765), .B2(G107), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n951), .B2(new_n770), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT115), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n265), .B1(new_n768), .B2(new_n365), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT116), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n1143), .C2(new_n1142), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1138), .B1(new_n835), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n793), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n749), .B1(new_n1066), .B2(new_n852), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(KEYINPUT113), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(KEYINPUT113), .B2(new_n1150), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1119), .A2(new_n992), .B1(new_n1127), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1126), .A2(new_n1153), .ZN(G378));
  NOR2_X1   g0954(.A1(new_n337), .A2(new_n672), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n364), .A2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n364), .A2(new_n1155), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1157), .B2(new_n1156), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1160), .A2(KEYINPUT118), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT118), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1164), .A2(new_n744), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n774), .A2(G58), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n754), .A2(G283), .B1(G97), .B2(new_n765), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(new_n565), .C2(new_n786), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n294), .B(new_n265), .C1(new_n768), .C2(new_n348), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n763), .A2(new_n625), .B1(new_n770), .B2(new_n467), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1168), .A2(new_n941), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1173));
  AOI21_X1  g0973(.A(G50), .B1(new_n546), .B2(new_n294), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n261), .B2(G41), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n946), .A2(new_n832), .B1(new_n768), .B2(new_n1129), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n943), .A2(G125), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n786), .A2(new_n838), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n763), .A2(new_n1180), .B1(new_n759), .B2(new_n1033), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n774), .A2(new_n756), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT59), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n1182), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n793), .B1(new_n1176), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT117), .Z(new_n1191));
  NAND2_X1  g0991(.A1(new_n852), .A2(new_n202), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n739), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1165), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n925), .A2(new_n1164), .A3(G330), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n919), .A2(KEYINPUT40), .B1(new_n921), .B2(new_n923), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n741), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n910), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n910), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1194), .B1(new_n1204), .B2(new_n992), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1105), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1204), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1123), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT112), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1119), .A2(new_n1113), .A3(new_n1123), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1120), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n910), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n910), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n698), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1205), .B1(new_n1207), .B2(new_n1215), .ZN(G375));
  NOR2_X1   g1016(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1120), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n1017), .A3(new_n1111), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n261), .B1(new_n763), .B2(new_n838), .C1(new_n946), .C2(new_n1129), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G50), .B2(new_n760), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n770), .A2(new_n832), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT120), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n786), .A2(new_n1033), .B1(new_n768), .B2(new_n1035), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G128), .B2(new_n754), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1221), .A2(new_n1166), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n261), .B1(new_n775), .B2(G77), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT119), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G107), .A2(new_n766), .B1(new_n765), .B2(G116), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n471), .B2(new_n768), .C1(new_n784), .C2(new_n753), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1037), .B1(new_n951), .B2(new_n763), .C1(new_n547), .C2(new_n770), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1226), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n793), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n749), .B1(new_n253), .B2(new_n852), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n914), .C2(new_n745), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1217), .B2(new_n737), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1219), .A2(new_n1238), .ZN(G381));
  INV_X1    g1039(.A(new_n1205), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n697), .B1(new_n1206), .B2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1241), .B1(new_n1211), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1240), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT121), .ZN(new_n1247));
  INV_X1    g1047(.A(G378), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1058), .A2(new_n805), .A3(new_n1060), .ZN(new_n1252));
  NOR4_X1   g1052(.A1(new_n1251), .A2(new_n1252), .A3(G387), .A4(G381), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1247), .A2(new_n1248), .A3(new_n1253), .ZN(G407));
  NAND2_X1  g1054(.A1(new_n673), .A2(G213), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT122), .Z(new_n1256));
  NAND3_X1  g1056(.A1(new_n1247), .A2(new_n1248), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G407), .A2(new_n1257), .A3(G213), .ZN(G409));
  INV_X1    g1058(.A(KEYINPUT127), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G390), .B(new_n967), .C1(new_n991), .C2(new_n1018), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT124), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n986), .A2(new_n972), .A3(new_n987), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(new_n988), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1052), .A2(new_n993), .A3(new_n1006), .A4(new_n1005), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1016), .B1(new_n1265), .B2(new_n993), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1266), .B2(new_n992), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(KEYINPUT124), .A3(new_n967), .A4(G390), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(new_n1249), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1252), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n805), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1270), .A2(new_n1276), .A3(new_n1273), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1269), .B(new_n1260), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1259), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1270), .A2(new_n1276), .A3(new_n1273), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1276), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1279), .B(new_n1259), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1256), .A2(G2897), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1218), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1217), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n698), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT123), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n697), .B1(new_n1287), .B2(new_n1218), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT123), .A3(new_n1289), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G384), .B1(new_n1295), .B2(new_n1238), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1250), .B(new_n1237), .C1(new_n1292), .C2(new_n1294), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1286), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  AND4_X1   g1098(.A1(KEYINPUT123), .A2(new_n1288), .A3(new_n698), .A4(new_n1289), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT123), .B1(new_n1293), .B2(new_n1289), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1238), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1250), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1295), .A2(G384), .A3(new_n1238), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1255), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1302), .A2(new_n1303), .A3(G2897), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1298), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1206), .A2(new_n1017), .A3(new_n1204), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G378), .B1(new_n1307), .B2(new_n1205), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1246), .B2(G378), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1306), .B1(new_n1309), .B2(new_n1256), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G378), .B(new_n1205), .C1(new_n1207), .C2(new_n1215), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1211), .A2(new_n1244), .A3(new_n1016), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1248), .B1(new_n1312), .B2(new_n1240), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1255), .A4(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1310), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1256), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1315), .B1(new_n1320), .B2(new_n1316), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1285), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1314), .A2(new_n1255), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1316), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1323), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1306), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1320), .A2(KEYINPUT63), .A3(new_n1316), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1322), .A2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1248), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1311), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1316), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1325), .A2(new_n1332), .A3(new_n1311), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1337));
  XNOR2_X1  g1137(.A(new_n1336), .B(new_n1337), .ZN(G402));
endmodule


