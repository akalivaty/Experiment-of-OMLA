//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n191), .B2(G134), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n189), .A3(G137), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT11), .B1(new_n189), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n191), .A3(G134), .ZN(new_n199));
  AOI22_X1  g013(.A1(new_n194), .A2(new_n196), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n193), .B1(new_n200), .B2(new_n188), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  AND4_X1   g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .A4(G128), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(KEYINPUT65), .A3(KEYINPUT1), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n201), .B(KEYINPUT67), .C1(new_n207), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n211), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(G128), .A3(new_n213), .ZN(new_n218));
  INV_X1    g032(.A(new_n208), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n207), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n194), .A2(new_n196), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n197), .A2(new_n199), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n188), .ZN(new_n223));
  INV_X1    g037(.A(new_n193), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n216), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT0), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n208), .B1(new_n227), .B2(new_n209), .ZN(new_n228));
  XOR2_X1   g042(.A(KEYINPUT0), .B(G128), .Z(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n208), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n221), .A2(new_n222), .A3(new_n188), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n188), .B1(new_n221), .B2(new_n222), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n215), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT30), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n223), .B(new_n224), .C1(new_n214), .C2(new_n207), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT30), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n236), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT2), .B(G113), .Z(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT66), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n245), .A3(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n242), .B2(new_n241), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(KEYINPUT68), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n238), .B1(new_n234), .B2(KEYINPUT30), .ZN(new_n251));
  INV_X1    g065(.A(new_n248), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G237), .ZN(new_n254));
  INV_X1    g068(.A(G953), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G210), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(KEYINPUT27), .Z(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT26), .ZN(new_n258));
  INV_X1    g072(.A(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n234), .A2(new_n248), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n249), .A2(new_n253), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n236), .A2(new_n233), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n248), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n252), .A2(new_n233), .A3(new_n236), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n266), .B(new_n269), .C1(new_n261), .C2(new_n268), .ZN(new_n270));
  INV_X1    g084(.A(new_n260), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n262), .B2(KEYINPUT31), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT69), .B1(new_n262), .B2(KEYINPUT31), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n264), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(G472), .A2(G902), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n187), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n270), .A2(new_n271), .ZN(new_n279));
  AND4_X1   g093(.A1(new_n260), .A2(new_n249), .A3(new_n253), .A4(new_n261), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT31), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n262), .A2(KEYINPUT31), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n285), .A3(new_n263), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n276), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n270), .A2(new_n271), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n249), .A2(new_n253), .A3(new_n261), .ZN(new_n289));
  AOI211_X1 g103(.A(KEYINPUT29), .B(new_n288), .C1(new_n271), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n269), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n234), .B(new_n248), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT29), .A3(new_n260), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G472), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n278), .A2(new_n287), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G128), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n300), .A2(KEYINPUT23), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n209), .A2(G119), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(KEYINPUT23), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G110), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT72), .B(G125), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT16), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(G125), .A2(G140), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n308), .B2(G140), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n313), .B2(new_n309), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n314), .A2(new_n203), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n203), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n302), .A2(new_n300), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT24), .B(G110), .Z(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n307), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G125), .B(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n203), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n305), .A2(G110), .B1(new_n318), .B2(new_n319), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(KEYINPUT73), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT22), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(G137), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT73), .B1(new_n321), .B2(new_n325), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT73), .B(new_n330), .C1(new_n321), .C2(new_n325), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n295), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT25), .ZN(new_n336));
  INV_X1    g150(.A(G234), .ZN(new_n337));
  OAI21_X1  g151(.A(G217), .B1(new_n337), .B2(G902), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n338), .B(KEYINPUT70), .Z(new_n339));
  INV_X1    g153(.A(new_n332), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n326), .A3(new_n330), .ZN(new_n341));
  INV_X1    g155(.A(new_n334), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n295), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n339), .A2(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n298), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n230), .A2(new_n308), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n220), .B2(new_n308), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n255), .A2(G224), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n353), .A2(new_n354), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(G110), .B(G122), .Z(new_n359));
  INV_X1    g173(.A(G104), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G107), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n360), .A2(G107), .ZN(new_n363));
  OAI21_X1  g177(.A(G101), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(new_n360), .B2(G107), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G104), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n365), .A2(new_n368), .A3(new_n259), .A4(new_n361), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT5), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n299), .A3(G116), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT80), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(G113), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n247), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n365), .A2(new_n368), .A3(new_n361), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(G101), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(G101), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(new_n386), .A3(G101), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT76), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT76), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n384), .A2(new_n385), .A3(new_n390), .A4(new_n387), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n382), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI211_X1 g206(.A(KEYINPUT81), .B(new_n378), .C1(new_n392), .C2(new_n248), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n394));
  INV_X1    g208(.A(new_n382), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n379), .A2(new_n386), .A3(G101), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n386), .B1(new_n379), .B2(G101), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n390), .B1(new_n398), .B2(new_n385), .ZN(new_n399));
  INV_X1    g213(.A(new_n391), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n395), .B(new_n248), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n394), .B1(new_n401), .B2(new_n377), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n359), .B1(new_n393), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n377), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n403), .B(KEYINPUT6), .C1(new_n359), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n406));
  INV_X1    g220(.A(new_n359), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n394), .A3(new_n377), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n411), .B(new_n359), .C1(new_n393), .C2(new_n402), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT82), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n358), .B(new_n405), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n404), .A2(new_n359), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n355), .A2(KEYINPUT7), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n359), .B(KEYINPUT8), .Z(new_n419));
  AOI21_X1  g233(.A(new_n371), .B1(new_n247), .B2(new_n376), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n378), .B2(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n353), .A2(KEYINPUT7), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n418), .A2(new_n421), .A3(new_n357), .A4(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n416), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n423), .A2(new_n417), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G210), .B1(G237), .B2(G902), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT84), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G469), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n255), .A2(G227), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT74), .Z(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(G110), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(new_n310), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n395), .B(new_n230), .C1(new_n399), .C2(new_n400), .ZN(new_n438));
  INV_X1    g252(.A(new_n207), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n210), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n219), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n370), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n442), .A2(KEYINPUT10), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n371), .B(KEYINPUT10), .C1(new_n214), .C2(new_n207), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n218), .A2(new_n219), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n439), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n448), .A2(KEYINPUT79), .A3(KEYINPUT10), .A4(new_n371), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n438), .A2(new_n443), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n231), .A2(new_n232), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n438), .A2(new_n452), .A3(new_n443), .A4(new_n450), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n437), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n448), .A2(new_n371), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n453), .B1(new_n457), .B2(new_n442), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT12), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n458), .A2(KEYINPUT12), .ZN(new_n460));
  AND4_X1   g274(.A1(new_n455), .A2(new_n437), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n432), .B(new_n295), .C1(new_n456), .C2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n432), .A2(new_n295), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n459), .A3(new_n460), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n436), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n454), .A2(new_n455), .A3(new_n437), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(G469), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G221), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT9), .B(G234), .Z(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n295), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G214), .B1(G237), .B2(G902), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n415), .A2(new_n429), .A3(new_n426), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n431), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G475), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n254), .A2(new_n255), .A3(G214), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(new_n205), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT17), .A3(G131), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(G131), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n480), .B(G143), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n188), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n315), .A2(new_n316), .A3(new_n482), .A4(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n313), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n323), .B1(new_n489), .B2(new_n203), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT18), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n484), .B1(new_n491), .B2(new_n188), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n490), .B(new_n492), .C1(new_n491), .C2(new_n483), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n360), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n488), .A2(new_n496), .A3(new_n493), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n479), .B1(new_n500), .B2(new_n295), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n483), .A2(new_n485), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT19), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n322), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(KEYINPUT19), .B2(new_n313), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n203), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n315), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n493), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n497), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n499), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT85), .ZN(new_n511));
  AOI21_X1  g325(.A(G475), .B1(new_n509), .B2(new_n499), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n295), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n488), .A2(new_n496), .A3(new_n493), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n496), .B1(new_n507), .B2(new_n493), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n479), .B(new_n295), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n509), .B2(new_n499), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n519), .B2(KEYINPUT20), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n501), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(G902), .B(G953), .C1(new_n337), .C2(new_n254), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT88), .Z(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT21), .B(G898), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(KEYINPUT87), .A2(G952), .ZN(new_n526));
  NOR2_X1   g340(.A1(KEYINPUT87), .A2(G952), .ZN(new_n527));
  OAI221_X1 g341(.A(new_n255), .B1(new_n337), .B2(new_n254), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n471), .A2(G217), .A3(new_n255), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT86), .Z(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n205), .A2(G128), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT13), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n209), .A2(G143), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  OAI21_X1  g353(.A(G134), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n534), .A2(new_n537), .A3(new_n189), .ZN(new_n541));
  XNOR2_X1  g355(.A(G116), .B(G122), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n367), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n367), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n540), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G116), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(new_n546), .B2(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(KEYINPUT14), .B2(new_n367), .ZN(new_n549));
  INV_X1    g363(.A(new_n541), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n189), .B1(new_n534), .B2(new_n537), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n533), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n532), .A2(new_n545), .A3(new_n552), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n295), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n557), .B(new_n559), .Z(new_n560));
  NAND3_X1  g374(.A1(new_n521), .A2(new_n530), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n478), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n351), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G101), .ZN(G3));
  INV_X1    g378(.A(G472), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(KEYINPUT89), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n286), .A2(new_n295), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n286), .B2(new_n295), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n350), .A4(new_n475), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n286), .A2(new_n295), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n566), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n575), .A2(new_n350), .A3(new_n568), .A4(new_n475), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT90), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n557), .A2(new_n558), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT91), .B(KEYINPUT33), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n554), .A2(new_n555), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n558), .A2(G902), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT33), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n582), .B(new_n583), .C1(new_n556), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n521), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n431), .A2(new_n477), .ZN(new_n590));
  INV_X1    g404(.A(new_n476), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n590), .A2(new_n529), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n578), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT34), .B(G104), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n501), .B(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n560), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n517), .B(KEYINPUT20), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NOR4_X1   g414(.A1(new_n590), .A2(new_n529), .A3(new_n591), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n578), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G107), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NAND2_X1  g418(.A1(new_n575), .A2(new_n568), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n478), .A2(new_n605), .A3(new_n561), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n321), .A2(new_n325), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n330), .A2(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n347), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n346), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT93), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT37), .B(G110), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G12));
  INV_X1    g429(.A(new_n478), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n528), .B(KEYINPUT94), .Z(new_n617));
  INV_X1    g431(.A(G900), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n523), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n600), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(new_n298), .A3(new_n611), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G128), .ZN(G30));
  XOR2_X1   g436(.A(new_n619), .B(KEYINPUT39), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n475), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT40), .Z(new_n625));
  NOR2_X1   g439(.A1(new_n521), .A2(new_n560), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n611), .A2(new_n627), .A3(new_n591), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT95), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n415), .A2(new_n429), .A3(new_n426), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n429), .B1(new_n415), .B2(new_n426), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n431), .A2(KEYINPUT38), .A3(new_n477), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n289), .A2(new_n260), .ZN(new_n637));
  INV_X1    g451(.A(new_n292), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n638), .B2(new_n271), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n565), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n278), .A2(new_n287), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n625), .A2(new_n629), .A3(new_n636), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n205), .ZN(G45));
  INV_X1    g459(.A(new_n589), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n619), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n616), .A2(new_n298), .A3(new_n611), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G146), .ZN(G48));
  OAI21_X1  g463(.A(new_n295), .B1(new_n456), .B2(new_n461), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(G469), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n473), .A3(new_n462), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n298), .A2(new_n350), .A3(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n631), .A2(new_n632), .A3(new_n591), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n530), .A3(new_n589), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT97), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT41), .B(G113), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G15));
  NAND3_X1  g474(.A1(new_n601), .A2(new_n351), .A3(new_n653), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  INV_X1    g476(.A(new_n561), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n298), .A2(new_n663), .A3(new_n611), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n655), .A2(new_n653), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G119), .ZN(G21));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n631), .A2(new_n632), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n530), .A3(new_n476), .A4(new_n626), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n565), .B1(new_n286), .B2(new_n295), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n276), .B(KEYINPUT98), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n293), .A2(new_n260), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(KEYINPUT31), .B2(new_n262), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n280), .A2(new_n281), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n672), .A2(new_n350), .A3(new_n653), .A4(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n668), .B1(new_n670), .B2(new_n680), .ZN(new_n681));
  NOR4_X1   g495(.A1(new_n671), .A2(new_n349), .A3(new_n652), .A4(new_n678), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n631), .A2(new_n632), .A3(new_n627), .A4(new_n591), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT99), .A4(new_n530), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G122), .ZN(G24));
  AND2_X1   g500(.A1(new_n346), .A2(new_n610), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n671), .A3(new_n678), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(new_n655), .A3(new_n647), .A4(new_n653), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G125), .ZN(G27));
  AND2_X1   g504(.A1(new_n462), .A2(new_n464), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n466), .A2(KEYINPUT100), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n465), .A2(new_n693), .A3(new_n436), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n692), .A2(G469), .A3(new_n467), .A4(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n472), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n590), .A2(new_n476), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n699), .B1(KEYINPUT101), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n699), .B2(new_n700), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n351), .A2(new_n698), .A3(new_n647), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n591), .B1(new_n431), .B2(new_n477), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n298), .A2(new_n704), .A3(new_n350), .A4(new_n696), .ZN(new_n705));
  INV_X1    g519(.A(new_n647), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G131), .ZN(G33));
  INV_X1    g523(.A(new_n705), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n620), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G134), .ZN(G36));
  NAND4_X1  g526(.A1(new_n692), .A2(KEYINPUT45), .A3(new_n467), .A4(new_n694), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n466), .A2(new_n467), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(G469), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT46), .B1(new_n717), .B2(new_n464), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n462), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(KEYINPUT46), .A3(new_n464), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI211_X1 g536(.A(KEYINPUT103), .B(KEYINPUT46), .C1(new_n717), .C2(new_n464), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n472), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n623), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT104), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(KEYINPUT43), .ZN(new_n729));
  INV_X1    g543(.A(new_n501), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n511), .A2(new_n513), .B1(new_n512), .B2(new_n295), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT20), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n730), .B(new_n587), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n728), .A2(KEYINPUT43), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n729), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n521), .B2(new_n587), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT106), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n735), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n605), .B(new_n611), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n704), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n744), .B2(new_n743), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n725), .A2(new_n747), .A3(new_n623), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n727), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT107), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  NAND2_X1  g565(.A1(new_n717), .A2(new_n464), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT103), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n718), .A2(new_n719), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n462), .A3(new_n721), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n758), .A3(new_n473), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n757), .B2(new_n473), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n298), .A2(new_n350), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n647), .A3(new_n704), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT108), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n310), .ZN(G42));
  NAND3_X1  g579(.A1(new_n590), .A2(new_n476), .A3(new_n653), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n617), .B1(new_n735), .B2(new_n738), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n351), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT48), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n255), .B1(new_n526), .B2(new_n527), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n766), .A2(new_n642), .A3(new_n349), .A4(new_n528), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(new_n589), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n651), .A2(new_n472), .A3(new_n462), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n759), .B2(new_n760), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n767), .A2(new_n671), .A3(new_n349), .A4(new_n678), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n704), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(KEYINPUT114), .A3(new_n704), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n635), .A2(KEYINPUT115), .A3(new_n591), .A4(new_n653), .ZN(new_n784));
  NOR2_X1   g598(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n633), .A2(new_n634), .A3(new_n591), .A4(new_n653), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n784), .A2(new_n777), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n768), .A2(new_n688), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n784), .A2(new_n777), .A3(new_n788), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n766), .ZN(new_n795));
  INV_X1    g609(.A(new_n642), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n349), .A2(new_n528), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n795), .A2(new_n521), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT117), .B1(new_n798), .B2(new_n587), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n772), .A2(new_n800), .A3(new_n521), .A4(new_n588), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n783), .A2(new_n789), .A3(new_n794), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n774), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n777), .A2(new_n655), .A3(new_n653), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n780), .A2(new_n781), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT47), .B1(new_n724), .B2(new_n472), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n757), .A2(new_n758), .A3(new_n473), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n807), .B1(new_n810), .B2(new_n775), .ZN(new_n811));
  INV_X1    g625(.A(new_n788), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n777), .B1(new_n786), .B2(new_n787), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n793), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n790), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT51), .A3(new_n789), .A4(new_n802), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n805), .A2(new_n806), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n619), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n560), .A2(new_n597), .A3(new_n599), .A4(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n476), .C1(new_n631), .C2(new_n632), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n590), .A2(KEYINPUT109), .A3(new_n476), .A4(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n298), .A2(new_n475), .A3(new_n611), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(KEYINPUT110), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n620), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n688), .A2(new_n647), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n705), .A2(new_n832), .B1(new_n833), .B2(new_n697), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n708), .A3(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n656), .A2(new_n654), .B1(new_n664), .B2(new_n665), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n655), .A2(new_n530), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n654), .A2(new_n838), .A3(new_n600), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n606), .A2(new_n611), .B1(new_n351), .B2(new_n562), .ZN(new_n841));
  INV_X1    g655(.A(new_n521), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n646), .B1(new_n560), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n573), .A2(new_n577), .A3(new_n592), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n840), .A2(new_n685), .A3(new_n841), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT111), .B1(new_n836), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n685), .A3(new_n844), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n657), .A2(new_n666), .A3(new_n661), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n834), .B1(new_n829), .B2(new_n830), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n708), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n611), .A2(new_n619), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n683), .A2(new_n642), .A3(new_n696), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n621), .A2(new_n648), .A3(new_n855), .A4(new_n689), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n856), .B(new_n857), .C1(new_n859), .C2(new_n860), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n859), .B1(new_n856), .B2(new_n860), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n846), .A2(new_n852), .A3(new_n853), .A4(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n841), .A2(new_n685), .A3(new_n844), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n851), .A2(new_n867), .A3(new_n708), .A4(new_n840), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n856), .B(KEYINPUT52), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT53), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n866), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n831), .A2(new_n708), .A3(new_n835), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n865), .A2(new_n872), .A3(KEYINPUT53), .A4(new_n849), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n853), .B1(new_n868), .B2(new_n869), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n818), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n818), .A2(new_n871), .A3(KEYINPUT118), .A4(new_n876), .ZN(new_n880));
  NOR2_X1   g694(.A1(G952), .A2(G953), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT119), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n651), .A2(new_n462), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n349), .B1(KEYINPUT49), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(KEYINPUT49), .B2(new_n884), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n642), .A2(new_n886), .A3(new_n472), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n733), .A2(new_n591), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n635), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n883), .A2(new_n889), .ZN(G75));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n873), .A2(new_n874), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(G902), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(new_n430), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n405), .B1(new_n412), .B2(new_n414), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n358), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT55), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n255), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n897), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n891), .B(new_n901), .C1(new_n893), .C2(new_n430), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n900), .A3(new_n902), .ZN(G51));
  XNOR2_X1  g717(.A(new_n463), .B(KEYINPUT57), .ZN(new_n904));
  INV_X1    g718(.A(new_n876), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n875), .B1(new_n873), .B2(new_n874), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n456), .B2(new_n461), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n893), .A2(new_n717), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  INV_X1    g725(.A(new_n510), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n899), .ZN(G60));
  NOR2_X1   g729(.A1(new_n556), .A2(new_n585), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n556), .B2(new_n581), .ZN(new_n917));
  XNOR2_X1  g731(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n558), .A2(new_n295), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n917), .B(new_n920), .C1(new_n905), .C2(new_n906), .ZN(new_n921));
  INV_X1    g735(.A(new_n920), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n871), .B2(new_n876), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n921), .B(new_n900), .C1(new_n917), .C2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT60), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n892), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n343), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n899), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n927), .B1(new_n873), .B2(new_n874), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n609), .B(KEYINPUT121), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n931), .A2(new_n933), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n900), .B1(new_n935), .B2(new_n343), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n892), .A2(new_n928), .A3(new_n936), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n932), .B(KEYINPUT61), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n524), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n849), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n895), .B1(G898), .B2(new_n255), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  XNOR2_X1  g761(.A(new_n251), .B(KEYINPUT123), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(new_n505), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(G900), .A2(G953), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n727), .A2(new_n351), .A3(new_n683), .A4(new_n748), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n952), .A2(new_n708), .A3(new_n711), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n749), .A2(new_n763), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n621), .A2(new_n648), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n689), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n950), .B(new_n951), .C1(new_n957), .C2(G953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n643), .A2(new_n955), .A3(new_n689), .A4(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n624), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n351), .A2(new_n964), .A3(new_n704), .A4(new_n843), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n749), .A2(new_n763), .A3(new_n963), .A4(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n969));
  AOI22_X1  g783(.A1(new_n956), .A2(new_n643), .B1(new_n962), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n965), .A2(new_n966), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n949), .B1(new_n972), .B2(G953), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n958), .A2(new_n961), .A3(new_n973), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n959), .A2(new_n960), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G72));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n972), .B2(new_n849), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n289), .A2(new_n260), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n866), .A2(new_n870), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n637), .A2(new_n978), .ZN(new_n983));
  OAI22_X1  g797(.A1(new_n980), .A2(new_n637), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n953), .A2(new_n954), .A3(new_n956), .A4(new_n849), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n981), .B1(new_n985), .B2(new_n978), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n987));
  OR3_X1    g801(.A1(new_n986), .A2(new_n987), .A3(new_n899), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n986), .B2(new_n899), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(G57));
endmodule


