

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596;

  NOR2_X1 U319 ( .A1(n563), .A2(n562), .ZN(n575) );
  AND2_X1 U320 ( .A1(G227GAT), .A2(G233GAT), .ZN(n287) );
  XOR2_X1 U321 ( .A(n557), .B(n556), .Z(n288) );
  XNOR2_X1 U322 ( .A(n387), .B(n386), .ZN(n563) );
  NOR2_X1 U323 ( .A1(n574), .A2(n517), .ZN(n518) );
  XNOR2_X1 U324 ( .A(n443), .B(n287), .ZN(n370) );
  INV_X1 U325 ( .A(G64GAT), .ZN(n444) );
  XNOR2_X1 U326 ( .A(n370), .B(n389), .ZN(n373) );
  XNOR2_X1 U327 ( .A(n445), .B(n444), .ZN(n446) );
  NOR2_X1 U328 ( .A1(n511), .A2(n559), .ZN(n403) );
  XNOR2_X1 U329 ( .A(n447), .B(n446), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n525), .B(n524), .ZN(n554) );
  XNOR2_X1 U331 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U332 ( .A(n590), .B(KEYINPUT109), .ZN(n570) );
  XNOR2_X1 U333 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(n590) );
  XNOR2_X1 U335 ( .A(n461), .B(n460), .ZN(n488) );
  XNOR2_X1 U336 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U337 ( .A(n465), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT67), .B(G8GAT), .Z(n290) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(G15GAT), .ZN(n289) );
  XNOR2_X1 U340 ( .A(n290), .B(n289), .ZN(n311) );
  XOR2_X1 U341 ( .A(G113GAT), .B(G141GAT), .Z(n292) );
  XNOR2_X1 U342 ( .A(G197GAT), .B(G22GAT), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n294) );
  XOR2_X1 U344 ( .A(G36GAT), .B(G50GAT), .Z(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n302) );
  XNOR2_X1 U346 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n295), .B(KEYINPUT29), .ZN(n296) );
  XOR2_X1 U348 ( .A(n296), .B(KEYINPUT71), .Z(n301) );
  XOR2_X1 U349 ( .A(G29GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U350 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n342) );
  XNOR2_X1 U352 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n299), .B(KEYINPUT70), .ZN(n453) );
  XNOR2_X1 U354 ( .A(n342), .B(n453), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n303) );
  NAND2_X1 U356 ( .A1(n302), .A2(n303), .ZN(n307) );
  INV_X1 U357 ( .A(n302), .ZN(n305) );
  INV_X1 U358 ( .A(n303), .ZN(n304) );
  NAND2_X1 U359 ( .A1(n305), .A2(n304), .ZN(n306) );
  NAND2_X1 U360 ( .A1(n307), .A2(n306), .ZN(n309) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X2 U363 ( .A(n311), .B(n310), .Z(n564) );
  XOR2_X1 U364 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n313) );
  NAND2_X1 U365 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U367 ( .A(n314), .B(KEYINPUT74), .Z(n319) );
  XNOR2_X1 U368 ( .A(G71GAT), .B(G57GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n315), .B(KEYINPUT13), .ZN(n452) );
  XOR2_X1 U370 ( .A(G64GAT), .B(G92GAT), .Z(n317) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n390) );
  XNOR2_X1 U373 ( .A(n452), .B(n390), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U375 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n321) );
  XNOR2_X1 U376 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U378 ( .A(n323), .B(n322), .Z(n327) );
  XNOR2_X1 U379 ( .A(G106GAT), .B(G78GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n324), .B(G148GAT), .ZN(n361) );
  XNOR2_X1 U381 ( .A(G99GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n325), .B(KEYINPUT73), .ZN(n341) );
  XNOR2_X1 U383 ( .A(n361), .B(n341), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n587) );
  NAND2_X1 U385 ( .A1(n564), .A2(n587), .ZN(n471) );
  XOR2_X1 U386 ( .A(KEYINPUT66), .B(KEYINPUT77), .Z(n329) );
  XNOR2_X1 U387 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U389 ( .A(KEYINPUT64), .B(KEYINPUT65), .Z(n331) );
  XNOR2_X1 U390 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n346) );
  XOR2_X1 U393 ( .A(G36GAT), .B(G190GAT), .Z(n397) );
  XNOR2_X1 U394 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n334), .B(G162GAT), .ZN(n352) );
  XOR2_X1 U396 ( .A(n397), .B(n352), .Z(n336) );
  NAND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U399 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n338) );
  XNOR2_X1 U400 ( .A(G134GAT), .B(G106GAT), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U402 ( .A(n340), .B(n339), .Z(n344) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n574) );
  XOR2_X1 U406 ( .A(KEYINPUT36), .B(n574), .Z(n593) );
  XOR2_X1 U407 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XNOR2_X1 U408 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT2), .ZN(n418) );
  XOR2_X1 U410 ( .A(n436), .B(n418), .Z(n349) );
  NAND2_X1 U411 ( .A1(G228GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n351) );
  INV_X1 U413 ( .A(G204GAT), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n352), .B(G211GAT), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U417 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n356) );
  XNOR2_X1 U418 ( .A(KEYINPUT84), .B(KEYINPUT23), .ZN(n355) );
  XOR2_X1 U419 ( .A(n356), .B(n355), .Z(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U421 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n360) );
  XNOR2_X1 U422 ( .A(G197GAT), .B(G218GAT), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n391) );
  XNOR2_X1 U424 ( .A(n361), .B(n391), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n559) );
  XOR2_X1 U426 ( .A(G15GAT), .B(G127GAT), .Z(n443) );
  INV_X1 U427 ( .A(KEYINPUT18), .ZN(n364) );
  NAND2_X1 U428 ( .A1(n364), .A2(KEYINPUT19), .ZN(n367) );
  INV_X1 U429 ( .A(KEYINPUT19), .ZN(n365) );
  NAND2_X1 U430 ( .A1(n365), .A2(KEYINPUT18), .ZN(n366) );
  NAND2_X1 U431 ( .A1(n367), .A2(n366), .ZN(n369) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n389) );
  INV_X1 U434 ( .A(n373), .ZN(n371) );
  NAND2_X1 U435 ( .A1(n371), .A2(G71GAT), .ZN(n375) );
  INV_X1 U436 ( .A(G71GAT), .ZN(n372) );
  NAND2_X1 U437 ( .A1(n373), .A2(n372), .ZN(n374) );
  NAND2_X1 U438 ( .A1(n375), .A2(n374), .ZN(n387) );
  XOR2_X1 U439 ( .A(KEYINPUT20), .B(G99GAT), .Z(n377) );
  XNOR2_X1 U440 ( .A(G43GAT), .B(G190GAT), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U442 ( .A(G183GAT), .B(KEYINPUT83), .Z(n379) );
  XNOR2_X1 U443 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U445 ( .A(n381), .B(n380), .Z(n385) );
  XOR2_X1 U446 ( .A(G120GAT), .B(KEYINPUT0), .Z(n383) );
  XNOR2_X1 U447 ( .A(G113GAT), .B(G134GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n419) );
  XNOR2_X1 U449 ( .A(n419), .B(G176GAT), .ZN(n384) );
  INV_X1 U450 ( .A(n563), .ZN(n511) );
  XNOR2_X1 U451 ( .A(G8GAT), .B(G183GAT), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n388), .B(G211GAT), .ZN(n437) );
  XNOR2_X1 U453 ( .A(n389), .B(n437), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n393) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U458 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n555) );
  NAND2_X1 U461 ( .A1(n511), .A2(n555), .ZN(n400) );
  XOR2_X1 U462 ( .A(KEYINPUT93), .B(n400), .Z(n401) );
  NAND2_X1 U463 ( .A1(n559), .A2(n401), .ZN(n402) );
  XNOR2_X1 U464 ( .A(KEYINPUT25), .B(n402), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n403), .B(KEYINPUT26), .ZN(n405) );
  INV_X1 U466 ( .A(KEYINPUT91), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n580) );
  XNOR2_X1 U468 ( .A(n555), .B(KEYINPUT90), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n406), .B(KEYINPUT27), .ZN(n430) );
  NAND2_X1 U470 ( .A1(n580), .A2(n430), .ZN(n542) );
  INV_X1 U471 ( .A(KEYINPUT92), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n542), .B(n407), .ZN(n408) );
  NOR2_X1 U473 ( .A1(n409), .A2(n408), .ZN(n428) );
  XOR2_X1 U474 ( .A(KEYINPUT6), .B(KEYINPUT86), .Z(n411) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(G57GAT), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n427) );
  XOR2_X1 U477 ( .A(G155GAT), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U478 ( .A(G127GAT), .B(G148GAT), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U480 ( .A(G29GAT), .B(G85GAT), .Z(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n423) );
  XNOR2_X1 U482 ( .A(KEYINPUT5), .B(KEYINPUT87), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n416), .B(KEYINPUT4), .ZN(n417) );
  XOR2_X1 U484 ( .A(n417), .B(KEYINPUT1), .Z(n421) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n425) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n558) );
  NOR2_X1 U491 ( .A1(n428), .A2(n558), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n429), .B(KEYINPUT94), .ZN(n434) );
  XOR2_X1 U493 ( .A(n559), .B(KEYINPUT28), .Z(n506) );
  INV_X1 U494 ( .A(n430), .ZN(n431) );
  NOR2_X1 U495 ( .A1(n506), .A2(n431), .ZN(n432) );
  NAND2_X1 U496 ( .A1(n432), .A2(n558), .ZN(n512) );
  NOR2_X1 U497 ( .A1(n512), .A2(n511), .ZN(n433) );
  NOR2_X1 U498 ( .A1(n434), .A2(n433), .ZN(n469) );
  NOR2_X1 U499 ( .A1(n593), .A2(n469), .ZN(n456) );
  INV_X1 U500 ( .A(n437), .ZN(n435) );
  NAND2_X1 U501 ( .A1(n436), .A2(n435), .ZN(n440) );
  INV_X1 U502 ( .A(n436), .ZN(n438) );
  NAND2_X1 U503 ( .A1(n438), .A2(n437), .ZN(n439) );
  NAND2_X1 U504 ( .A1(n440), .A2(n439), .ZN(n442) );
  NAND2_X1 U505 ( .A1(G231GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n443), .B(G78GAT), .ZN(n445) );
  XOR2_X1 U508 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n449) );
  XNOR2_X1 U509 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U511 ( .A(n451), .B(n450), .Z(n455) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U513 ( .A1(n456), .A2(n590), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT37), .B(n457), .Z(n501) );
  NOR2_X1 U515 ( .A1(n471), .A2(n501), .ZN(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n459) );
  INV_X1 U517 ( .A(KEYINPUT100), .ZN(n458) );
  AND2_X1 U518 ( .A1(n488), .A2(n511), .ZN(n465) );
  XNOR2_X1 U519 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n463) );
  INV_X1 U520 ( .A(G43GAT), .ZN(n462) );
  XNOR2_X1 U521 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n574), .A2(n590), .ZN(n466) );
  XOR2_X1 U523 ( .A(n467), .B(n466), .Z(n468) );
  NOR2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U525 ( .A(KEYINPUT95), .B(n470), .ZN(n491) );
  NOR2_X1 U526 ( .A1(n471), .A2(n491), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT96), .ZN(n479) );
  NAND2_X1 U528 ( .A1(n479), .A2(n558), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n473), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n474), .ZN(G1324GAT) );
  XOR2_X1 U531 ( .A(G8GAT), .B(KEYINPUT97), .Z(n476) );
  NAND2_X1 U532 ( .A1(n555), .A2(n479), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U535 ( .A1(n511), .A2(n479), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NAND2_X1 U537 ( .A1(n479), .A2(n506), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT98), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(G29GAT), .B(KEYINPUT99), .Z(n483) );
  NAND2_X1 U541 ( .A1(n488), .A2(n558), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n485) );
  XOR2_X1 U543 ( .A(KEYINPUT39), .B(KEYINPUT102), .Z(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  XOR2_X1 U545 ( .A(G36GAT), .B(KEYINPUT103), .Z(n487) );
  NAND2_X1 U546 ( .A1(n488), .A2(n555), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(G1329GAT) );
  XOR2_X1 U548 ( .A(G50GAT), .B(KEYINPUT105), .Z(n490) );
  NAND2_X1 U549 ( .A1(n488), .A2(n506), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(G1331GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n493) );
  INV_X1 U552 ( .A(n564), .ZN(n582) );
  XNOR2_X1 U553 ( .A(n587), .B(KEYINPUT41), .ZN(n566) );
  NAND2_X1 U554 ( .A1(n582), .A2(n566), .ZN(n500) );
  NOR2_X1 U555 ( .A1(n491), .A2(n500), .ZN(n497) );
  NAND2_X1 U556 ( .A1(n497), .A2(n558), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U558 ( .A(G57GAT), .B(n494), .Z(G1332GAT) );
  NAND2_X1 U559 ( .A1(n497), .A2(n555), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n495), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U561 ( .A1(n497), .A2(n511), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n496), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U563 ( .A(G78GAT), .B(KEYINPUT43), .Z(n499) );
  NAND2_X1 U564 ( .A1(n497), .A2(n506), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(G1335GAT) );
  NOR2_X1 U566 ( .A1(n501), .A2(n500), .ZN(n507) );
  NAND2_X1 U567 ( .A1(n507), .A2(n558), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G85GAT), .B(n502), .ZN(G1336GAT) );
  XOR2_X1 U569 ( .A(G92GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U570 ( .A1(n507), .A2(n555), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1337GAT) );
  NAND2_X1 U572 ( .A1(n507), .A2(n511), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n509) );
  NAND2_X1 U575 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U577 ( .A(G106GAT), .B(n510), .Z(G1339GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n529) );
  NOR2_X1 U579 ( .A1(n563), .A2(n512), .ZN(n526) );
  AND2_X1 U580 ( .A1(n566), .A2(n564), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n513), .B(KEYINPUT46), .ZN(n514) );
  NOR2_X1 U582 ( .A1(n570), .A2(n514), .ZN(n516) );
  INV_X1 U583 ( .A(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(KEYINPUT47), .ZN(n523) );
  NOR2_X1 U586 ( .A1(n593), .A2(n590), .ZN(n519) );
  XOR2_X1 U587 ( .A(KEYINPUT45), .B(n519), .Z(n520) );
  NOR2_X1 U588 ( .A1(n564), .A2(n520), .ZN(n521) );
  NAND2_X1 U589 ( .A1(n521), .A2(n587), .ZN(n522) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n525) );
  XOR2_X1 U591 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n524) );
  NAND2_X1 U592 ( .A1(n526), .A2(n554), .ZN(n527) );
  XOR2_X1 U593 ( .A(KEYINPUT112), .B(n527), .Z(n537) );
  NAND2_X1 U594 ( .A1(n564), .A2(n537), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U598 ( .A1(n537), .A2(n566), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n535) );
  NAND2_X1 U602 ( .A1(n537), .A2(n570), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n539) );
  NAND2_X1 U606 ( .A1(n574), .A2(n537), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n540), .Z(G1343GAT) );
  NAND2_X1 U609 ( .A1(n554), .A2(n558), .ZN(n541) );
  NOR2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n552), .A2(n564), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n543), .B(KEYINPUT118), .ZN(n544) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n546) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(n547), .Z(n549) );
  NAND2_X1 U618 ( .A1(n552), .A2(n566), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  INV_X1 U620 ( .A(n590), .ZN(n550) );
  NAND2_X1 U621 ( .A1(n552), .A2(n550), .ZN(n551) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n552), .A2(n574), .ZN(n553) );
  XNOR2_X1 U624 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n555), .A2(n554), .ZN(n557) );
  XOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n556) );
  INV_X1 U627 ( .A(n558), .ZN(n579) );
  AND2_X1 U628 ( .A1(n559), .A2(n579), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n288), .A2(n560), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT55), .B(n561), .Z(n562) );
  NAND2_X1 U631 ( .A1(n564), .A2(n575), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  NAND2_X1 U634 ( .A1(n575), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n572) );
  NAND2_X1 U638 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(n573), .ZN(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n577) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(G190GAT), .B(n578), .Z(G1351GAT) );
  AND2_X1 U645 ( .A1(n288), .A2(n579), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n592) );
  NOR2_X1 U647 ( .A1(n592), .A2(n582), .ZN(n586) );
  XOR2_X1 U648 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  NOR2_X1 U652 ( .A1(n587), .A2(n592), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1353GAT) );
  NOR2_X1 U655 ( .A1(n590), .A2(n592), .ZN(n591) );
  XOR2_X1 U656 ( .A(G211GAT), .B(n591), .Z(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XOR2_X1 U660 ( .A(G218GAT), .B(n596), .Z(G1355GAT) );
endmodule

