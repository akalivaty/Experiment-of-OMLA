//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  AND2_X1   g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n209), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT0), .Z(new_n234));
  NOR4_X1   g0034(.A1(new_n225), .A2(new_n226), .A3(new_n231), .A4(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n202), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n211), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT84), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G257), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G303), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(G1698), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n260), .B(new_n264), .C1(new_n265), .C2(new_n220), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n229), .B1(KEYINPUT66), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n206), .A2(G45), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT5), .A2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT5), .A2(G41), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n272), .A2(G274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n276), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(new_n272), .A3(G270), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n268), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT83), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n268), .A2(KEYINPUT83), .A3(new_n277), .A4(new_n279), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G200), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n285), .A2(new_n207), .A3(G1), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G116), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n229), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n290), .B(new_n286), .C1(new_n206), .C2(G33), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(new_n291), .B2(G116), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G283), .ZN(new_n293));
  INV_X1    g0093(.A(G97), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(new_n207), .C1(G33), .C2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n290), .C1(new_n207), .C2(G116), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT20), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n296), .B(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n284), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n282), .B2(new_n283), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n253), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n302), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n304), .A2(KEYINPUT84), .A3(new_n284), .A4(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n258), .A2(new_n207), .A3(G87), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT22), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT22), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n258), .A2(new_n309), .A3(new_n207), .A4(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G116), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G20), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n207), .B2(G107), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n219), .A2(KEYINPUT23), .A3(G20), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n311), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n312), .B1(new_n311), .B2(new_n318), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n290), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT25), .B1(new_n286), .B2(new_n219), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n291), .A2(G107), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n258), .A2(G257), .A3(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G33), .A2(G294), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n258), .A2(new_n259), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n214), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n267), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n278), .A2(new_n272), .A3(G264), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n277), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n333), .A2(G179), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n326), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n292), .B2(new_n298), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n282), .A2(new_n283), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT21), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n268), .A2(G179), .A3(new_n277), .A4(new_n279), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n299), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n282), .A2(KEYINPUT21), .A3(new_n338), .A4(new_n283), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n337), .A2(new_n341), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n306), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n258), .A2(G250), .A3(G1698), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n258), .A2(G244), .A3(new_n259), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT4), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n293), .B(new_n347), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n263), .A2(G1698), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT4), .B1(new_n351), .B2(G244), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n267), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n278), .A2(new_n272), .A3(G257), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n354), .A2(new_n277), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT81), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(KEYINPUT81), .A3(new_n355), .ZN(new_n359));
  AOI21_X1  g0159(.A(G169), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n356), .A2(G179), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n287), .A2(G97), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n291), .B2(G97), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(G97), .A3(new_n219), .ZN(new_n366));
  XOR2_X1   g0166(.A(G97), .B(G107), .Z(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G20), .A2(G33), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(G20), .B1(G77), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n256), .A2(new_n207), .A3(new_n257), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n257), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT76), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(G107), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT80), .B1(new_n380), .B2(new_n290), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT80), .ZN(new_n382));
  INV_X1    g0182(.A(new_n290), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n382), .B(new_n383), .C1(new_n370), .C2(new_n379), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n364), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n362), .A2(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n381), .A2(new_n384), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n356), .A2(G200), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n358), .A2(G190), .A3(new_n359), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n387), .A2(new_n364), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n331), .A2(new_n332), .A3(G190), .A4(new_n277), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n333), .A2(G200), .ZN(new_n392));
  AND4_X1   g0192(.A1(new_n321), .A2(new_n325), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n258), .A2(G238), .A3(new_n259), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n313), .C1(new_n265), .C2(new_n218), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n267), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n273), .A2(new_n214), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n272), .B(new_n397), .C1(G274), .C2(new_n273), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G200), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n207), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n213), .A2(new_n294), .A3(new_n219), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n258), .A2(new_n207), .A3(G68), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n207), .A2(G33), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n401), .B1(new_n294), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT15), .B(G87), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n409), .A2(new_n290), .B1(new_n286), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n291), .A2(G87), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n396), .A2(G190), .A3(new_n398), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n400), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n290), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(new_n286), .ZN(new_n416));
  INV_X1    g0216(.A(new_n410), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n291), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n399), .A2(new_n334), .ZN(new_n420));
  INV_X1    g0220(.A(G179), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n396), .A2(new_n421), .A3(new_n398), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n393), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n386), .A2(new_n390), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n346), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n428));
  INV_X1    g0228(.A(G222), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n428), .B1(new_n217), .B2(new_n258), .C1(new_n329), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n267), .ZN(new_n431));
  INV_X1    g0231(.A(G41), .ZN(new_n432));
  INV_X1    g0232(.A(G45), .ZN(new_n433));
  AOI21_X1  g0233(.A(G1), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n272), .A2(G274), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n270), .B2(new_n271), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G226), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G200), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT10), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n431), .A2(G190), .A3(new_n435), .A4(new_n437), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT9), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n407), .B(KEYINPUT67), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT8), .B(G58), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n369), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n383), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n286), .A2(new_n290), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT68), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n207), .B2(G1), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n206), .A2(KEYINPUT68), .A3(G20), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n202), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n450), .A2(new_n454), .B1(new_n202), .B2(new_n286), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n443), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n448), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n444), .B2(new_n446), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT9), .B(new_n455), .C1(new_n459), .C2(new_n383), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n442), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n441), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT72), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n442), .A2(new_n457), .A3(KEYINPUT72), .A4(new_n460), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(new_n439), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT10), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT73), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT73), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n469), .A3(KEYINPUT10), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n462), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G232), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G1698), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(G226), .B2(G1698), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n402), .B1(new_n474), .B2(new_n263), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n267), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n436), .A2(G238), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n435), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT13), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n478), .A2(KEYINPUT13), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT14), .B1(new_n482), .B2(new_n334), .ZN(new_n483));
  INV_X1    g0283(.A(new_n481), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n479), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT14), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(G169), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n483), .B(new_n487), .C1(new_n421), .C2(new_n485), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n369), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n489));
  INV_X1    g0289(.A(new_n444), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n217), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT11), .A3(new_n290), .ZN(new_n492));
  OR3_X1    g0292(.A1(new_n287), .A2(KEYINPUT12), .A3(G68), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT12), .B1(new_n287), .B2(G68), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n452), .A2(new_n453), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n211), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n493), .A2(new_n494), .B1(new_n497), .B2(new_n450), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT11), .B1(new_n491), .B2(new_n290), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT75), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n488), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n485), .B2(new_n301), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT74), .ZN(new_n505));
  INV_X1    g0305(.A(G200), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n505), .B1(new_n482), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n485), .A2(KEYINPUT74), .A3(G200), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n438), .A2(new_n334), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n455), .B1(new_n459), .B2(new_n383), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(G179), .C2(new_n438), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT69), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n446), .A2(new_n369), .B1(G20), .B2(G77), .ZN(new_n515));
  INV_X1    g0315(.A(new_n407), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n417), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n383), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n450), .A2(G77), .A3(new_n495), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G77), .B2(new_n287), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n436), .A2(G244), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n522), .A2(new_n435), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n263), .A2(G107), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n265), .B2(new_n212), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT70), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n329), .B2(new_n472), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n351), .A2(KEYINPUT70), .A3(G232), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n267), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n521), .B1(new_n531), .B2(new_n334), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n527), .A2(new_n528), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n267), .B1(new_n533), .B2(new_n525), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n534), .A2(KEYINPUT71), .A3(new_n421), .A4(new_n523), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n421), .B(new_n523), .C1(new_n529), .C2(new_n530), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n532), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n534), .A2(G190), .A3(new_n523), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n531), .A2(G200), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(new_n521), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n503), .A2(new_n510), .A3(new_n514), .A4(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n496), .A2(new_n445), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n450), .B1(new_n286), .B2(new_n445), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n376), .A2(G68), .A3(new_n378), .ZN(new_n547));
  INV_X1    g0347(.A(G58), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n211), .ZN(new_n549));
  OAI21_X1  g0349(.A(G20), .B1(new_n549), .B2(new_n201), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n369), .A2(G159), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT16), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT7), .B1(new_n263), .B2(new_n207), .ZN(new_n555));
  OAI21_X1  g0355(.A(G68), .B1(new_n555), .B2(new_n377), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(KEYINPUT16), .A3(new_n553), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n290), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n546), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(KEYINPUT77), .B(new_n546), .C1(new_n554), .C2(new_n558), .ZN(new_n562));
  INV_X1    g0362(.A(new_n434), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n272), .A2(G232), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n435), .A2(new_n564), .ZN(new_n565));
  OR2_X1    g0365(.A1(G223), .A2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(G226), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(G1698), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n566), .B(new_n568), .C1(new_n261), .C2(new_n262), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT78), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n569), .A2(new_n573), .A3(new_n570), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n267), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G169), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n421), .B2(new_n576), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n561), .A2(new_n562), .A3(new_n578), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n579), .A2(KEYINPUT18), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n506), .B1(new_n565), .B2(new_n575), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n565), .A2(new_n575), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(G190), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n546), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n547), .A2(new_n553), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT16), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n373), .A2(new_n375), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n552), .B1(new_n588), .B2(G68), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n383), .B1(new_n589), .B2(KEYINPUT16), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n584), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT17), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n579), .A2(KEYINPUT18), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n580), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR4_X1   g0395(.A1(new_n427), .A2(new_n471), .A3(new_n544), .A4(new_n595), .ZN(G372));
  INV_X1    g0396(.A(new_n514), .ZN(new_n597));
  INV_X1    g0397(.A(new_n462), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n466), .A2(new_n469), .A3(KEYINPUT10), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n469), .B1(new_n466), .B2(KEYINPUT10), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT88), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n603), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n565), .A2(new_n575), .A3(G179), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n334), .B1(new_n565), .B2(new_n575), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT87), .B1(new_n591), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n578), .A2(new_n610), .A3(new_n559), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n609), .A2(new_n611), .A3(KEYINPUT18), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n509), .A2(new_n539), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n502), .B2(new_n488), .ZN(new_n618));
  INV_X1    g0418(.A(new_n593), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n597), .B1(new_n605), .B2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n471), .A2(new_n544), .A3(new_n595), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n345), .A2(new_n386), .A3(new_n390), .A4(new_n425), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n423), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n414), .A2(new_n423), .ZN(new_n625));
  AND4_X1   g0425(.A1(KEYINPUT26), .A2(new_n362), .A3(new_n625), .A4(new_n385), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n358), .A2(new_n359), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n334), .ZN(new_n629));
  INV_X1    g0429(.A(new_n361), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(KEYINPUT86), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT86), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n360), .B2(new_n361), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n631), .A2(new_n633), .A3(new_n385), .A4(new_n625), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n626), .B1(new_n627), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n622), .B1(new_n624), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n621), .A2(new_n636), .ZN(G369));
  NAND3_X1  g0437(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(KEYINPUT27), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G213), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n299), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT89), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n306), .A2(new_n638), .A3(new_n645), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n644), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n393), .B1(new_n326), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n337), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n337), .A2(new_n652), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n638), .A2(new_n644), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n656), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n232), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n404), .A2(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n227), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n331), .A2(new_n332), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n342), .A2(new_n399), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n358), .A3(new_n359), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n671), .A2(KEYINPUT30), .A3(new_n358), .A4(new_n359), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n356), .A2(new_n333), .ZN(new_n677));
  AOI21_X1  g0477(.A(G179), .B1(new_n396), .B2(new_n398), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n282), .A2(new_n283), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT90), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n282), .A2(new_n681), .A3(new_n283), .A4(new_n678), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n652), .B1(new_n676), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT31), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT31), .B(new_n652), .C1(new_n676), .C2(new_n683), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n686), .B(new_n687), .C1(new_n427), .C2(new_n652), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n424), .B1(new_n387), .B2(new_n364), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(KEYINPUT26), .A3(new_n633), .A4(new_n631), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n625), .A2(new_n385), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n629), .A2(new_n630), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n627), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n423), .A3(new_n623), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .A3(new_n644), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n644), .B1(new_n635), .B2(new_n624), .ZN(new_n699));
  XOR2_X1   g0499(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n690), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n669), .B1(new_n702), .B2(G1), .ZN(G364));
  NOR2_X1   g0503(.A1(new_n285), .A2(G20), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n206), .B1(new_n704), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n664), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n232), .A2(new_n258), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT92), .Z(new_n710));
  INV_X1    g0510(.A(G116), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n710), .A2(G355), .B1(new_n711), .B2(new_n663), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n251), .A2(new_n433), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n663), .A2(new_n258), .ZN(new_n714));
  INV_X1    g0514(.A(new_n228), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(G45), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n712), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n229), .B1(G20), .B2(new_n334), .ZN(new_n718));
  NOR3_X1   g0518(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n708), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n718), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n207), .A2(new_n421), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n724), .A2(new_n506), .A3(G190), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n301), .A2(G179), .A3(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n207), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(G68), .A2(new_n725), .B1(new_n728), .B2(G97), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT93), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n301), .A2(new_n506), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n207), .A2(G179), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G87), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n724), .A2(new_n301), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n737), .B2(new_n548), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(new_n301), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G107), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G190), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT32), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n258), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n723), .A2(new_n731), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n723), .A2(new_n742), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n747), .A2(new_n202), .B1(new_n748), .B2(new_n217), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n743), .A2(KEYINPUT32), .A3(new_n744), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n738), .A2(new_n746), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n743), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n736), .A2(G322), .B1(G329), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n747), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n258), .B1(new_n754), .B2(G326), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(G294), .B2(new_n728), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n739), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G303), .ZN(new_n760));
  INV_X1    g0560(.A(G311), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n733), .B1(new_n748), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n759), .B(new_n762), .C1(new_n725), .C2(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n730), .A2(new_n751), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n721), .B1(new_n722), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT94), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n719), .B(KEYINPUT95), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n649), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT96), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n649), .A2(G330), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n771), .A2(new_n650), .A3(new_n708), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(G396));
  NAND2_X1  g0574(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n623), .A2(new_n423), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n634), .A2(new_n627), .ZN(new_n777));
  INV_X1    g0577(.A(new_n626), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n652), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT100), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n652), .B1(new_n518), .B2(new_n520), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n539), .A2(new_n542), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT99), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n539), .A2(new_n785), .A3(new_n542), .A4(new_n782), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n532), .A2(new_n535), .A3(new_n538), .A4(new_n652), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n781), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n783), .A2(KEYINPUT99), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n790), .A2(KEYINPUT100), .A3(new_n787), .A4(new_n786), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n780), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n789), .A2(new_n791), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n699), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n775), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT101), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n689), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n798), .A3(new_n689), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n707), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n794), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n748), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n736), .A2(G143), .B1(G159), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n725), .A2(G150), .B1(new_n754), .B2(G137), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT34), .Z(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n258), .B1(new_n743), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT98), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n740), .A2(G68), .B1(new_n734), .B2(G50), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n728), .A2(G58), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n737), .A2(new_n818), .B1(new_n294), .B2(new_n727), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G107), .A2(new_n734), .B1(new_n752), .B2(G311), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n760), .B2(new_n747), .ZN(new_n822));
  INV_X1    g0622(.A(new_n725), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n823), .A2(new_n758), .B1(new_n748), .B2(new_n711), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n263), .B1(new_n739), .B2(new_n213), .ZN(new_n825));
  OR3_X1    g0625(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n809), .A2(new_n817), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n718), .A2(new_n803), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n827), .A2(new_n718), .B1(new_n217), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n708), .B1(new_n804), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(KEYINPUT102), .B1(new_n802), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n799), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n796), .B2(new_n775), .ZN(new_n833));
  INV_X1    g0633(.A(new_n801), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n708), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT102), .ZN(new_n836));
  INV_X1    g0636(.A(new_n830), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n831), .A2(new_n838), .ZN(G384));
  OR2_X1    g0639(.A1(new_n368), .A2(KEYINPUT35), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n368), .A2(KEYINPUT35), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n840), .A2(G116), .A3(new_n230), .A4(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT36), .Z(new_n843));
  OR3_X1    g0643(.A1(new_n549), .A2(new_n227), .A3(new_n217), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n206), .B(G13), .C1(new_n844), .C2(new_n247), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT39), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT37), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n589), .A2(KEYINPUT16), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n546), .B1(new_n558), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n578), .B2(new_n643), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n848), .B1(new_n851), .B2(new_n592), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT103), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n561), .A2(new_n562), .A3(new_n643), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT104), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n561), .A2(KEYINPUT104), .A3(new_n562), .A4(new_n643), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n579), .A2(new_n848), .A3(new_n592), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n859), .A2(KEYINPUT105), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT105), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n854), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n850), .A2(new_n643), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n595), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n565), .A2(new_n575), .A3(G190), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n582), .B2(new_n506), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT106), .B1(new_n868), .B2(new_n559), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT106), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n583), .A2(new_n591), .A3(new_n870), .ZN(new_n871));
  AND4_X1   g0671(.A1(new_n611), .A2(new_n609), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n861), .B2(new_n862), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n593), .A2(new_n614), .A3(new_n615), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n857), .A3(new_n858), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n847), .B1(new_n866), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n852), .B(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n859), .A2(new_n860), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT105), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n865), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n880), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n488), .A2(new_n502), .A3(new_n644), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n879), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n616), .A2(new_n643), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n502), .A2(new_n652), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n503), .A2(new_n510), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n502), .B(new_n652), .C1(new_n509), .C2(new_n488), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n539), .A2(new_n652), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n793), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n888), .A2(new_n889), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n894), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n893), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n700), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n698), .B(new_n622), .C1(new_n780), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n621), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT107), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n905), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT108), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n866), .B2(new_n878), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n859), .B1(new_n616), .B2(new_n593), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n884), .A2(new_n885), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n874), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n889), .B(KEYINPUT108), .C1(new_n916), .C2(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n686), .A2(new_n687), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n386), .A2(new_n390), .A3(new_n425), .ZN(new_n919));
  NOR4_X1   g0719(.A1(new_n919), .A2(new_n306), .A3(new_n345), .A4(new_n652), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n898), .B(new_n792), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n913), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n921), .B1(new_n888), .B2(new_n889), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(KEYINPUT40), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n688), .A2(new_n622), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  INV_X1    g0729(.A(G330), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n911), .A2(new_n931), .B1(new_n206), .B2(new_n704), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n911), .A2(new_n931), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n846), .B1(new_n932), .B2(new_n933), .ZN(G367));
  NAND2_X1  g0734(.A1(new_n385), .A2(new_n652), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n386), .A2(new_n390), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n631), .A2(new_n633), .A3(new_n385), .A4(new_n652), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(KEYINPUT111), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(KEYINPUT111), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n660), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT42), .Z(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n938), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n386), .B1(new_n942), .B2(new_n337), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n644), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n644), .B1(new_n411), .B2(new_n412), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT109), .ZN(new_n947));
  INV_X1    g0747(.A(new_n423), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT110), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n949), .B(KEYINPUT110), .C1(new_n424), .C2(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n945), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n941), .A2(new_n953), .A3(new_n944), .A4(new_n952), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n658), .A2(new_n942), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n664), .B(KEYINPUT41), .Z(new_n962));
  NAND3_X1  g0762(.A1(new_n661), .A2(new_n938), .A3(new_n939), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT45), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n661), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n968), .A2(new_n942), .A3(KEYINPUT44), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT44), .B1(new_n968), .B2(new_n942), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n967), .A2(new_n971), .A3(new_n658), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n965), .A2(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  INV_X1    g0773(.A(new_n658), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n657), .B(new_n659), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n650), .B(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n975), .A3(new_n702), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n962), .B1(new_n978), .B2(new_n702), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n961), .B1(new_n979), .B2(new_n706), .ZN(new_n980));
  INV_X1    g0780(.A(new_n714), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n720), .B1(new_n232), .B2(new_n410), .C1(new_n981), .C2(new_n242), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n982), .A2(new_n707), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n739), .A2(new_n217), .B1(new_n733), .B2(new_n548), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n263), .B(new_n984), .C1(G159), .C2(new_n725), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n736), .A2(G150), .B1(G50), .B2(new_n805), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n754), .A2(G143), .B1(new_n752), .B2(G137), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n728), .A2(G68), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n823), .A2(new_n818), .B1(new_n748), .B2(new_n758), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G317), .B2(new_n752), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n728), .A2(G107), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n258), .B1(new_n754), .B2(G311), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n736), .A2(G303), .B1(G97), .B2(new_n740), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT112), .B1(new_n733), .B2(new_n711), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT46), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n989), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT47), .Z(new_n999));
  OAI221_X1 g0799(.A(new_n983), .B1(new_n722), .B2(new_n999), .C1(new_n955), .C2(new_n768), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n980), .A2(new_n1000), .ZN(G387));
  OR2_X1    g0801(.A1(new_n657), .A2(new_n768), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n714), .B1(new_n239), .B2(new_n433), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n710), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n666), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n445), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT50), .B1(new_n445), .B2(G50), .ZN(new_n1007));
  AOI21_X1  g0807(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n666), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1005), .A2(new_n1009), .B1(new_n219), .B2(new_n663), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n720), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n707), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n737), .A2(new_n202), .B1(new_n748), .B2(new_n211), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n446), .B2(new_n725), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n728), .A2(new_n417), .ZN(new_n1015));
  INV_X1    g0815(.A(G150), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n733), .A2(new_n217), .B1(new_n743), .B2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n263), .B(new_n1017), .C1(G97), .C2(new_n740), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n754), .A2(G159), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT113), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n258), .B1(new_n752), .B2(G326), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n736), .A2(G317), .B1(G303), .B2(new_n805), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n725), .A2(G311), .B1(new_n754), .B2(G322), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT114), .Z(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n728), .A2(G283), .B1(new_n734), .B2(G294), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1022), .B1(new_n711), .B2(new_n739), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1021), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1012), .B1(new_n1035), .B2(new_n718), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n977), .A2(new_n706), .B1(new_n1002), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n977), .A2(new_n702), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(KEYINPUT115), .A3(new_n664), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n702), .B2(new_n977), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT115), .B1(new_n1038), .B2(new_n664), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT116), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(KEYINPUT116), .B(new_n1037), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(G393));
  INV_X1    g0846(.A(new_n975), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n973), .A2(new_n974), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n705), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n942), .A2(new_n719), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n720), .B1(new_n294), .B2(new_n232), .C1(new_n981), .C2(new_n246), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n707), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n736), .A2(G159), .B1(new_n754), .B2(G150), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  AOI22_X1  g0854(.A1(new_n446), .A2(new_n805), .B1(new_n734), .B2(G68), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n725), .A2(G50), .B1(G143), .B2(new_n752), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n727), .A2(new_n217), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n263), .B(new_n1057), .C1(G87), .C2(new_n740), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n736), .A2(G311), .B1(new_n754), .B2(G317), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT52), .Z(new_n1061));
  AOI22_X1  g0861(.A1(new_n725), .A2(G303), .B1(G294), .B2(new_n805), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n711), .C2(new_n727), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G283), .A2(new_n734), .B1(new_n752), .B2(G322), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(new_n263), .A3(new_n741), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT117), .Z(new_n1066));
  OAI21_X1  g0866(.A(new_n1059), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1052), .B1(new_n1067), .B2(new_n718), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1049), .B1(new_n1050), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1038), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n664), .A3(new_n978), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(G390));
  NAND4_X1  g0872(.A1(new_n688), .A2(G330), .A3(new_n792), .A4(new_n898), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n697), .A2(new_n792), .A3(new_n644), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n901), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n892), .B1(new_n1076), .B2(new_n898), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n913), .A2(new_n1077), .A3(new_n917), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n901), .B1(new_n699), .B2(new_n794), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n892), .B1(new_n1079), .B2(new_n898), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n879), .B2(new_n890), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1074), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1080), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n890), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n875), .A2(new_n877), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n880), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n1086), .B2(new_n889), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n913), .A2(new_n1077), .A3(new_n917), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n1089), .A3(new_n1073), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n803), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n828), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n707), .B1(new_n446), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n733), .A2(new_n1016), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n736), .A2(G132), .B1(G125), .B2(new_n752), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT54), .B(G143), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1097), .B(new_n1098), .C1(new_n748), .C2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n725), .A2(G137), .B1(new_n754), .B2(G128), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n263), .B1(new_n740), .B2(G50), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n744), .C2(new_n727), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n725), .A2(G107), .B1(G97), .B2(new_n805), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n711), .B2(new_n737), .C1(new_n818), .C2(new_n743), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n754), .A2(G283), .B1(new_n740), .B2(G68), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1057), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1106), .A2(new_n263), .A3(new_n735), .A4(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1100), .A2(new_n1103), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1095), .B1(new_n1109), .B2(new_n718), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1092), .A2(new_n706), .B1(new_n1093), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n688), .A2(new_n622), .A3(G330), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n907), .A2(new_n621), .A3(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(G330), .B(new_n792), .C1(new_n918), .C2(new_n920), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n899), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n1073), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1079), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1115), .A2(new_n1073), .A3(new_n901), .A4(new_n1075), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1082), .A2(new_n1090), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT118), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n664), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1119), .A2(KEYINPUT119), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT119), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1124), .B(new_n1113), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1091), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1121), .B1(new_n1120), .B2(new_n664), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1111), .B1(new_n1128), .B2(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(new_n1113), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1120), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT57), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n921), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT38), .B1(new_n863), .B2(new_n865), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n866), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n930), .B1(new_n1136), .B2(new_n922), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n602), .A2(new_n513), .A3(new_n604), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n512), .A2(new_n643), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n602), .A2(new_n604), .A3(new_n513), .A4(new_n1139), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1137), .A2(new_n924), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1137), .B2(new_n924), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1147), .A2(new_n1148), .A3(new_n905), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n893), .A2(new_n904), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n913), .A2(new_n917), .A3(new_n923), .ZN(new_n1152));
  OAI21_X1  g0952(.A(G330), .B1(new_n925), .B2(KEYINPUT40), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1137), .A2(new_n924), .A3(new_n1146), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT120), .B1(new_n1149), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n905), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1133), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1154), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1158), .A2(new_n1162), .B1(new_n1120), .B2(new_n1131), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n664), .B1(new_n1163), .B2(KEYINPUT57), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1146), .A2(new_n803), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n707), .B1(G50), .B2(new_n1094), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n733), .A2(new_n1099), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G128), .A2(new_n736), .B1(new_n725), .B2(G132), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G125), .A2(new_n754), .B1(new_n805), .B2(G137), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n728), .A2(G150), .ZN(new_n1172));
  AND4_X1   g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT59), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n255), .B(new_n432), .C1(new_n739), .C2(new_n744), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G124), .B2(new_n752), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n417), .A2(new_n805), .B1(new_n752), .B2(G283), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n263), .A2(new_n432), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G77), .B2(new_n734), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1182), .A3(new_n988), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n737), .A2(new_n219), .B1(new_n548), .B2(new_n739), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n823), .A2(new_n294), .B1(new_n747), .B2(new_n711), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT58), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1181), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1186), .A2(KEYINPUT58), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1179), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1168), .B1(new_n1190), .B2(new_n718), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1166), .A2(new_n706), .B1(new_n1167), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1165), .A2(new_n1192), .ZN(G375));
  INV_X1    g0993(.A(new_n962), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1126), .B(new_n1194), .C1(new_n1131), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n706), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n707), .B1(G68), .B2(new_n1094), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n736), .A2(G137), .B1(G159), .B2(new_n734), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n1016), .B2(new_n748), .C1(new_n823), .C2(new_n1099), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n754), .A2(G132), .B1(new_n752), .B2(G128), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n263), .B1(new_n740), .B2(G58), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n202), .C2(new_n727), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G116), .A2(new_n725), .B1(new_n736), .B2(G283), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G294), .A2(new_n754), .B1(new_n805), .B2(G107), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n258), .B1(new_n740), .B2(G77), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1204), .A2(new_n1015), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n733), .A2(new_n294), .B1(new_n743), .B2(new_n760), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT121), .Z(new_n1209));
  OAI22_X1  g1009(.A1(new_n1200), .A2(new_n1203), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1198), .B1(new_n1210), .B2(new_n718), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n803), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n898), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1197), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1196), .A2(new_n1215), .ZN(G381));
  INV_X1    g1016(.A(G375), .ZN(new_n1217));
  INV_X1    g1017(.A(G378), .ZN(new_n1218));
  INV_X1    g1018(.A(G390), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n831), .A2(new_n838), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1044), .A2(new_n773), .A3(new_n1045), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1221), .A2(G387), .A3(new_n1222), .A4(G381), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1217), .A2(new_n1218), .A3(new_n1223), .ZN(G407));
  INV_X1    g1024(.A(G213), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(G343), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1217), .A2(new_n1218), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(G407), .A2(new_n1227), .A3(G213), .ZN(G409));
  OAI211_X1 g1028(.A(G378), .B(new_n1192), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1129), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1127), .A3(new_n1122), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1166), .A2(new_n1132), .A3(new_n1194), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1167), .A2(new_n1191), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n705), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1231), .B(new_n1111), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1229), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1226), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1119), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n664), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT122), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1195), .B2(new_n1131), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1241), .B(KEYINPUT60), .C1(new_n1195), .C2(new_n1131), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1240), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(G384), .A3(new_n1215), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1220), .B1(new_n1246), .B2(new_n1214), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1237), .A2(new_n1238), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1226), .B1(new_n1229), .B2(new_n1236), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1251), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1219), .A2(G387), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(G390), .A2(new_n980), .A3(new_n1000), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G393), .A2(G396), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1222), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1257), .A2(new_n1260), .A3(new_n1222), .A4(new_n1258), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1254), .A2(new_n1256), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1226), .A2(KEYINPUT124), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1248), .A2(new_n1249), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1226), .A2(G2897), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1269), .B(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1255), .B2(KEYINPUT123), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT123), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1273), .B(new_n1226), .C1(new_n1229), .C2(new_n1236), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT125), .B1(new_n1267), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1273), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1255), .A2(KEYINPUT123), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1271), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1265), .B1(new_n1253), .B2(new_n1252), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .A4(new_n1256), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1276), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1277), .B2(new_n1271), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1252), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1252), .B2(new_n1286), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1285), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1284), .A2(new_n1292), .ZN(G405));
  NAND3_X1  g1093(.A1(new_n1262), .A2(new_n1251), .A3(new_n1264), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1251), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT127), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1250), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1294), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1218), .ZN(new_n1301));
  AND4_X1   g1101(.A1(new_n1229), .A2(new_n1297), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1297), .A2(new_n1300), .B1(new_n1229), .B2(new_n1301), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(G402));
endmodule


