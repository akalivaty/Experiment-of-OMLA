//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  OAI21_X1  g005(.A(G214), .B1(G237), .B2(G902), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n197), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G116), .ZN(new_n205));
  INV_X1    g019(.A(G116), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  INV_X1    g021(.A(G113), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n205), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(new_n207), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT2), .B(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n199), .A2(new_n216), .A3(G101), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n203), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n206), .A2(G119), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n221), .B(new_n222), .C1(new_n212), .C2(new_n219), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT5), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT86), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT86), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n220), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(G113), .C1(new_n212), .C2(new_n219), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT87), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n223), .A2(new_n230), .A3(new_n211), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n196), .A2(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n193), .A2(G107), .ZN(new_n233));
  OAI21_X1  g047(.A(G101), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n202), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT81), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n202), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n218), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n241), .B(new_n218), .C1(new_n231), .C2(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(KEYINPUT6), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT6), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n246), .A3(new_n242), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(KEYINPUT1), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n249), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n252), .B(G146), .C1(new_n248), .C2(KEYINPUT1), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n250), .A3(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G125), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n251), .A2(new_n253), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G143), .B(G146), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT0), .B(G128), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G125), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G224), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G953), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n245), .A2(new_n247), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(G210), .B1(G237), .B2(G902), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT88), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n265), .B2(G125), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT7), .B1(new_n268), .B2(G953), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n267), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n260), .A2(new_n273), .A3(new_n266), .A4(new_n275), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n241), .B(KEYINPUT8), .Z(new_n279));
  OAI21_X1  g093(.A(new_n221), .B1(new_n224), .B2(new_n212), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n211), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n202), .A2(new_n234), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n223), .A2(new_n230), .A3(new_n211), .A4(new_n235), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n277), .A2(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n285), .B2(new_n244), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n271), .A2(new_n272), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n272), .B(KEYINPUT89), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n271), .B2(new_n286), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n192), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G953), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G227), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(KEYINPUT79), .ZN(new_n295));
  XNOR2_X1  g109(.A(G110), .B(G140), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n199), .A2(G101), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n265), .B1(new_n299), .B2(new_n216), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n249), .A2(new_n251), .A3(new_n253), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT80), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n255), .A2(new_n256), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n263), .A2(new_n304), .A3(new_n249), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n282), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n203), .A2(new_n300), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT66), .B1(new_n254), .B2(new_n257), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n301), .A2(new_n311), .A3(new_n255), .A4(new_n256), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n202), .A2(new_n234), .A3(new_n237), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n237), .B1(new_n202), .B2(new_n234), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT11), .B1(new_n318), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT11), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G134), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT64), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n321), .B2(G134), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(KEYINPUT64), .A3(G137), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G131), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n319), .A2(new_n322), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n325), .A4(new_n326), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n309), .A2(new_n317), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n331), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n318), .A2(KEYINPUT64), .A3(G137), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT64), .B1(new_n318), .B2(G137), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n330), .B1(new_n336), .B2(new_n329), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT82), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n328), .A2(new_n339), .A3(new_n331), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n265), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n342), .B(new_n217), .C1(new_n299), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n307), .A2(new_n308), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n317), .A2(new_n341), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT83), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n309), .A2(new_n348), .A3(new_n317), .A4(new_n341), .ZN(new_n349));
  AOI211_X1 g163(.A(new_n298), .B(new_n332), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n258), .A2(new_n235), .ZN(new_n352));
  AOI221_X4 g166(.A(new_n351), .B1(new_n328), .B2(new_n331), .C1(new_n307), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n307), .A2(new_n352), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n328), .A2(new_n331), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT12), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n347), .B2(new_n349), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n297), .B1(new_n358), .B2(KEYINPUT84), .ZN(new_n359));
  INV_X1    g173(.A(new_n357), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n257), .B1(KEYINPUT80), .B2(new_n301), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n235), .B1(new_n361), .B2(new_n305), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n344), .B1(new_n362), .B2(KEYINPUT10), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n312), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n239), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n348), .B1(new_n366), .B2(new_n341), .ZN(new_n367));
  INV_X1    g181(.A(new_n349), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n360), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n350), .B1(new_n359), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G469), .B1(new_n372), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n332), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n367), .B2(new_n368), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n298), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n332), .B1(new_n347), .B2(new_n349), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT85), .B1(new_n378), .B2(new_n297), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n298), .B1(new_n347), .B2(new_n349), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n360), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n190), .ZN(new_n384));
  AOI211_X1 g198(.A(new_n191), .B(new_n292), .C1(new_n373), .C2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G472), .A2(G902), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n318), .A2(G137), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n321), .A2(G134), .ZN(new_n388));
  OAI21_X1  g202(.A(G131), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n331), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT65), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n258), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n331), .A2(KEYINPUT65), .A3(new_n389), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n342), .B1(new_n333), .B2(new_n337), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT30), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n310), .A2(new_n331), .A3(new_n312), .A4(new_n389), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n215), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n211), .A2(new_n214), .A3(KEYINPUT67), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT67), .B1(new_n211), .B2(new_n214), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n396), .A3(new_n398), .ZN(new_n405));
  NOR2_X1   g219(.A1(G237), .A2(G953), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G210), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT27), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G101), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT68), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n265), .B1(new_n328), .B2(new_n331), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n258), .B1(new_n390), .B2(new_n391), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(new_n394), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n215), .B(new_n399), .C1(new_n415), .C2(KEYINPUT30), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n410), .A4(new_n405), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n412), .A2(KEYINPUT31), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n400), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n331), .A2(KEYINPUT65), .A3(new_n389), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT65), .B1(new_n331), .B2(new_n389), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n422), .A2(new_n423), .A3(new_n258), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n421), .B1(new_n424), .B2(new_n413), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n411), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT31), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n405), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n215), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n405), .B1(new_n415), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n428), .B1(new_n435), .B2(new_n410), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n386), .B1(new_n419), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n405), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n404), .A2(new_n396), .A3(KEYINPUT72), .A4(new_n398), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n396), .A2(new_n398), .ZN(new_n445));
  INV_X1    g259(.A(new_n404), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT73), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT73), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n431), .B1(new_n451), .B2(KEYINPUT28), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n410), .A2(KEYINPUT29), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n432), .B1(new_n395), .B2(new_n396), .ZN(new_n455));
  INV_X1    g269(.A(new_n405), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n434), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n410), .A3(new_n430), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT71), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n435), .A2(new_n460), .A3(new_n410), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n416), .A2(new_n405), .ZN(new_n462));
  INV_X1    g276(.A(new_n410), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT29), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G472), .ZN(new_n467));
  INV_X1    g281(.A(new_n386), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n457), .A2(new_n430), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n469), .A2(new_n463), .B1(new_n426), .B2(new_n427), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n412), .A2(KEYINPUT31), .A3(new_n418), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT70), .B1(new_n472), .B2(KEYINPUT32), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n440), .A2(new_n467), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G234), .ZN(new_n476));
  OAI21_X1  g290(.A(G217), .B1(new_n476), .B2(G902), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT74), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n204), .B2(G128), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n204), .A2(G128), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n484), .A2(KEYINPUT76), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(KEYINPUT76), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(G110), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(KEYINPUT77), .A2(G125), .ZN(new_n488));
  INV_X1    g302(.A(G140), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(KEYINPUT77), .A2(G125), .A3(G140), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT16), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n259), .B2(G140), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G146), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n250), .A3(new_n494), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT24), .B(G110), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT75), .B1(new_n204), .B2(G128), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT75), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n248), .A3(G119), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n502), .A3(new_n483), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n487), .B(new_n498), .C1(new_n499), .C2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G125), .B(G140), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n505), .A2(new_n250), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n495), .B2(G146), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n503), .A2(new_n499), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(G110), .B2(new_n484), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n507), .A2(KEYINPUT78), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT78), .B1(new_n507), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n187), .A2(new_n476), .A3(G953), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n513), .B(new_n514), .Z(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n504), .B(new_n515), .C1(new_n510), .C2(new_n511), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n190), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT25), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(KEYINPUT25), .A3(new_n190), .A4(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n479), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n518), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n478), .A2(G902), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n193), .ZN(new_n529));
  INV_X1    g343(.A(G237), .ZN(new_n530));
  AND4_X1   g344(.A1(G143), .A2(new_n530), .A3(new_n293), .A4(G214), .ZN(new_n531));
  AOI21_X1  g345(.A(G143), .B1(new_n406), .B2(G214), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT18), .B(G131), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n293), .A3(G214), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n252), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n406), .A2(G143), .A3(G214), .ZN(new_n536));
  NAND2_X1  g350(.A1(KEYINPUT18), .A2(G131), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n490), .A2(new_n491), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(new_n250), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n533), .B(new_n538), .C1(new_n506), .C2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT17), .B(G131), .C1(new_n531), .C2(new_n532), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n496), .A2(new_n497), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G131), .B1(new_n531), .B2(new_n532), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n535), .A2(new_n330), .A3(new_n536), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n529), .B(new_n541), .C1(new_n543), .C2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n551), .A2(new_n496), .A3(new_n497), .A4(new_n542), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n552), .A2(KEYINPUT90), .A3(new_n529), .A4(new_n541), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n552), .A2(new_n541), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n529), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n190), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT20), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT91), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n544), .A2(new_n546), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT19), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n505), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n562), .B2(new_n539), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n561), .B(new_n496), .C1(G146), .C2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n529), .B1(new_n565), .B2(new_n541), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n560), .B1(new_n554), .B2(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(KEYINPUT91), .B(new_n566), .C1(new_n550), .C2(new_n553), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G475), .A2(G902), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n559), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  AOI211_X1 g387(.A(KEYINPUT20), .B(new_n573), .C1(new_n554), .C2(new_n567), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n558), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G952), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(G953), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n476), .B2(new_n530), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT21), .B(G898), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT96), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n190), .B(new_n293), .C1(G234), .C2(G237), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n585), .A2(new_n586), .B1(new_n248), .B2(G143), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n585), .B2(new_n586), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G134), .ZN(new_n589));
  XNOR2_X1  g403(.A(G128), .B(G143), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(G134), .A3(new_n590), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n206), .A2(G122), .ZN(new_n595));
  INV_X1    g409(.A(G122), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n596), .A2(KEYINPUT92), .A3(G116), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT92), .B1(new_n596), .B2(G116), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G107), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n196), .B(new_n595), .C1(new_n597), .C2(new_n598), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n591), .A2(new_n318), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n590), .A2(G134), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n595), .A2(KEYINPUT14), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT14), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n206), .A3(G122), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n608), .B(new_n610), .C1(new_n597), .C2(new_n598), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(KEYINPUT94), .A3(G107), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT94), .B1(new_n611), .B2(G107), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n607), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n189), .A2(G217), .A3(new_n293), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n603), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT95), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n603), .A2(new_n615), .A3(new_n620), .A4(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n603), .A2(new_n615), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n616), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n619), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n190), .ZN(new_n625));
  INV_X1    g439(.A(G478), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(KEYINPUT15), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n624), .B(new_n190), .C1(KEYINPUT15), .C2(new_n626), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n575), .A2(new_n584), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n385), .A2(new_n475), .A3(new_n527), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NAND2_X1  g447(.A1(new_n625), .A2(new_n626), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n624), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n635), .B1(new_n637), .B2(new_n617), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n622), .A2(KEYINPUT97), .A3(new_n616), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n626), .A2(G902), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n634), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n575), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n192), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n271), .A2(new_n286), .ZN(new_n647));
  INV_X1    g461(.A(new_n272), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n649), .B2(new_n287), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n645), .A2(new_n584), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n191), .B1(new_n373), .B2(new_n384), .ZN(new_n653));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  AOI21_X1  g468(.A(G902), .B1(new_n470), .B2(new_n471), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n437), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n527), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n652), .A2(new_n653), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  NOR4_X1   g476(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT20), .A4(new_n573), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n558), .B(new_n630), .C1(new_n572), .C2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n664), .B2(new_n584), .ZN(new_n665));
  INV_X1    g479(.A(new_n558), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n554), .A2(new_n567), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT91), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n554), .A2(new_n560), .A3(new_n567), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n571), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT20), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n570), .A2(new_n559), .A3(new_n571), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n666), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n584), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n673), .A2(KEYINPUT98), .A3(new_n674), .A4(new_n630), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n665), .A2(new_n650), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n653), .A3(new_n658), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NAND2_X1  g493(.A1(new_n521), .A2(new_n522), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n478), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n516), .A2(KEYINPUT36), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n512), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n512), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n685), .A2(G902), .A3(new_n478), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT99), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n681), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT99), .B1(new_n523), .B2(new_n686), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n656), .ZN(new_n692));
  INV_X1    g506(.A(new_n292), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n653), .A3(new_n631), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  AOI21_X1  g510(.A(new_n438), .B1(new_n437), .B2(new_n439), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n472), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n466), .A2(G472), .B1(new_n472), .B2(KEYINPUT32), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n691), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n653), .A2(new_n650), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n579), .B1(new_n583), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n664), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n248), .ZN(G30));
  XOR2_X1   g523(.A(new_n705), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n653), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n451), .A2(new_n463), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n412), .A2(new_n418), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n190), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G472), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n699), .A2(new_n474), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n291), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n287), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT38), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n575), .A2(new_n630), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n523), .A2(new_n686), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n646), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n721), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n712), .A2(new_n713), .A3(new_n718), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  INV_X1    g543(.A(new_n705), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n574), .B1(new_n670), .B2(KEYINPUT20), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n644), .B(new_n730), .C1(new_n731), .C2(new_n666), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n575), .A2(KEYINPUT100), .A3(new_n644), .A4(new_n730), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n703), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n250), .ZN(G48));
  NAND2_X1  g552(.A1(new_n382), .A2(new_n190), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G469), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(KEYINPUT101), .A3(new_n384), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT101), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n742), .A3(G469), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n191), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n657), .B1(new_n699), .B2(new_n700), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n652), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT102), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n747), .B(new_n749), .ZN(G15));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n676), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G116), .ZN(G18));
  NAND4_X1  g566(.A1(new_n744), .A2(new_n701), .A3(new_n631), .A4(new_n650), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  NAND2_X1  g568(.A1(new_n470), .A2(new_n471), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n654), .B1(new_n755), .B2(new_n190), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n471), .B(new_n428), .C1(new_n452), .C2(new_n410), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n386), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n759), .A3(new_n527), .A4(new_n674), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n575), .A2(new_n630), .A3(new_n650), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n744), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  AND2_X1   g578(.A1(new_n734), .A2(new_n735), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n757), .A2(new_n759), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n724), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n744), .A2(new_n650), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  NOR2_X1   g583(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n700), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n527), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n719), .A2(new_n192), .A3(new_n287), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n191), .B(new_n775), .C1(new_n373), .C2(new_n384), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT42), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n774), .A2(new_n777), .A3(new_n736), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  INV_X1    g593(.A(new_n775), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n475), .A2(new_n653), .A3(new_n527), .A4(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n779), .B1(new_n781), .B2(new_n736), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT103), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT103), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n779), .C1(new_n781), .C2(new_n736), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n778), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n330), .ZN(G33));
  NOR2_X1   g601(.A1(new_n781), .A2(new_n707), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n318), .ZN(G36));
  INV_X1    g603(.A(new_n644), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n575), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT105), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT43), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n795), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n656), .A3(new_n725), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT44), .Z(new_n799));
  INV_X1    g613(.A(new_n191), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n359), .A2(new_n371), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n350), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n372), .A2(KEYINPUT45), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(G469), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(G469), .A2(G902), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT46), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n384), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n800), .B(new_n710), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n775), .B(KEYINPUT106), .Z(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n799), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n321), .ZN(G39));
  OAI21_X1  g630(.A(new_n800), .B1(new_n810), .B2(new_n811), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n736), .A2(new_n475), .A3(new_n527), .A4(new_n775), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(new_n489), .ZN(G42));
  AND2_X1   g636(.A1(new_n797), .A2(new_n579), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n766), .A2(new_n657), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT115), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n721), .A2(new_n192), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n826), .A2(new_n744), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n744), .A2(new_n829), .ZN(new_n831));
  OAI211_X1 g645(.A(KEYINPUT115), .B(new_n827), .C1(new_n825), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n744), .A2(new_n780), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n823), .A2(new_n767), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n718), .A2(new_n657), .A3(new_n578), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n731), .A2(new_n666), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n834), .A2(new_n836), .A3(new_n837), .A4(new_n790), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n833), .A2(KEYINPUT51), .A3(new_n835), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n741), .A2(new_n743), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n800), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n819), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(KEYINPUT116), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n826), .A2(new_n813), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n843), .B2(KEYINPUT116), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n839), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n833), .A2(new_n835), .A3(new_n838), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(new_n813), .A3(new_n826), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT51), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n823), .A2(new_n834), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n774), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT48), .Z(new_n853));
  NAND4_X1  g667(.A1(new_n834), .A2(new_n836), .A3(new_n575), .A4(new_n644), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n826), .A2(new_n650), .A3(new_n744), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n577), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n847), .A2(new_n850), .A3(new_n856), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n774), .A2(new_n777), .A3(new_n736), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n745), .A2(new_n765), .A3(new_n776), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n784), .B1(new_n859), .B2(new_n779), .ZN(new_n860));
  INV_X1    g674(.A(new_n785), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n745), .B(new_n744), .C1(new_n676), .C2(new_n652), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n753), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n575), .A2(KEYINPUT107), .A3(new_n644), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT107), .B1(new_n575), .B2(new_n644), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n674), .B(new_n192), .C1(new_n288), .C2(new_n291), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n867), .A2(new_n653), .A3(new_n658), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n763), .A2(new_n870), .A3(new_n632), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n837), .A3(KEYINPUT108), .A4(new_n630), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT108), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n558), .B(new_n630), .C1(new_n572), .C2(new_n574), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n875), .B2(new_n868), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n873), .A2(new_n658), .A3(new_n653), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n694), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT109), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n694), .A3(KEYINPUT109), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n653), .A2(new_n780), .ZN(new_n883));
  INV_X1    g697(.A(new_n630), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n673), .A2(new_n884), .A3(new_n730), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n691), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n475), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n756), .B1(new_n386), .B2(new_n758), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n734), .A2(new_n889), .A3(new_n735), .A4(new_n725), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n883), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n788), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n862), .A2(new_n872), .A3(new_n882), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT110), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n891), .A2(new_n788), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n783), .A2(new_n785), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n896), .B2(new_n858), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n877), .A2(new_n694), .A3(KEYINPUT109), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT109), .B1(new_n877), .B2(new_n694), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n900), .A2(new_n864), .A3(new_n871), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT110), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT111), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT53), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n701), .B(new_n702), .C1(new_n765), .C2(new_n706), .ZN(new_n907));
  INV_X1    g721(.A(new_n761), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n725), .A2(new_n705), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n718), .A2(new_n653), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n768), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT113), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT112), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT52), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(KEYINPUT112), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT52), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT112), .B1(new_n911), .B2(new_n912), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT114), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT114), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n916), .B(new_n922), .C1(new_n918), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n894), .A2(KEYINPUT111), .A3(new_n903), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n906), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n911), .B(new_n915), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n763), .A2(new_n870), .A3(new_n632), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n882), .A2(new_n928), .A3(new_n753), .A4(new_n863), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n929), .A2(new_n786), .A3(KEYINPUT110), .A4(new_n895), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n902), .B1(new_n897), .B2(new_n901), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT53), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n926), .A2(KEYINPUT54), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT53), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n897), .A2(new_n901), .A3(KEYINPUT53), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n923), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n913), .A2(new_n914), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n915), .B1(new_n911), .B2(KEYINPUT112), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n922), .B1(new_n942), .B2(new_n916), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT54), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n936), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n857), .A2(new_n934), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT117), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT117), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n857), .A2(new_n934), .A3(new_n949), .A4(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n576), .A2(new_n293), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n841), .A2(KEYINPUT49), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n527), .A2(new_n800), .A3(new_n192), .ZN(new_n954));
  NOR4_X1   g768(.A1(new_n718), .A2(new_n721), .A3(new_n792), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n841), .A2(KEYINPUT49), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n952), .A2(new_n957), .ZN(G75));
  NOR2_X1   g772(.A1(new_n293), .A2(G952), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT53), .B1(new_n904), .B2(new_n927), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n937), .B1(new_n921), .B2(new_n923), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n963), .A2(new_n190), .A3(new_n290), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n245), .A2(new_n247), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(new_n270), .Z(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT55), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(KEYINPUT56), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n960), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n963), .A2(new_n190), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(G210), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT118), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT56), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT118), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n970), .A2(new_n974), .A3(G210), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n969), .B1(new_n976), .B2(new_n967), .ZN(G51));
  INV_X1    g791(.A(KEYINPUT119), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n963), .A2(new_n190), .A3(new_n805), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n806), .B(KEYINPUT57), .Z(new_n980));
  NOR3_X1   g794(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT54), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n945), .B1(new_n936), .B2(new_n944), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n979), .B1(new_n983), .B2(new_n382), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n984), .B2(new_n959), .ZN(new_n985));
  INV_X1    g799(.A(new_n382), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT54), .B1(new_n961), .B2(new_n962), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n946), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(new_n980), .ZN(new_n989));
  OAI211_X1 g803(.A(KEYINPUT119), .B(new_n960), .C1(new_n989), .C2(new_n979), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n985), .A2(new_n990), .ZN(G54));
  NAND2_X1  g805(.A1(KEYINPUT58), .A2(G475), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT120), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n970), .A2(new_n570), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n570), .B1(new_n970), .B2(new_n993), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n994), .A2(new_n995), .A3(new_n959), .ZN(G60));
  NAND2_X1  g810(.A1(G478), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT59), .Z(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n934), .B2(new_n946), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n636), .B2(new_n640), .ZN(new_n1000));
  INV_X1    g814(.A(new_n988), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n641), .A2(new_n998), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n960), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1000), .A2(new_n1003), .ZN(G63));
  INV_X1    g818(.A(new_n685), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G217), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT60), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n1005), .B(new_n1008), .C1(new_n961), .C2(new_n962), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT121), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1009), .A2(new_n960), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n936), .A2(new_n944), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n525), .B1(new_n1015), .B2(new_n1008), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1014), .A2(new_n1016), .A3(KEYINPUT122), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT122), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1007), .B1(new_n936), .B2(new_n944), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n959), .B1(new_n1019), .B2(new_n1005), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n524), .B1(new_n963), .B2(new_n1007), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1013), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(KEYINPUT122), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1020), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1024), .A2(new_n1025), .A3(new_n1012), .A4(new_n1011), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1023), .A2(new_n1026), .ZN(G66));
  NOR2_X1   g841(.A1(new_n901), .A2(G953), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT123), .ZN(new_n1029));
  OAI21_X1  g843(.A(G953), .B1(new_n582), .B2(new_n268), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n965), .B1(G898), .B2(new_n293), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(G69));
  AOI21_X1  g847(.A(new_n293), .B1(G227), .B2(G900), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n425), .A2(new_n399), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT124), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1036), .B(KEYINPUT125), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(new_n564), .ZN(new_n1038));
  NAND2_X1  g852(.A1(G900), .A2(G953), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n815), .A2(new_n821), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n812), .A2(new_n761), .A3(new_n774), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n907), .A2(new_n768), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1041), .A2(new_n788), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1040), .A2(new_n862), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1038), .B(new_n1039), .C1(new_n1045), .C2(G953), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1034), .B1(new_n1046), .B2(KEYINPUT126), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n875), .B1(new_n865), .B2(new_n866), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n745), .A2(new_n1048), .A3(new_n710), .A4(new_n776), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1042), .A2(new_n728), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1050), .B(KEYINPUT62), .Z(new_n1051));
  NAND3_X1  g865(.A1(new_n1040), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n1052), .A2(new_n293), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1046), .B1(new_n1053), .B2(new_n1038), .ZN(new_n1054));
  XOR2_X1   g868(.A(new_n1047), .B(new_n1054), .Z(G72));
  NAND2_X1  g869(.A1(G472), .A2(G902), .ZN(new_n1056));
  XOR2_X1   g870(.A(new_n1056), .B(KEYINPUT63), .Z(new_n1057));
  OAI21_X1  g871(.A(new_n1057), .B1(new_n1052), .B2(new_n929), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1058), .A2(new_n410), .A3(new_n462), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1057), .B1(new_n1045), .B2(new_n929), .ZN(new_n1060));
  INV_X1    g874(.A(new_n462), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1060), .A2(new_n463), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n1059), .A2(new_n1062), .A3(new_n960), .ZN(new_n1063));
  AND2_X1   g877(.A1(new_n926), .A2(new_n933), .ZN(new_n1064));
  INV_X1    g878(.A(new_n1057), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n1061), .A2(KEYINPUT127), .A3(new_n410), .ZN(new_n1066));
  NOR2_X1   g880(.A1(new_n1066), .A2(new_n715), .ZN(new_n1067));
  OAI21_X1  g881(.A(KEYINPUT127), .B1(new_n1061), .B2(new_n410), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1063), .B1(new_n1064), .B2(new_n1069), .ZN(G57));
endmodule


