

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734;

  NOR2_X1 U361 ( .A1(n574), .A2(n573), .ZN(n582) );
  BUF_X1 U362 ( .A(G107), .Z(n341) );
  XNOR2_X2 U363 ( .A(n485), .B(n342), .ZN(n632) );
  XNOR2_X2 U364 ( .A(n486), .B(n347), .ZN(n342) );
  XNOR2_X2 U365 ( .A(n403), .B(n468), .ZN(n485) );
  INV_X1 U366 ( .A(G953), .ZN(n726) );
  XNOR2_X2 U367 ( .A(n477), .B(n476), .ZN(n669) );
  INV_X2 U368 ( .A(G128), .ZN(n388) );
  AND2_X2 U369 ( .A1(n528), .A2(n561), .ZN(n540) );
  NOR2_X1 U370 ( .A1(n652), .A2(n597), .ZN(n600) );
  XNOR2_X2 U371 ( .A(n402), .B(n410), .ZN(n486) );
  XNOR2_X2 U372 ( .A(G110), .B(G107), .ZN(n402) );
  XNOR2_X1 U373 ( .A(n559), .B(KEYINPUT107), .ZN(n624) );
  NOR2_X1 U374 ( .A1(n713), .A2(n680), .ZN(n583) );
  NAND2_X1 U375 ( .A1(n357), .A2(n659), .ZN(n372) );
  NOR2_X1 U376 ( .A1(n624), .A2(n560), .ZN(n352) );
  XNOR2_X1 U377 ( .A(n539), .B(n409), .ZN(n625) );
  NOR2_X1 U378 ( .A1(n365), .A2(n366), .ZN(n539) );
  NAND2_X1 U379 ( .A1(n525), .A2(n524), .ZN(n527) );
  AND2_X1 U380 ( .A1(n587), .A2(n567), .ZN(n568) );
  XNOR2_X1 U381 ( .A(n535), .B(n534), .ZN(n674) );
  NOR2_X1 U382 ( .A1(n573), .A2(n658), .ZN(n543) );
  AND2_X1 U383 ( .A1(n378), .A2(n377), .ZN(n376) );
  BUF_X1 U384 ( .A(n530), .Z(n659) );
  BUF_X1 U385 ( .A(n542), .Z(n573) );
  XNOR2_X1 U386 ( .A(n510), .B(KEYINPUT91), .ZN(n511) );
  XNOR2_X1 U387 ( .A(n475), .B(n474), .ZN(n618) );
  XOR2_X1 U388 ( .A(KEYINPUT59), .B(n606), .Z(n607) );
  XNOR2_X1 U389 ( .A(n469), .B(n467), .ZN(n403) );
  XNOR2_X1 U390 ( .A(n371), .B(G146), .ZN(n493) );
  XNOR2_X1 U391 ( .A(G116), .B(G113), .ZN(n468) );
  INV_X1 U392 ( .A(G119), .ZN(n467) );
  INV_X1 U393 ( .A(n603), .ZN(n343) );
  NAND2_X1 U394 ( .A1(n376), .A2(n373), .ZN(n581) );
  NOR2_X1 U395 ( .A1(n372), .A2(n556), .ZN(n557) );
  XNOR2_X1 U396 ( .A(n372), .B(n523), .ZN(n525) );
  BUF_X1 U397 ( .A(n486), .Z(n344) );
  XNOR2_X1 U398 ( .A(n500), .B(n499), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n500), .B(n499), .ZN(n506) );
  XNOR2_X2 U400 ( .A(G146), .B(n725), .ZN(n475) );
  XNOR2_X2 U401 ( .A(n423), .B(n408), .ZN(n725) );
  XNOR2_X1 U402 ( .A(n493), .B(n370), .ZN(n446) );
  INV_X1 U403 ( .A(KEYINPUT10), .ZN(n370) );
  XOR2_X1 U404 ( .A(G137), .B(G140), .Z(n447) );
  INV_X1 U405 ( .A(KEYINPUT45), .ZN(n396) );
  XNOR2_X1 U406 ( .A(n426), .B(n425), .ZN(n537) );
  XNOR2_X1 U407 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U408 ( .A(n380), .B(n592), .ZN(n596) );
  BUF_X1 U409 ( .A(n652), .Z(n626) );
  XNOR2_X1 U410 ( .A(n404), .B(n384), .ZN(n383) );
  XNOR2_X1 U411 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n384) );
  XNOR2_X1 U412 ( .A(n405), .B(KEYINPUT93), .ZN(n404) );
  INV_X1 U413 ( .A(G110), .ZN(n405) );
  XNOR2_X1 U414 ( .A(n443), .B(n442), .ZN(n382) );
  XNOR2_X1 U415 ( .A(G119), .B(G128), .ZN(n443) );
  XNOR2_X1 U416 ( .A(n387), .B(n385), .ZN(n419) );
  XNOR2_X1 U417 ( .A(KEYINPUT8), .B(KEYINPUT66), .ZN(n387) );
  NOR2_X1 U418 ( .A1(n386), .A2(G953), .ZN(n385) );
  XNOR2_X1 U419 ( .A(n422), .B(n392), .ZN(n391) );
  XNOR2_X1 U420 ( .A(n424), .B(n393), .ZN(n392) );
  INV_X1 U421 ( .A(n341), .ZN(n424) );
  XNOR2_X1 U422 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n488) );
  XNOR2_X1 U423 ( .A(KEYINPUT18), .B(KEYINPUT74), .ZN(n487) );
  INV_X1 U424 ( .A(G125), .ZN(n371) );
  NAND2_X1 U425 ( .A1(n364), .A2(n361), .ZN(n365) );
  AND2_X1 U426 ( .A1(n367), .A2(n368), .ZN(n364) );
  NAND2_X1 U427 ( .A1(n363), .A2(n362), .ZN(n361) );
  INV_X1 U428 ( .A(n589), .ZN(n368) );
  AND2_X1 U429 ( .A1(n674), .A2(n351), .ZN(n366) );
  INV_X1 U430 ( .A(KEYINPUT46), .ZN(n406) );
  XNOR2_X1 U431 ( .A(n418), .B(G469), .ZN(n542) );
  INV_X1 U432 ( .A(G234), .ZN(n386) );
  INV_X1 U433 ( .A(G116), .ZN(n393) );
  XNOR2_X1 U434 ( .A(n542), .B(KEYINPUT1), .ZN(n530) );
  NOR2_X1 U435 ( .A1(n369), .A2(n351), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n389), .B(KEYINPUT106), .ZN(n678) );
  NAND2_X1 U437 ( .A1(n537), .A2(n536), .ZN(n389) );
  INV_X1 U438 ( .A(KEYINPUT108), .ZN(n523) );
  XOR2_X1 U439 ( .A(G140), .B(G104), .Z(n428) );
  XNOR2_X1 U440 ( .A(G131), .B(G143), .ZN(n432) );
  INV_X1 U441 ( .A(G104), .ZN(n410) );
  XNOR2_X1 U442 ( .A(n447), .B(n411), .ZN(n412) );
  NAND2_X1 U443 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U444 ( .A1(n505), .A2(KEYINPUT19), .ZN(n374) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n444) );
  NAND2_X1 U446 ( .A1(n395), .A2(G217), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n632), .B(n358), .ZN(n613) );
  XNOR2_X1 U448 ( .A(n359), .B(n494), .ZN(n358) );
  NOR2_X1 U449 ( .A1(n726), .A2(G952), .ZN(n650) );
  XNOR2_X1 U450 ( .A(n654), .B(n355), .ZN(n354) );
  INV_X1 U451 ( .A(KEYINPUT80), .ZN(n355) );
  OR2_X1 U452 ( .A1(n653), .A2(KEYINPUT2), .ZN(n654) );
  AND2_X1 U453 ( .A1(n528), .A2(n562), .ZN(n346) );
  XOR2_X1 U454 ( .A(KEYINPUT16), .B(G122), .Z(n347) );
  XOR2_X1 U455 ( .A(n583), .B(KEYINPUT47), .Z(n348) );
  AND2_X1 U456 ( .A1(n625), .A2(n561), .ZN(n349) );
  XOR2_X1 U457 ( .A(n711), .B(KEYINPUT82), .Z(n350) );
  XOR2_X1 U458 ( .A(KEYINPUT69), .B(KEYINPUT34), .Z(n351) );
  XNOR2_X1 U459 ( .A(n399), .B(KEYINPUT68), .ZN(n398) );
  XNOR2_X2 U460 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U461 ( .A1(n353), .A2(n352), .ZN(n401) );
  NAND2_X1 U462 ( .A1(n541), .A2(KEYINPUT44), .ZN(n353) );
  NOR2_X1 U463 ( .A1(n354), .A2(n655), .ZN(n656) );
  XNOR2_X1 U464 ( .A(n356), .B(n622), .ZN(G57) );
  NOR2_X2 U465 ( .A1(n621), .A2(n650), .ZN(n356) );
  NAND2_X1 U466 ( .A1(n346), .A2(n349), .ZN(n399) );
  NAND2_X1 U467 ( .A1(n519), .A2(n357), .ZN(n522) );
  XNOR2_X2 U468 ( .A(n515), .B(n514), .ZN(n357) );
  XNOR2_X1 U469 ( .A(n492), .B(n493), .ZN(n359) );
  OR2_X2 U470 ( .A1(n613), .A2(n598), .ZN(n500) );
  INV_X1 U471 ( .A(n674), .ZN(n362) );
  NAND2_X1 U472 ( .A1(n369), .A2(n351), .ZN(n367) );
  INV_X1 U473 ( .A(n544), .ZN(n369) );
  INV_X1 U474 ( .A(n345), .ZN(n375) );
  NAND2_X1 U475 ( .A1(n505), .A2(KEYINPUT19), .ZN(n377) );
  NAND2_X1 U476 ( .A1(n506), .A2(KEYINPUT19), .ZN(n378) );
  XNOR2_X2 U477 ( .A(n379), .B(n512), .ZN(n548) );
  NAND2_X1 U478 ( .A1(n581), .A2(n511), .ZN(n379) );
  NAND2_X1 U479 ( .A1(n585), .A2(n381), .ZN(n380) );
  AND2_X1 U480 ( .A1(n584), .A2(n350), .ZN(n381) );
  XNOR2_X1 U481 ( .A(n401), .B(KEYINPUT87), .ZN(n400) );
  XNOR2_X2 U482 ( .A(n388), .B(G143), .ZN(n490) );
  NOR2_X1 U483 ( .A1(n678), .A2(n504), .ZN(n513) );
  XNOR2_X1 U484 ( .A(n394), .B(n390), .ZN(n641) );
  XNOR2_X1 U485 ( .A(n391), .B(n423), .ZN(n390) );
  INV_X1 U486 ( .A(n441), .ZN(n395) );
  XNOR2_X2 U487 ( .A(n397), .B(n396), .ZN(n652) );
  NAND2_X1 U488 ( .A1(n400), .A2(n398), .ZN(n397) );
  NAND2_X1 U489 ( .A1(n636), .A2(G469), .ZN(n649) );
  NAND2_X1 U490 ( .A1(n636), .A2(G478), .ZN(n643) );
  NAND2_X1 U491 ( .A1(n636), .A2(G217), .ZN(n639) );
  XNOR2_X1 U492 ( .A(n407), .B(n406), .ZN(n585) );
  NAND2_X1 U493 ( .A1(n733), .A2(n734), .ZN(n407) );
  XNOR2_X1 U494 ( .A(n576), .B(n577), .ZN(n734) );
  XNOR2_X1 U495 ( .A(n570), .B(n569), .ZN(n733) );
  NOR2_X2 U496 ( .A1(n616), .A2(n650), .ZN(n617) );
  NOR2_X2 U497 ( .A1(n609), .A2(n650), .ZN(n610) );
  XOR2_X1 U498 ( .A(G131), .B(KEYINPUT4), .Z(n408) );
  XOR2_X1 U499 ( .A(n538), .B(KEYINPUT76), .Z(n409) );
  NOR2_X1 U500 ( .A1(n720), .A2(n348), .ZN(n584) );
  INV_X1 U501 ( .A(KEYINPUT48), .ZN(n592) );
  INV_X1 U502 ( .A(KEYINPUT73), .ZN(n413) );
  INV_X1 U503 ( .A(G134), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n413), .B(G101), .ZN(n414) );
  BUF_X1 U505 ( .A(n674), .Z(n691) );
  INV_X1 U506 ( .A(KEYINPUT71), .ZN(n531) );
  XNOR2_X1 U507 ( .A(n415), .B(n414), .ZN(n417) );
  AND2_X1 U508 ( .A1(n669), .A2(n571), .ZN(n572) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n448) );
  NAND2_X1 U510 ( .A1(G227), .A2(n726), .ZN(n411) );
  XNOR2_X1 U511 ( .A(n344), .B(n412), .ZN(n415) );
  XNOR2_X2 U512 ( .A(n490), .B(n416), .ZN(n423) );
  XNOR2_X1 U513 ( .A(n417), .B(n475), .ZN(n645) );
  NOR2_X1 U514 ( .A1(n645), .A2(G902), .ZN(n418) );
  XNOR2_X1 U515 ( .A(KEYINPUT83), .B(n419), .ZN(n441) );
  XOR2_X1 U516 ( .A(KEYINPUT104), .B(KEYINPUT7), .Z(n421) );
  XNOR2_X1 U517 ( .A(G122), .B(KEYINPUT9), .ZN(n420) );
  XNOR2_X1 U518 ( .A(n421), .B(n420), .ZN(n422) );
  INV_X1 U519 ( .A(G902), .ZN(n481) );
  NAND2_X1 U520 ( .A1(n641), .A2(n481), .ZN(n426) );
  INV_X1 U521 ( .A(G478), .ZN(n425) );
  INV_X1 U522 ( .A(n537), .ZN(n553) );
  XNOR2_X1 U523 ( .A(G113), .B(G122), .ZN(n427) );
  XNOR2_X1 U524 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U525 ( .A(n446), .B(n429), .ZN(n437) );
  XOR2_X1 U526 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n431) );
  NOR2_X1 U527 ( .A1(G953), .A2(G237), .ZN(n470) );
  NAND2_X1 U528 ( .A1(G214), .A2(n470), .ZN(n430) );
  XNOR2_X1 U529 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U530 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n433) );
  XNOR2_X1 U531 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U532 ( .A(n435), .B(n434), .Z(n436) );
  XNOR2_X1 U533 ( .A(n437), .B(n436), .ZN(n606) );
  NOR2_X1 U534 ( .A1(n606), .A2(G902), .ZN(n439) );
  XNOR2_X1 U535 ( .A(KEYINPUT13), .B(G475), .ZN(n438) );
  XNOR2_X1 U536 ( .A(n439), .B(n438), .ZN(n503) );
  XNOR2_X1 U537 ( .A(n503), .B(KEYINPUT103), .ZN(n552) );
  OR2_X1 U538 ( .A1(n553), .A2(n552), .ZN(n715) );
  INV_X1 U539 ( .A(G221), .ZN(n440) );
  NOR2_X1 U540 ( .A1(n441), .A2(n440), .ZN(n445) );
  INV_X1 U541 ( .A(KEYINPUT23), .ZN(n442) );
  XOR2_X1 U542 ( .A(n447), .B(n446), .Z(n723) );
  XNOR2_X1 U543 ( .A(n448), .B(n723), .ZN(n637) );
  NOR2_X1 U544 ( .A1(G902), .A2(n637), .ZN(n455) );
  XNOR2_X1 U545 ( .A(G902), .B(KEYINPUT15), .ZN(n495) );
  NAND2_X1 U546 ( .A1(n495), .A2(G234), .ZN(n450) );
  XNOR2_X1 U547 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n449) );
  XNOR2_X1 U548 ( .A(n450), .B(n449), .ZN(n456) );
  AND2_X1 U549 ( .A1(n456), .A2(G217), .ZN(n451) );
  XNOR2_X1 U550 ( .A(n451), .B(KEYINPUT95), .ZN(n453) );
  XNOR2_X1 U551 ( .A(KEYINPUT25), .B(KEYINPUT72), .ZN(n452) );
  XNOR2_X1 U552 ( .A(n455), .B(n454), .ZN(n529) );
  BUF_X1 U553 ( .A(n529), .Z(n662) );
  AND2_X1 U554 ( .A1(n456), .A2(G221), .ZN(n457) );
  XNOR2_X1 U555 ( .A(KEYINPUT21), .B(n457), .ZN(n661) );
  NAND2_X1 U556 ( .A1(G234), .A2(G237), .ZN(n458) );
  XNOR2_X1 U557 ( .A(n458), .B(KEYINPUT14), .ZN(n461) );
  NAND2_X1 U558 ( .A1(n461), .A2(G952), .ZN(n459) );
  XNOR2_X1 U559 ( .A(n459), .B(KEYINPUT88), .ZN(n688) );
  NOR2_X1 U560 ( .A1(n688), .A2(G953), .ZN(n460) );
  XNOR2_X1 U561 ( .A(n460), .B(KEYINPUT89), .ZN(n509) );
  NAND2_X1 U562 ( .A1(n461), .A2(G902), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n462), .B(KEYINPUT90), .ZN(n507) );
  NOR2_X1 U564 ( .A1(n507), .A2(G900), .ZN(n463) );
  NAND2_X1 U565 ( .A1(G953), .A2(n463), .ZN(n464) );
  NAND2_X1 U566 ( .A1(n509), .A2(n464), .ZN(n586) );
  AND2_X1 U567 ( .A1(n661), .A2(n586), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n465), .B(KEYINPUT67), .ZN(n466) );
  NOR2_X1 U569 ( .A1(n662), .A2(n466), .ZN(n571) );
  XNOR2_X2 U570 ( .A(G101), .B(KEYINPUT3), .ZN(n469) );
  XOR2_X1 U571 ( .A(G137), .B(KEYINPUT5), .Z(n472) );
  NAND2_X1 U572 ( .A1(n470), .A2(G210), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U574 ( .A(n485), .B(n473), .ZN(n474) );
  NAND2_X1 U575 ( .A1(n618), .A2(n481), .ZN(n477) );
  XNOR2_X1 U576 ( .A(G472), .B(KEYINPUT98), .ZN(n476) );
  INV_X1 U577 ( .A(KEYINPUT6), .ZN(n478) );
  XNOR2_X1 U578 ( .A(n669), .B(n478), .ZN(n556) );
  NAND2_X1 U579 ( .A1(n571), .A2(n556), .ZN(n479) );
  NOR2_X1 U580 ( .A1(n715), .A2(n479), .ZN(n482) );
  INV_X1 U581 ( .A(G237), .ZN(n480) );
  NAND2_X1 U582 ( .A1(n481), .A2(n480), .ZN(n496) );
  NAND2_X1 U583 ( .A1(n496), .A2(G214), .ZN(n675) );
  NAND2_X1 U584 ( .A1(n482), .A2(n675), .ZN(n578) );
  INV_X1 U585 ( .A(n578), .ZN(n483) );
  NAND2_X1 U586 ( .A1(n659), .A2(n483), .ZN(n484) );
  XNOR2_X1 U587 ( .A(n484), .B(KEYINPUT43), .ZN(n501) );
  XNOR2_X1 U588 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U589 ( .A(n490), .B(n489), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n726), .A2(G224), .ZN(n491) );
  XNOR2_X1 U591 ( .A(n491), .B(KEYINPUT75), .ZN(n492) );
  INV_X1 U592 ( .A(n495), .ZN(n598) );
  NAND2_X1 U593 ( .A1(n496), .A2(G210), .ZN(n498) );
  INV_X1 U594 ( .A(KEYINPUT79), .ZN(n497) );
  XNOR2_X1 U595 ( .A(n498), .B(n497), .ZN(n499) );
  BUF_X2 U596 ( .A(n345), .Z(n588) );
  AND2_X1 U597 ( .A1(n501), .A2(n588), .ZN(n594) );
  XNOR2_X1 U598 ( .A(G140), .B(KEYINPUT118), .ZN(n502) );
  XOR2_X1 U599 ( .A(n594), .B(n502), .Z(G42) );
  INV_X1 U600 ( .A(n503), .ZN(n536) );
  INV_X1 U601 ( .A(n661), .ZN(n504) );
  INV_X1 U602 ( .A(n675), .ZN(n505) );
  OR2_X1 U603 ( .A1(G898), .A2(n726), .ZN(n631) );
  OR2_X1 U604 ( .A1(n631), .A2(n507), .ZN(n508) );
  AND2_X1 U605 ( .A1(n509), .A2(n508), .ZN(n510) );
  INV_X1 U606 ( .A(KEYINPUT0), .ZN(n512) );
  NAND2_X1 U607 ( .A1(n513), .A2(n548), .ZN(n515) );
  XNOR2_X1 U608 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n514) );
  OR2_X1 U609 ( .A1(n662), .A2(n659), .ZN(n516) );
  OR2_X1 U610 ( .A1(n556), .A2(n516), .ZN(n518) );
  INV_X1 U611 ( .A(KEYINPUT78), .ZN(n517) );
  XNOR2_X1 U612 ( .A(n518), .B(n517), .ZN(n519) );
  INV_X1 U613 ( .A(KEYINPUT77), .ZN(n520) );
  XNOR2_X1 U614 ( .A(n520), .B(KEYINPUT32), .ZN(n521) );
  XNOR2_X1 U615 ( .A(n522), .B(n521), .ZN(n561) );
  XNOR2_X1 U616 ( .A(n561), .B(G119), .ZN(G21) );
  NOR2_X1 U617 ( .A1(n669), .A2(n662), .ZN(n524) );
  INV_X1 U618 ( .A(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U619 ( .A(n528), .B(G110), .ZN(G12) );
  NAND2_X1 U620 ( .A1(n529), .A2(n661), .ZN(n658) );
  NOR2_X1 U621 ( .A1(n530), .A2(n658), .ZN(n532) );
  XNOR2_X1 U622 ( .A(n532), .B(n531), .ZN(n547) );
  NAND2_X1 U623 ( .A1(n547), .A2(n556), .ZN(n535) );
  INV_X1 U624 ( .A(KEYINPUT110), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n533), .B(KEYINPUT33), .ZN(n534) );
  XNOR2_X1 U626 ( .A(n548), .B(KEYINPUT92), .ZN(n544) );
  OR2_X1 U627 ( .A1(n537), .A2(n536), .ZN(n589) );
  XNOR2_X1 U628 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n538) );
  NAND2_X1 U629 ( .A1(n540), .A2(n625), .ZN(n541) );
  XNOR2_X1 U630 ( .A(KEYINPUT97), .B(n543), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n565), .A2(n669), .ZN(n545) );
  NAND2_X1 U632 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U633 ( .A(KEYINPUT99), .B(n546), .Z(n704) );
  AND2_X1 U634 ( .A1(n547), .A2(n669), .ZN(n671) );
  BUF_X1 U635 ( .A(n548), .Z(n549) );
  NAND2_X1 U636 ( .A1(n671), .A2(n549), .ZN(n551) );
  XOR2_X1 U637 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n550) );
  XNOR2_X1 U638 ( .A(n551), .B(n550), .ZN(n718) );
  AND2_X1 U639 ( .A1(n704), .A2(n718), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n553), .A2(n552), .ZN(n717) );
  NAND2_X1 U641 ( .A1(n715), .A2(n717), .ZN(n554) );
  XNOR2_X1 U642 ( .A(KEYINPUT105), .B(n554), .ZN(n680) );
  NOR2_X1 U643 ( .A1(n555), .A2(n680), .ZN(n560) );
  XNOR2_X1 U644 ( .A(n557), .B(KEYINPUT86), .ZN(n558) );
  NAND2_X1 U645 ( .A1(n558), .A2(n662), .ZN(n559) );
  INV_X1 U646 ( .A(KEYINPUT44), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n675), .A2(n669), .ZN(n563) );
  XNOR2_X1 U648 ( .A(KEYINPUT30), .B(n563), .ZN(n564) );
  NOR2_X1 U649 ( .A1(n565), .A2(n564), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n566) );
  XNOR2_X1 U651 ( .A(n588), .B(n566), .ZN(n676) );
  AND2_X1 U652 ( .A1(n676), .A2(n586), .ZN(n567) );
  XNOR2_X1 U653 ( .A(KEYINPUT39), .B(n568), .ZN(n593) );
  NOR2_X1 U654 ( .A1(n593), .A2(n715), .ZN(n570) );
  INV_X1 U655 ( .A(KEYINPUT40), .ZN(n569) );
  XOR2_X1 U656 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n577) );
  XOR2_X1 U657 ( .A(KEYINPUT28), .B(n572), .Z(n574) );
  NAND2_X1 U658 ( .A1(n675), .A2(n676), .ZN(n679) );
  NOR2_X1 U659 ( .A1(n678), .A2(n679), .ZN(n575) );
  XOR2_X1 U660 ( .A(KEYINPUT41), .B(n575), .Z(n657) );
  NAND2_X1 U661 ( .A1(n582), .A2(n657), .ZN(n576) );
  NOR2_X1 U662 ( .A1(n578), .A2(n588), .ZN(n579) );
  XOR2_X1 U663 ( .A(KEYINPUT36), .B(n579), .Z(n580) );
  NOR2_X1 U664 ( .A1(n659), .A2(n580), .ZN(n720) );
  NAND2_X1 U665 ( .A1(n582), .A2(n581), .ZN(n713) );
  AND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n591) );
  NOR2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n711) );
  NOR2_X1 U669 ( .A1(n593), .A2(n717), .ZN(n722) );
  NOR2_X1 U670 ( .A1(n722), .A2(n594), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n602) );
  OR2_X2 U672 ( .A1(n602), .A2(n495), .ZN(n597) );
  AND2_X1 U673 ( .A1(n598), .A2(KEYINPUT2), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT64), .ZN(n605) );
  INV_X1 U676 ( .A(n602), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  NOR2_X1 U678 ( .A1(n604), .A2(n626), .ZN(n655) );
  NOR2_X2 U679 ( .A1(n605), .A2(n655), .ZN(n635) );
  NAND2_X1 U680 ( .A1(n635), .A2(G475), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U683 ( .A1(n635), .A2(G210), .ZN(n615) );
  XNOR2_X1 U684 ( .A(KEYINPUT81), .B(KEYINPUT54), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT55), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U689 ( .A(KEYINPUT63), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n635), .A2(G472), .ZN(n620) );
  XOR2_X1 U691 ( .A(KEYINPUT62), .B(n618), .Z(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(n621) );
  XOR2_X1 U693 ( .A(G101), .B(KEYINPUT112), .Z(n623) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(G3) );
  XNOR2_X1 U695 ( .A(n625), .B(G122), .ZN(G24) );
  NOR2_X1 U696 ( .A1(n626), .A2(G953), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G953), .A2(G224), .ZN(n627) );
  XNOR2_X1 U698 ( .A(KEYINPUT61), .B(n627), .ZN(n628) );
  AND2_X1 U699 ( .A1(n628), .A2(G898), .ZN(n629) );
  NOR2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(G69) );
  BUF_X1 U703 ( .A(n635), .Z(n636) );
  XNOR2_X1 U704 ( .A(n637), .B(KEYINPUT126), .ZN(n638) );
  XNOR2_X1 U705 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U706 ( .A1(n640), .A2(n650), .ZN(G66) );
  XNOR2_X1 U707 ( .A(n641), .B(KEYINPUT125), .ZN(n642) );
  XNOR2_X1 U708 ( .A(n643), .B(n642), .ZN(n644) );
  NOR2_X1 U709 ( .A1(n644), .A2(n650), .ZN(G63) );
  XOR2_X1 U710 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n646) );
  XNOR2_X1 U711 ( .A(n646), .B(KEYINPUT58), .ZN(n647) );
  XNOR2_X1 U712 ( .A(n645), .B(n647), .ZN(n648) );
  XNOR2_X1 U713 ( .A(n649), .B(n648), .ZN(n651) );
  NOR2_X1 U714 ( .A1(n651), .A2(n650), .ZN(G54) );
  NOR2_X1 U715 ( .A1(n652), .A2(n602), .ZN(n653) );
  XNOR2_X1 U716 ( .A(n656), .B(KEYINPUT84), .ZN(n698) );
  INV_X1 U717 ( .A(n657), .ZN(n692) );
  NAND2_X1 U718 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U719 ( .A(KEYINPUT50), .B(n660), .ZN(n667) );
  NOR2_X1 U720 ( .A1(n662), .A2(n661), .ZN(n664) );
  XNOR2_X1 U721 ( .A(KEYINPUT120), .B(KEYINPUT49), .ZN(n663) );
  XNOR2_X1 U722 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U723 ( .A(KEYINPUT119), .B(n665), .Z(n666) );
  NAND2_X1 U724 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U725 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U726 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U727 ( .A(KEYINPUT51), .B(n672), .Z(n673) );
  NOR2_X1 U728 ( .A1(n692), .A2(n673), .ZN(n686) );
  NOR2_X1 U729 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U730 ( .A1(n678), .A2(n677), .ZN(n683) );
  NOR2_X1 U731 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U732 ( .A(KEYINPUT121), .B(n681), .Z(n682) );
  NOR2_X1 U733 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U734 ( .A1(n691), .A2(n684), .ZN(n685) );
  NOR2_X1 U735 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U736 ( .A(n687), .B(KEYINPUT52), .ZN(n689) );
  NOR2_X1 U737 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U738 ( .A(KEYINPUT122), .B(n690), .Z(n696) );
  NOR2_X1 U739 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U740 ( .A(KEYINPUT123), .B(n693), .Z(n694) );
  NOR2_X1 U741 ( .A1(n694), .A2(G953), .ZN(n695) );
  NAND2_X1 U742 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U743 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U744 ( .A(n699), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U745 ( .A1(n715), .A2(n704), .ZN(n701) );
  XNOR2_X1 U746 ( .A(G104), .B(KEYINPUT113), .ZN(n700) );
  XNOR2_X1 U747 ( .A(n701), .B(n700), .ZN(G6) );
  XOR2_X1 U748 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n703) );
  XNOR2_X1 U749 ( .A(n341), .B(KEYINPUT26), .ZN(n702) );
  XNOR2_X1 U750 ( .A(n703), .B(n702), .ZN(n706) );
  NOR2_X1 U751 ( .A1(n717), .A2(n704), .ZN(n705) );
  XOR2_X1 U752 ( .A(n706), .B(n705), .Z(G9) );
  NOR2_X1 U753 ( .A1(n713), .A2(n717), .ZN(n710) );
  XOR2_X1 U754 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n708) );
  XNOR2_X1 U755 ( .A(G128), .B(KEYINPUT116), .ZN(n707) );
  XNOR2_X1 U756 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U757 ( .A(n710), .B(n709), .ZN(G30) );
  XNOR2_X1 U758 ( .A(G143), .B(n711), .ZN(n712) );
  XNOR2_X1 U759 ( .A(n712), .B(KEYINPUT117), .ZN(G45) );
  NOR2_X1 U760 ( .A1(n713), .A2(n715), .ZN(n714) );
  XOR2_X1 U761 ( .A(G146), .B(n714), .Z(G48) );
  NOR2_X1 U762 ( .A1(n718), .A2(n715), .ZN(n716) );
  XOR2_X1 U763 ( .A(G113), .B(n716), .Z(G15) );
  NOR2_X1 U764 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U765 ( .A(G116), .B(n719), .Z(G18) );
  XNOR2_X1 U766 ( .A(G125), .B(n720), .ZN(n721) );
  XNOR2_X1 U767 ( .A(n721), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U768 ( .A(G134), .B(n722), .Z(G36) );
  XOR2_X1 U769 ( .A(n723), .B(KEYINPUT127), .Z(n724) );
  XNOR2_X1 U770 ( .A(n725), .B(n724), .ZN(n728) );
  XNOR2_X1 U771 ( .A(n343), .B(n728), .ZN(n727) );
  NAND2_X1 U772 ( .A1(n727), .A2(n726), .ZN(n732) );
  XNOR2_X1 U773 ( .A(G227), .B(n728), .ZN(n729) );
  NAND2_X1 U774 ( .A1(n729), .A2(G900), .ZN(n730) );
  NAND2_X1 U775 ( .A1(n730), .A2(G953), .ZN(n731) );
  NAND2_X1 U776 ( .A1(n732), .A2(n731), .ZN(G72) );
  XNOR2_X1 U777 ( .A(G131), .B(n733), .ZN(G33) );
  XNOR2_X1 U778 ( .A(G137), .B(n734), .ZN(G39) );
endmodule

