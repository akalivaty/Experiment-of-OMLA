//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1221,
    new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n459), .B1(new_n449), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  NOR3_X1   g047(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n467), .B2(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT69), .A4(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n468), .A3(new_n466), .ZN(new_n478));
  OR2_X1    g053(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(G137), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n477), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n464), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(G113), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n468), .ZN(new_n486));
  INV_X1    g061(.A(G125), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n470), .A2(new_n471), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G160));
  NOR2_X1   g068(.A1(new_n478), .A2(new_n489), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  OAI221_X1 g070(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n489), .C2(G112), .ZN(new_n496));
  INV_X1    g071(.A(G136), .ZN(new_n497));
  INV_X1    g072(.A(new_n478), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(new_n462), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT71), .ZN(G162));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(G126), .A2(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n475), .A2(new_n466), .A3(new_n468), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n507), .A2(new_n508), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n479), .A2(G138), .A3(new_n480), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n512), .B(KEYINPUT4), .C1(new_n478), .C2(new_n513), .ZN(new_n514));
  NOR3_X1   g089(.A1(new_n513), .A2(new_n486), .A3(KEYINPUT4), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT4), .B1(new_n478), .B2(new_n513), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT73), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n511), .B1(new_n514), .B2(new_n517), .ZN(G164));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT5), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G62), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n521), .B2(new_n523), .ZN(new_n532));
  NAND2_X1  g107(.A1(G75), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(G651), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g113(.A(KEYINPUT76), .B(G651), .C1(new_n532), .C2(new_n535), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n530), .B1(new_n538), .B2(new_n539), .ZN(G166));
  INV_X1    g115(.A(new_n526), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n541), .A2(G89), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  INV_X1    g120(.A(G51), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n543), .B(new_n545), .C1(new_n546), .C2(new_n528), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n542), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  INV_X1    g127(.A(G52), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n526), .A2(new_n552), .B1(new_n528), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  AOI22_X1  g130(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n550), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT77), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n525), .A2(G543), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n541), .A2(G81), .B1(new_n559), .B2(G43), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT78), .ZN(G188));
  XOR2_X1   g144(.A(KEYINPUT79), .B(KEYINPUT9), .Z(new_n570));
  NAND3_X1  g145(.A1(new_n559), .A2(G53), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n528), .A2(new_n572), .B1(new_n573), .B2(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n524), .A2(KEYINPUT81), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n521), .B2(new_n523), .ZN(new_n580));
  OAI21_X1  g155(.A(G65), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G78), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n519), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n550), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n541), .A2(G91), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n577), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  INV_X1    g165(.A(G168), .ZN(G286));
  INV_X1    g166(.A(G166), .ZN(G303));
  OAI21_X1  g167(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n593));
  INV_X1    g168(.A(G49), .ZN(new_n594));
  INV_X1    g169(.A(G87), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n594), .B2(new_n528), .C1(new_n595), .C2(new_n526), .ZN(G288));
  AOI22_X1  g171(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n550), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  INV_X1    g174(.A(G48), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n526), .A2(new_n599), .B1(new_n528), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(new_n559), .A2(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OAI221_X1 g181(.A(new_n604), .B1(new_n605), .B2(new_n526), .C1(new_n550), .C2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT82), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n524), .B(KEYINPUT81), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n610), .A2(G66), .ZN(new_n611));
  AND2_X1   g186(.A1(G79), .A2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n541), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n526), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n614), .A2(new_n617), .B1(G54), .B2(new_n559), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n609), .B1(G868), .B2(new_n620), .ZN(G284));
  OAI21_X1  g196(.A(new_n609), .B1(G868), .B2(new_n620), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n577), .A2(new_n588), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(G148));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n561), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n619), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g208(.A(new_n486), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n465), .A2(G2105), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT13), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n637), .A2(new_n638), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n498), .A2(G135), .A3(new_n462), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT84), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n494), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n489), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(G2096), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n642), .A2(new_n649), .A3(new_n650), .ZN(G156));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n655), .B(new_n661), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n663), .ZN(G401));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT17), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(new_n670), .B2(new_n668), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT85), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(new_n670), .A3(new_n668), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n670), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n669), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  AOI211_X1 g268(.A(new_n691), .B(new_n693), .C1(new_n686), .C2(new_n690), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT86), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n695), .B(new_n700), .ZN(G229));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT26), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n704), .A2(new_n705), .B1(G105), .B2(new_n635), .ZN(new_n706));
  INV_X1    g281(.A(G141), .ZN(new_n707));
  INV_X1    g282(.A(G129), .ZN(new_n708));
  INV_X1    g283(.A(new_n494), .ZN(new_n709));
  OAI221_X1 g284(.A(new_n706), .B1(new_n499), .B2(new_n707), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(KEYINPUT97), .C1(G29), .C2(G32), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(KEYINPUT97), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G2084), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(KEYINPUT24), .B2(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(KEYINPUT24), .B2(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n492), .B2(G29), .ZN(new_n721));
  OAI22_X1  g296(.A1(new_n714), .A2(new_n716), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT96), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n489), .A2(G103), .A3(G2104), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT94), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT25), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(KEYINPUT25), .ZN(new_n727));
  INV_X1    g302(.A(G139), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n726), .A2(new_n727), .B1(new_n728), .B2(new_n499), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI221_X1 g306(.A(KEYINPUT95), .B1(new_n728), .B2(new_n499), .C1(new_n726), .C2(new_n727), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n634), .A2(G127), .ZN(new_n734));
  NAND2_X1  g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n489), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n723), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(KEYINPUT96), .B(new_n736), .C1(new_n731), .C2(new_n732), .ZN(new_n739));
  OAI21_X1  g314(.A(G29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G33), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(G29), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2072), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n722), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT98), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n718), .A2(G25), .ZN(new_n749));
  OAI221_X1 g324(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n489), .C2(G107), .ZN(new_n750));
  INV_X1    g325(.A(G119), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n709), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n499), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(G131), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(new_n718), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT35), .B(G1991), .Z(new_n756));
  XOR2_X1   g331(.A(new_n755), .B(new_n756), .Z(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G24), .ZN(new_n758));
  XNOR2_X1  g333(.A(G290), .B(KEYINPUT87), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT88), .B(G1986), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n757), .B(new_n762), .C1(KEYINPUT90), .C2(KEYINPUT36), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G23), .ZN(new_n765));
  INV_X1    g340(.A(G288), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(new_n764), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT33), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1976), .ZN(new_n769));
  NOR2_X1   g344(.A1(G6), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n602), .B2(G16), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT32), .B(G1981), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n764), .A2(G22), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT89), .Z(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G166), .B2(new_n764), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G1971), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(G1971), .ZN(new_n778));
  AND3_X1   g353(.A1(new_n773), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n769), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT34), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT34), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n763), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n746), .B2(new_n747), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n561), .A2(G16), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n764), .A2(G19), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G1341), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT91), .B(G1348), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n620), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n791), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n764), .A2(G20), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT23), .Z(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G299), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1956), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n718), .A2(G27), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G164), .B2(new_n718), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2078), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n721), .A2(new_n717), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n789), .B2(new_n790), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n796), .A2(new_n801), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n795), .A2(new_n792), .B1(new_n714), .B2(new_n716), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n648), .A2(new_n718), .ZN(new_n809));
  NOR2_X1   g384(.A1(G171), .A2(new_n764), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G5), .B2(new_n764), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n764), .A2(G21), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G168), .B2(new_n764), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT99), .B(G1966), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n811), .A2(new_n812), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n809), .B(new_n817), .C1(new_n814), .C2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n718), .A2(G26), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT28), .ZN(new_n820));
  INV_X1    g395(.A(G140), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n489), .A2(G116), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n499), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(G128), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n709), .A2(KEYINPUT92), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT92), .B1(new_n709), .B2(new_n825), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n820), .B1(new_n828), .B2(new_n718), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT93), .B(G2067), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT31), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(G11), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(G11), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT30), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(G28), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n718), .B1(new_n835), .B2(G28), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n833), .B(new_n834), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n811), .B2(new_n812), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n808), .A2(new_n818), .A3(new_n831), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n718), .A2(G35), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G162), .B2(new_n718), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(G2090), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(G2090), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n840), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n807), .B(new_n847), .C1(new_n783), .C2(new_n784), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n748), .A2(new_n786), .A3(new_n848), .ZN(G311));
  INV_X1    g424(.A(G311), .ZN(G150));
  AOI22_X1  g425(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n550), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n526), .A2(new_n853), .B1(new_n528), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n620), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n561), .A2(new_n857), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n558), .A2(new_n560), .A3(new_n856), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n861), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT101), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n869));
  INV_X1    g444(.A(new_n865), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n870), .B2(KEYINPUT39), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n868), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n859), .B1(new_n872), .B2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n648), .B(G160), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  INV_X1    g452(.A(new_n738), .ZN(new_n878));
  INV_X1    g453(.A(new_n739), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n881));
  INV_X1    g456(.A(new_n515), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n514), .A3(new_n882), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n507), .A2(new_n508), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n507), .A2(new_n508), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n504), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT103), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n888), .A2(new_n828), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n828), .ZN(new_n890));
  OR3_X1    g465(.A1(new_n889), .A2(new_n890), .A3(new_n711), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n711), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n880), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n878), .A2(new_n879), .A3(new_n877), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT104), .B1(new_n738), .B2(new_n739), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n494), .A2(G130), .ZN(new_n898));
  OAI221_X1 g473(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n489), .C2(G118), .ZN(new_n899));
  INV_X1    g474(.A(G142), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n499), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(new_n637), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n754), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT105), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n893), .A2(new_n897), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n893), .B2(new_n897), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n876), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n893), .A2(new_n897), .A3(new_n903), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n876), .B(KEYINPUT106), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n893), .A2(new_n897), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n908), .B(new_n909), .C1(new_n910), .C2(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n907), .A2(new_n911), .A3(new_n912), .A4(new_n914), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(G395));
  NAND2_X1  g493(.A1(new_n624), .A2(new_n620), .ZN(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(new_n619), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n864), .B(new_n631), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n921), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n926), .ZN(new_n929));
  XNOR2_X1  g504(.A(G166), .B(G290), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n602), .B(G288), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n931), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n930), .B(new_n931), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT108), .B1(new_n932), .B2(new_n934), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n935), .B1(new_n940), .B2(new_n933), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n929), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n929), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(G868), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n857), .A2(new_n629), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(G295));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n947));
  XNOR2_X1  g522(.A(G295), .B(new_n947), .ZN(G331));
  INV_X1    g523(.A(new_n863), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n856), .B1(new_n558), .B2(new_n560), .ZN(new_n950));
  OAI21_X1  g525(.A(G171), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n862), .A2(G301), .A3(new_n863), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(G168), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G168), .B1(new_n951), .B2(new_n952), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n928), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n949), .A2(G171), .A3(new_n950), .ZN(new_n957));
  AOI21_X1  g532(.A(G301), .B1(new_n862), .B2(new_n863), .ZN(new_n958));
  OAI21_X1  g533(.A(G286), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(new_n923), .A3(new_n953), .A4(new_n924), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(KEYINPUT110), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n912), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n956), .A2(new_n940), .A3(new_n960), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n940), .B1(new_n956), .B2(new_n960), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(KEYINPUT110), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT112), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n956), .A2(new_n960), .ZN(new_n970));
  INV_X1    g545(.A(new_n940), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n956), .A2(new_n940), .A3(new_n960), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n966), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n962), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT43), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n972), .B2(new_n973), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n980), .B2(new_n968), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n969), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n974), .A2(new_n975), .A3(new_n983), .A4(new_n968), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n974), .A2(new_n968), .A3(new_n975), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT111), .B1(new_n980), .B2(new_n968), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n979), .B(new_n984), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n982), .A2(new_n987), .ZN(G397));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(G164), .B2(G1384), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n483), .A2(G40), .A3(new_n491), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n989), .B1(new_n994), .B2(G1996), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(KEYINPUT46), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G2067), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n828), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n993), .B1(new_n999), .B2(new_n710), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT127), .Z(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT47), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n710), .B(G1996), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n999), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n754), .B(new_n756), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n993), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G290), .A2(G1986), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n993), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT48), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(KEYINPUT48), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n828), .A2(new_n998), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n754), .A2(new_n756), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n993), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1003), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  NOR3_X1   g595(.A1(G166), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1971), .ZN(new_n1024));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n887), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(new_n990), .ZN(new_n1027));
  INV_X1    g602(.A(new_n992), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n883), .B2(new_n886), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(KEYINPUT45), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1024), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1032));
  INV_X1    g607(.A(G2090), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .A4(new_n1028), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1023), .B1(new_n1037), .B2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n602), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G1981), .B1(new_n598), .B2(new_n601), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT114), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G305), .A2(new_n1043), .A3(G1981), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT115), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1020), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1042), .A2(new_n1044), .A3(KEYINPUT115), .A4(new_n1046), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n766), .A2(G1976), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT52), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1038), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G168), .A2(G8), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n992), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n717), .A4(new_n1035), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n815), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1032), .A2(new_n717), .A3(new_n1035), .A4(new_n1028), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT116), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1061), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1037), .A2(G8), .A3(new_n1023), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1059), .A2(new_n1060), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1051), .A2(new_n1053), .A3(new_n766), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1040), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1051), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1020), .B(new_n1022), .C1(new_n1031), .C2(new_n1036), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1073), .A2(new_n1049), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1038), .A2(new_n1075), .A3(new_n1058), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1060), .B1(new_n1078), .B2(new_n1069), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1037), .A2(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1022), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1083));
  INV_X1    g658(.A(G2078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n991), .A2(new_n1084), .A3(new_n1085), .A4(new_n1028), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n992), .B1(new_n1026), .B2(new_n990), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT53), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1032), .A2(new_n1035), .A3(new_n1028), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n812), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1068), .A2(G168), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1096), .A2(new_n1097), .A3(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1028), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1100));
  AOI211_X1 g675(.A(KEYINPUT50), .B(G1384), .C1(new_n883), .C2(new_n886), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1100), .A2(new_n1101), .A3(G2084), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n1063), .ZN(new_n1103));
  OAI21_X1  g678(.A(G286), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(G8), .A3(new_n1096), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1105), .B2(KEYINPUT51), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1095), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G168), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1096), .A2(G8), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT51), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1098), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(KEYINPUT62), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1080), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT45), .B1(new_n887), .B2(new_n1025), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n476), .A2(new_n482), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT123), .B1(new_n1119), .B2(new_n464), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n483), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G40), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n488), .B2(new_n490), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1117), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1124), .B1(new_n483), .B2(new_n1121), .ZN(new_n1127));
  AOI211_X1 g702(.A(KEYINPUT123), .B(new_n464), .C1(new_n476), .C2(new_n482), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(KEYINPUT124), .C1(KEYINPUT45), .C2(new_n1029), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1084), .A2(KEYINPUT53), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n1029), .B2(KEYINPUT45), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1126), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1088), .A2(new_n1133), .A3(new_n1092), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1116), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1087), .A2(new_n1086), .B1(new_n1091), .B2(new_n812), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(G301), .A4(new_n1090), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1088), .A2(new_n1092), .A3(new_n1090), .A4(G301), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT125), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1136), .B2(new_n1090), .ZN(new_n1142));
  AND4_X1   g717(.A1(G301), .A2(new_n1088), .A3(new_n1133), .A4(new_n1092), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1116), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1144), .A3(new_n1078), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT126), .B1(new_n1145), .B2(new_n1106), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1136), .A2(G301), .A3(new_n1133), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT54), .B1(new_n1094), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(new_n1083), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1113), .A2(new_n1149), .A3(new_n1150), .A4(new_n1141), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n991), .A2(new_n1028), .A3(new_n1085), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(G1996), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(new_n790), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n562), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n562), .B(new_n1160), .C1(new_n1154), .C2(new_n1157), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1153), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT56), .B(G2072), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1166), .A2(new_n1167), .B1(new_n1091), .B2(new_n800), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n583), .B1(new_n610), .B2(G65), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1169), .B(new_n586), .C1(new_n1170), .C2(new_n550), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT117), .B1(new_n585), .B2(new_n587), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(new_n575), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT57), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n1175), .A2(KEYINPUT118), .B1(new_n1174), .B2(G299), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(KEYINPUT118), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1168), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(G299), .A2(new_n1174), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT118), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1167), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1184), .A2(G1956), .B1(new_n1153), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1183), .A2(new_n1186), .A3(new_n1177), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1179), .A2(new_n1187), .A3(KEYINPUT61), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT60), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1091), .A2(new_n792), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1029), .A2(new_n1028), .A3(new_n998), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1189), .B1(new_n1192), .B2(new_n619), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1193), .B1(new_n619), .B2(new_n1192), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1192), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1195), .A2(new_n1189), .A3(new_n620), .ZN(new_n1196));
  AND4_X1   g771(.A1(new_n1165), .A2(new_n1188), .A3(new_n1194), .A4(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1183), .A2(new_n1186), .A3(KEYINPUT121), .A4(new_n1177), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1179), .A2(new_n1187), .A3(new_n1201), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1200), .A2(KEYINPUT122), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(KEYINPUT122), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1197), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1187), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1195), .A2(new_n619), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1206), .B1(new_n1179), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1115), .B1(new_n1152), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1008), .A2(KEYINPUT113), .ZN(new_n1211));
  NAND2_X1  g786(.A1(G290), .A2(G1986), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1007), .B1(new_n994), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1017), .B1(new_n1210), .B2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g790(.A1(G229), .A2(G227), .A3(G401), .A4(new_n460), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n913), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g792(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n1219));
  NOR2_X1   g793(.A1(new_n1218), .A2(new_n1219), .ZN(G308));
  OAI21_X1  g794(.A(KEYINPUT43), .B1(new_n965), .B2(G37), .ZN(new_n1221));
  OAI211_X1 g795(.A(new_n1221), .B(KEYINPUT111), .C1(new_n976), .C2(KEYINPUT43), .ZN(new_n1222));
  NAND4_X1  g796(.A1(new_n1222), .A2(new_n913), .A3(new_n984), .A4(new_n1217), .ZN(G225));
endmodule


