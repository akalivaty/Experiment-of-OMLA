//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116, new_n1117;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(KEYINPUT68), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT67), .B(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(new_n461), .A3(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(G137), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n465), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(G160));
  AOI21_X1  g054(.A(KEYINPUT68), .B1(new_n473), .B2(KEYINPUT3), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n467), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n465), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  NOR3_X1   g061(.A1(new_n473), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n474), .A2(new_n466), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n469), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(new_n469), .B2(G114), .ZN(new_n493));
  NOR2_X1   g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT3), .B(G2104), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n465), .A3(G138), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(KEYINPUT4), .B(G138), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n489), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT69), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(G88), .B1(G50), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND2_X1  g102(.A1(new_n523), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n521), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n522), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n516), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(G651), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT71), .B(G81), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n523), .A2(new_n549), .B1(new_n524), .B2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n524), .A2(KEYINPUT72), .A3(G53), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n516), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n523), .A2(G91), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n559), .A2(new_n560), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  OAI21_X1  g143(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(KEYINPUT73), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n569), .A2(KEYINPUT73), .B1(new_n524), .B2(G49), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n523), .A2(G87), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n524), .A2(G48), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  OAI221_X1 g151(.A(new_n574), .B1(new_n575), .B2(new_n522), .C1(new_n576), .C2(new_n536), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT74), .ZN(G305));
  NAND2_X1  g153(.A1(new_n524), .A2(G47), .ZN(new_n579));
  XOR2_X1   g154(.A(KEYINPUT75), .B(G85), .Z(new_n580));
  AOI22_X1  g155(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n522), .B2(new_n580), .C1(new_n581), .C2(new_n536), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n522), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n516), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n584), .A2(new_n587), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n524), .A2(G54), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n583), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n583), .B1(new_n594), .B2(G868), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G299), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  XNOR2_X1  g174(.A(G297), .B(KEYINPUT76), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NOR2_X1   g177(.A1(new_n593), .A2(G559), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n483), .A2(G123), .ZN(new_n608));
  OAI221_X1 g183(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n465), .C2(G111), .ZN(new_n609));
  INV_X1    g184(.A(G135), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n490), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(KEYINPUT78), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2096), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  NAND2_X1  g191(.A1(KEYINPUT77), .A2(G2100), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n616), .B(new_n617), .Z(new_n618));
  OAI211_X1 g193(.A(new_n613), .B(new_n618), .C1(KEYINPUT77), .C2(G2100), .ZN(G156));
  XNOR2_X1  g194(.A(G2451), .B(G2454), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G1341), .B(G1348), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2435), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2438), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n625), .B(new_n630), .Z(new_n631));
  AND2_X1   g206(.A1(new_n631), .A2(G14), .ZN(G401));
  XNOR2_X1  g207(.A(G2067), .B(G2678), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n638), .B1(KEYINPUT17), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(new_n637), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n641), .B(new_n642), .C1(KEYINPUT17), .C2(new_n640), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n639), .B(KEYINPUT82), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n640), .A3(new_n633), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n643), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2100), .Z(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(KEYINPUT84), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G229));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n594), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G4), .B2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(G1348), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G35), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G162), .B2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT98), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G2090), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n552), .A2(new_n674), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n674), .B2(G19), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(G1341), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n676), .A2(new_n677), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n684), .B(new_n690), .C1(G1341), .C2(new_n687), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n683), .A2(G2090), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n679), .A2(G26), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G128), .ZN(new_n696));
  OAI221_X1 g271(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n465), .C2(G116), .ZN(new_n697));
  INV_X1    g272(.A(G140), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n490), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n695), .B1(new_n699), .B2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G2067), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n674), .A2(G20), .ZN(new_n703));
  OAI211_X1 g278(.A(KEYINPUT23), .B(new_n703), .C1(new_n598), .C2(new_n674), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(KEYINPUT23), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G1956), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR4_X1   g282(.A1(new_n691), .A2(new_n692), .A3(new_n702), .A4(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n490), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G139), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n496), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(new_n465), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT25), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT93), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G33), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(G29), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2072), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(KEYINPUT94), .A3(G2072), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n709), .A2(G141), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n483), .A2(G129), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n469), .A2(G105), .A3(G2104), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n727), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  MUX2_X1   g308(.A(G32), .B(new_n733), .S(G29), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n721), .A2(G2072), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n679), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n679), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2078), .ZN(new_n740));
  NAND2_X1  g315(.A1(G171), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G5), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT96), .B(KEYINPUT30), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G28), .Z(new_n745));
  AOI22_X1  g320(.A1(new_n742), .A2(new_n743), .B1(new_n679), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n743), .B2(new_n742), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n740), .B(new_n747), .C1(G29), .C2(new_n612), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G11), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n674), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n674), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1966), .ZN(new_n752));
  OR2_X1    g327(.A1(KEYINPUT24), .A2(G34), .ZN(new_n753));
  NAND2_X1  g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n753), .A2(new_n679), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G160), .B2(new_n679), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2084), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n748), .A2(new_n749), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n737), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n726), .A2(new_n736), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n708), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n679), .A2(G25), .ZN(new_n766));
  OAI221_X1 g341(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n465), .C2(G107), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT87), .Z(new_n768));
  AOI22_X1  g343(.A1(new_n709), .A2(G131), .B1(G119), .B2(new_n483), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(new_n679), .ZN(new_n772));
  MUX2_X1   g347(.A(new_n766), .B(new_n772), .S(KEYINPUT86), .Z(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT35), .B(G1991), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n773), .B(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G24), .B(G290), .S(G16), .Z(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1986), .Z(new_n778));
  MUX2_X1   g353(.A(G6), .B(G305), .S(G16), .Z(new_n779));
  XOR2_X1   g354(.A(KEYINPUT32), .B(G1981), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n674), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n674), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT33), .ZN(new_n785));
  INV_X1    g360(.A(G1976), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  INV_X1    g363(.A(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(KEYINPUT88), .B1(new_n789), .B2(G16), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n789), .A2(KEYINPUT88), .A3(G16), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n790), .B(new_n791), .C1(G166), .C2(new_n674), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1971), .Z(new_n793));
  NAND4_X1  g368(.A1(new_n781), .A2(new_n787), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n776), .B(new_n778), .C1(new_n794), .C2(KEYINPUT34), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT89), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(KEYINPUT90), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n795), .A2(new_n796), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n797), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n800), .A3(new_n801), .ZN(new_n803));
  INV_X1    g378(.A(new_n799), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n798), .A2(KEYINPUT90), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AND4_X1   g381(.A1(new_n678), .A2(new_n765), .A3(new_n802), .A4(new_n806), .ZN(G311));
  NAND4_X1  g382(.A1(new_n765), .A2(new_n802), .A3(new_n806), .A4(new_n678), .ZN(G150));
  NAND2_X1  g383(.A1(G80), .A2(G543), .ZN(new_n809));
  INV_X1    g384(.A(G67), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n516), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G651), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n524), .A2(G55), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n522), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(G860), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  AOI21_X1  g394(.A(new_n552), .B1(new_n817), .B2(new_n816), .ZN(new_n820));
  INV_X1    g395(.A(new_n815), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n551), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(KEYINPUT101), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n816), .A2(new_n817), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n551), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n826));
  INV_X1    g401(.A(new_n822), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n594), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT102), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n819), .B1(new_n835), .B2(G860), .ZN(G145));
  AOI22_X1  g411(.A1(new_n709), .A2(G142), .B1(G130), .B2(new_n483), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(KEYINPUT104), .ZN(new_n839));
  OR3_X1    g414(.A1(new_n465), .A2(KEYINPUT103), .A3(G118), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT103), .B1(new_n465), .B2(G118), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(KEYINPUT104), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n837), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n615), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n699), .B(new_n506), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n732), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n717), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n733), .B(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n718), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n771), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n851), .A2(new_n771), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n845), .A3(new_n852), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n612), .B(G160), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n491), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n860), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT40), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n861), .A2(new_n866), .A3(new_n862), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(G395));
  NAND2_X1  g443(.A1(new_n829), .A2(new_n603), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n823), .A2(new_n604), .A3(new_n828), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n594), .A2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n598), .A2(new_n593), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(KEYINPUT41), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n869), .A2(new_n874), .A3(new_n870), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(KEYINPUT42), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(G303), .B(G290), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G305), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G288), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n882), .A2(new_n883), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(G868), .B2(new_n824), .ZN(G295));
  OAI21_X1  g467(.A(new_n891), .B1(G868), .B2(new_n824), .ZN(G331));
  XOR2_X1   g468(.A(G286), .B(G171), .Z(new_n894));
  NAND3_X1  g469(.A1(new_n823), .A2(new_n828), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n823), .B2(new_n828), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n878), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n895), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n874), .B1(new_n899), .B2(new_n896), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n887), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n862), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n874), .A2(new_n876), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n897), .A2(new_n895), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n900), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT106), .B1(new_n908), .B2(new_n889), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  AOI211_X1 g485(.A(new_n910), .B(new_n887), .C1(new_n907), .C2(new_n900), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n903), .B(new_n904), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT107), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n887), .B1(new_n907), .B2(new_n900), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT106), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n904), .A4(new_n903), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n887), .B1(new_n898), .B2(new_n900), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n902), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(KEYINPUT43), .A3(new_n903), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n904), .B1(new_n902), .B2(new_n918), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(G397));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  OAI21_X1  g503(.A(G138), .B1(new_n500), .B2(new_n501), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n498), .B1(new_n929), .B2(new_n475), .ZN(new_n930));
  INV_X1    g505(.A(new_n495), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n482), .B1(new_n503), .B2(new_n502), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n477), .A2(new_n478), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT108), .B(G40), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n937), .A2(new_n470), .A3(new_n468), .A4(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n941), .A2(G1996), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(new_n733), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT109), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n699), .B(new_n701), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n732), .A2(G1996), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n770), .A2(new_n774), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n699), .A2(G2067), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n941), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n771), .A2(new_n775), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n940), .B1(new_n953), .B2(new_n949), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n941), .A2(G1986), .A3(G290), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT48), .Z(new_n956));
  AND3_X1   g531(.A1(new_n948), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n942), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(KEYINPUT46), .ZN(new_n959));
  INV_X1    g534(.A(new_n945), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n940), .B1(new_n960), .B2(new_n732), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(KEYINPUT46), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(KEYINPUT47), .Z(new_n964));
  NOR3_X1   g539(.A1(new_n952), .A2(new_n957), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n783), .A2(G1976), .ZN(new_n966));
  INV_X1    g541(.A(G8), .ZN(new_n967));
  INV_X1    g542(.A(new_n939), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n499), .B2(new_n505), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n783), .A2(G1976), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n971), .A2(KEYINPUT52), .A3(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT112), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(KEYINPUT52), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT111), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n577), .B(G1981), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n970), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n978), .B2(new_n977), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT113), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n939), .B1(new_n934), .B2(KEYINPUT50), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n969), .A2(KEYINPUT110), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT110), .B1(new_n969), .B2(new_n985), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n988), .A2(G2090), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n939), .B1(new_n934), .B2(new_n935), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT45), .B(new_n928), .C1(new_n932), .C2(new_n933), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(G1971), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n967), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G303), .A2(G8), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT55), .Z(new_n996));
  AND2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT63), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n974), .A2(new_n981), .A3(new_n1000), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n994), .A2(new_n996), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n983), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n969), .A2(KEYINPUT115), .A3(KEYINPUT45), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n991), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n990), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1966), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(G2084), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n984), .B(new_n1010), .C1(new_n986), .C2(new_n987), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n967), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G168), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT63), .B1(new_n1003), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n983), .A2(new_n997), .A3(new_n1001), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n980), .A2(G1976), .A3(G288), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n577), .A2(G1981), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n970), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G2078), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT53), .B1(new_n992), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT123), .B(G1961), .Z(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n988), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1007), .A2(new_n1024), .A3(G2078), .ZN(new_n1025));
  AOI21_X1  g600(.A(G301), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT126), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1009), .A2(G168), .A3(new_n1011), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT121), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1030), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1030), .A2(KEYINPUT121), .A3(G8), .A4(new_n1031), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1012), .A2(G286), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(KEYINPUT122), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT122), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1027), .A2(KEYINPUT126), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1049), .B2(new_n1041), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1029), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1003), .A2(G168), .A3(new_n1012), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n477), .B(KEYINPUT124), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n478), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n936), .A2(new_n1055), .A3(G40), .A4(new_n991), .ZN(new_n1056));
  OR4_X1    g631(.A1(new_n1024), .A2(new_n1056), .A3(G2078), .A4(new_n471), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1023), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1053), .B1(new_n1058), .B2(G171), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT125), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1023), .A2(G301), .A3(new_n1025), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1049), .A2(new_n1041), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1058), .A2(G171), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1053), .B1(new_n1066), .B2(new_n1026), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n988), .A2(new_n677), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n968), .A2(new_n969), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n1069), .B2(G2067), .ZN(new_n1070));
  OR3_X1    g645(.A1(new_n1069), .A2(KEYINPUT118), .A3(G2067), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n992), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n565), .B2(KEYINPUT117), .ZN(new_n1075));
  XNOR2_X1  g650(.A(G299), .B(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n984), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n706), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1072), .A2(new_n1080), .A3(new_n594), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1076), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1080), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT61), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1080), .A3(KEYINPUT61), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1072), .A2(KEYINPUT60), .A3(new_n594), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n593), .B(KEYINPUT60), .Z(new_n1090));
  OR2_X1    g665(.A1(new_n1072), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(G1996), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n992), .A2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1069), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n551), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT59), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1081), .B(new_n1084), .C1(new_n1092), .C2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .A4(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1051), .A2(new_n1052), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n993), .B1(G2090), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(new_n967), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n996), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1108), .A2(new_n997), .A3(new_n982), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1019), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(G290), .B(G1986), .Z(new_n1111));
  OAI211_X1 g686(.A(new_n948), .B(new_n954), .C1(new_n941), .C2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n965), .B1(new_n1110), .B2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g688(.A1(G227), .A2(G401), .ZN(new_n1115));
  NAND3_X1  g689(.A1(new_n1115), .A2(G319), .A3(new_n672), .ZN(new_n1116));
  XNOR2_X1  g690(.A(new_n1116), .B(KEYINPUT127), .ZN(new_n1117));
  AND3_X1   g691(.A1(new_n864), .A2(new_n920), .A3(new_n1117), .ZN(G308));
  NAND3_X1  g692(.A1(new_n864), .A2(new_n920), .A3(new_n1117), .ZN(G225));
endmodule


