

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(G8), .A2(n725), .ZN(n772) );
  BUF_X1 U551 ( .A(n548), .Z(n549) );
  INV_X1 U552 ( .A(n517), .ZN(n522) );
  XNOR2_X1 U553 ( .A(KEYINPUT64), .B(G2104), .ZN(n517) );
  NOR2_X1 U554 ( .A1(n759), .A2(n758), .ZN(n760) );
  INV_X1 U555 ( .A(KEYINPUT85), .ZN(n518) );
  NOR2_X2 U556 ( .A1(n536), .A2(n535), .ZN(G160) );
  NOR2_X1 U557 ( .A1(n772), .A2(n753), .ZN(n515) );
  INV_X1 U558 ( .A(KEYINPUT30), .ZN(n727) );
  XNOR2_X1 U559 ( .A(n734), .B(KEYINPUT31), .ZN(n742) );
  AND2_X1 U560 ( .A1(n522), .A2(G2105), .ZN(n532) );
  NOR2_X1 U561 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n649) );
  BUF_X1 U563 ( .A(n532), .Z(n889) );
  XNOR2_X1 U564 ( .A(n519), .B(n518), .ZN(n520) );
  NOR2_X1 U565 ( .A1(n526), .A2(n525), .ZN(G164) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n516), .Z(n548) );
  NAND2_X1 U568 ( .A1(n548), .A2(G138), .ZN(n521) );
  NAND2_X1 U569 ( .A1(G126), .A2(n532), .ZN(n519) );
  NAND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n526) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n890) );
  NAND2_X1 U572 ( .A1(G114), .A2(n890), .ZN(n524) );
  NOR2_X4 U573 ( .A1(n522), .A2(G2105), .ZN(n528) );
  NAND2_X1 U574 ( .A1(G102), .A2(n528), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U576 ( .A1(G137), .A2(n548), .ZN(n527) );
  XOR2_X1 U577 ( .A(n527), .B(KEYINPUT65), .Z(n531) );
  NAND2_X1 U578 ( .A1(G101), .A2(n528), .ZN(n529) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n536) );
  NAND2_X1 U581 ( .A1(G125), .A2(n889), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G113), .A2(n890), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U584 ( .A(G2438), .B(G2454), .Z(n538) );
  XNOR2_X1 U585 ( .A(G2435), .B(G2430), .ZN(n537) );
  XNOR2_X1 U586 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U587 ( .A(n539), .B(G2427), .Z(n541) );
  XNOR2_X1 U588 ( .A(G1341), .B(G1348), .ZN(n540) );
  XNOR2_X1 U589 ( .A(n541), .B(n540), .ZN(n545) );
  XOR2_X1 U590 ( .A(G2443), .B(G2446), .Z(n543) );
  XNOR2_X1 U591 ( .A(KEYINPUT106), .B(G2451), .ZN(n542) );
  XNOR2_X1 U592 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U593 ( .A(n545), .B(n544), .Z(n546) );
  AND2_X1 U594 ( .A1(G14), .A2(n546), .ZN(G401) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(G123), .A2(n889), .ZN(n547) );
  XNOR2_X1 U597 ( .A(n547), .B(KEYINPUT18), .ZN(n556) );
  NAND2_X1 U598 ( .A1(G135), .A2(n549), .ZN(n551) );
  NAND2_X1 U599 ( .A1(G111), .A2(n890), .ZN(n550) );
  NAND2_X1 U600 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U601 ( .A1(n528), .A2(G99), .ZN(n552) );
  XOR2_X1 U602 ( .A(KEYINPUT74), .B(n552), .Z(n553) );
  NOR2_X1 U603 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U604 ( .A1(n556), .A2(n555), .ZN(n926) );
  XNOR2_X1 U605 ( .A(G2096), .B(n926), .ZN(n557) );
  OR2_X1 U606 ( .A1(G2100), .A2(n557), .ZN(G156) );
  INV_X1 U607 ( .A(G132), .ZN(G219) );
  INV_X1 U608 ( .A(G82), .ZN(G220) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  INV_X1 U610 ( .A(G651), .ZN(n561) );
  NOR2_X1 U611 ( .A1(G543), .A2(n561), .ZN(n558) );
  XOR2_X1 U612 ( .A(KEYINPUT1), .B(n558), .Z(n650) );
  NAND2_X1 U613 ( .A1(G65), .A2(n650), .ZN(n560) );
  XOR2_X1 U614 ( .A(KEYINPUT0), .B(G543), .Z(n627) );
  NOR2_X2 U615 ( .A1(G651), .A2(n627), .ZN(n657) );
  NAND2_X1 U616 ( .A1(G53), .A2(n657), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U618 ( .A1(G91), .A2(n649), .ZN(n563) );
  NOR2_X1 U619 ( .A1(n627), .A2(n561), .ZN(n653) );
  NAND2_X1 U620 ( .A1(G78), .A2(n653), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n707) );
  INV_X1 U623 ( .A(n707), .ZN(G299) );
  NAND2_X1 U624 ( .A1(G64), .A2(n650), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G52), .A2(n657), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G90), .A2(n649), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G77), .A2(n653), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U631 ( .A1(n572), .A2(n571), .ZN(G171) );
  NAND2_X1 U632 ( .A1(n649), .A2(G89), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G76), .A2(n653), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U636 ( .A(KEYINPUT5), .B(n576), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G63), .A2(n650), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G51), .A2(n657), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT72), .B(KEYINPUT6), .Z(n579) );
  XNOR2_X1 U641 ( .A(n580), .B(n579), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U643 ( .A(KEYINPUT7), .B(n583), .ZN(G168) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n584) );
  XOR2_X1 U646 ( .A(n584), .B(KEYINPUT10), .Z(n829) );
  NAND2_X1 U647 ( .A1(n829), .A2(G567), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  XOR2_X1 U649 ( .A(G860), .B(KEYINPUT68), .Z(n611) );
  NAND2_X1 U650 ( .A1(G56), .A2(n650), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n586), .Z(n592) );
  NAND2_X1 U652 ( .A1(n649), .A2(G81), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G68), .A2(n653), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U656 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U658 ( .A1(n657), .A2(G43), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n967) );
  OR2_X1 U660 ( .A1(n611), .A2(n967), .ZN(G153) );
  INV_X1 U661 ( .A(G171), .ZN(G301) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U663 ( .A1(n657), .A2(G54), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT70), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n653), .A2(G79), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT71), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G66), .A2(n650), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G92), .A2(n649), .ZN(n601) );
  XNOR2_X1 U671 ( .A(KEYINPUT69), .B(n601), .ZN(n602) );
  XOR2_X1 U672 ( .A(KEYINPUT15), .B(n604), .Z(n979) );
  INV_X1 U673 ( .A(n979), .ZN(n840) );
  INV_X1 U674 ( .A(G868), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n840), .A2(n607), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(G284) );
  NOR2_X1 U677 ( .A1(G286), .A2(n607), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT73), .B(n608), .Z(n610) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U681 ( .A1(n611), .A2(G559), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n612), .A2(n979), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n967), .ZN(n616) );
  NAND2_X1 U685 ( .A1(G868), .A2(n979), .ZN(n614) );
  NOR2_X1 U686 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U687 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U688 ( .A1(n653), .A2(G80), .ZN(n617) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT76), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G67), .A2(n650), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U692 ( .A1(G93), .A2(n649), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G55), .A2(n657), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n661) );
  NAND2_X1 U696 ( .A1(G559), .A2(n979), .ZN(n624) );
  XNOR2_X1 U697 ( .A(n967), .B(n624), .ZN(n667) );
  NOR2_X1 U698 ( .A1(G860), .A2(n667), .ZN(n625) );
  XOR2_X1 U699 ( .A(KEYINPUT75), .B(n625), .Z(n626) );
  XNOR2_X1 U700 ( .A(n661), .B(n626), .ZN(G145) );
  NAND2_X1 U701 ( .A1(G49), .A2(n657), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G87), .A2(n627), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n650), .A2(n630), .ZN(n632) );
  NAND2_X1 U705 ( .A1(G651), .A2(G74), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U707 ( .A1(G88), .A2(n649), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G75), .A2(n653), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n640) );
  NAND2_X1 U710 ( .A1(G50), .A2(n657), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT78), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G62), .A2(n650), .ZN(n636) );
  XOR2_X1 U713 ( .A(KEYINPUT77), .B(n636), .Z(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(G166) );
  INV_X1 U716 ( .A(G166), .ZN(G303) );
  NAND2_X1 U717 ( .A1(G85), .A2(n649), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G72), .A2(n653), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U720 ( .A(KEYINPUT66), .B(n643), .ZN(n646) );
  NAND2_X1 U721 ( .A1(G60), .A2(n650), .ZN(n644) );
  XNOR2_X1 U722 ( .A(KEYINPUT67), .B(n644), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n657), .A2(G47), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(G290) );
  NAND2_X1 U726 ( .A1(G86), .A2(n649), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G61), .A2(n650), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n657), .A2(G48), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(G305) );
  NOR2_X1 U734 ( .A1(G868), .A2(n661), .ZN(n660) );
  XOR2_X1 U735 ( .A(KEYINPUT80), .B(n660), .Z(n671) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(G288), .ZN(n666) );
  XOR2_X1 U737 ( .A(G303), .B(G290), .Z(n662) );
  XOR2_X1 U738 ( .A(n662), .B(n661), .Z(n663) );
  XOR2_X1 U739 ( .A(G299), .B(n663), .Z(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(G305), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n666), .B(n665), .ZN(n838) );
  XOR2_X1 U742 ( .A(n838), .B(n667), .Z(n668) );
  NAND2_X1 U743 ( .A1(n668), .A2(G868), .ZN(n669) );
  XOR2_X1 U744 ( .A(KEYINPUT79), .B(n669), .Z(n670) );
  NAND2_X1 U745 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n675), .A2(G2072), .ZN(n676) );
  XOR2_X1 U751 ( .A(KEYINPUT81), .B(n676), .Z(G158) );
  XNOR2_X1 U752 ( .A(KEYINPUT82), .B(G44), .ZN(n677) );
  XNOR2_X1 U753 ( .A(n677), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U755 ( .A1(G237), .A2(n678), .ZN(n679) );
  XNOR2_X1 U756 ( .A(KEYINPUT84), .B(n679), .ZN(n680) );
  NAND2_X1 U757 ( .A1(n680), .A2(G108), .ZN(n835) );
  NAND2_X1 U758 ( .A1(n835), .A2(G567), .ZN(n686) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n681) );
  XNOR2_X1 U760 ( .A(KEYINPUT22), .B(n681), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n682), .A2(G96), .ZN(n683) );
  NOR2_X1 U762 ( .A1(n683), .A2(G218), .ZN(n684) );
  XNOR2_X1 U763 ( .A(n684), .B(KEYINPUT83), .ZN(n834) );
  NAND2_X1 U764 ( .A1(n834), .A2(G2106), .ZN(n685) );
  NAND2_X1 U765 ( .A1(n686), .A2(n685), .ZN(n912) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U767 ( .A1(n912), .A2(n687), .ZN(n831) );
  NAND2_X1 U768 ( .A1(n831), .A2(G36), .ZN(G176) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n776) );
  INV_X1 U770 ( .A(n776), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n775) );
  NOR2_X2 U772 ( .A1(n688), .A2(n775), .ZN(n714) );
  INV_X2 U773 ( .A(n714), .ZN(n725) );
  NAND2_X1 U774 ( .A1(G1348), .A2(n725), .ZN(n690) );
  NAND2_X1 U775 ( .A1(G2067), .A2(n714), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n697) );
  NOR2_X1 U777 ( .A1(n840), .A2(n697), .ZN(n696) );
  INV_X1 U778 ( .A(G1996), .ZN(n847) );
  NOR2_X1 U779 ( .A1(n725), .A2(n847), .ZN(n691) );
  XOR2_X1 U780 ( .A(n691), .B(KEYINPUT26), .Z(n693) );
  NAND2_X1 U781 ( .A1(n725), .A2(G1341), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n967), .A2(n694), .ZN(n695) );
  OR2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U785 ( .A1(n840), .A2(n697), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U787 ( .A1(G1956), .A2(n725), .ZN(n700) );
  XNOR2_X1 U788 ( .A(KEYINPUT95), .B(n700), .ZN(n703) );
  NAND2_X1 U789 ( .A1(n714), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U790 ( .A(KEYINPUT27), .B(n701), .ZN(n702) );
  NOR2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U792 ( .A1(n707), .A2(n706), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U795 ( .A(n708), .B(KEYINPUT28), .Z(n709) );
  NAND2_X1 U796 ( .A1(n710), .A2(n709), .ZN(n712) );
  XOR2_X1 U797 ( .A(KEYINPUT29), .B(KEYINPUT96), .Z(n711) );
  XNOR2_X1 U798 ( .A(n712), .B(n711), .ZN(n718) );
  XOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .Z(n713) );
  XNOR2_X1 U800 ( .A(KEYINPUT94), .B(n713), .ZN(n944) );
  NOR2_X1 U801 ( .A1(n725), .A2(n944), .ZN(n716) );
  XOR2_X1 U802 ( .A(G1961), .B(KEYINPUT93), .Z(n996) );
  NOR2_X1 U803 ( .A1(n714), .A2(n996), .ZN(n715) );
  NOR2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n731) );
  OR2_X1 U805 ( .A1(n731), .A2(G301), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n741) );
  INV_X1 U807 ( .A(G8), .ZN(n724) );
  NOR2_X1 U808 ( .A1(G1971), .A2(n772), .ZN(n720) );
  NOR2_X1 U809 ( .A1(G2090), .A2(n725), .ZN(n719) );
  NOR2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U811 ( .A1(n721), .A2(G303), .ZN(n722) );
  XNOR2_X1 U812 ( .A(n722), .B(KEYINPUT98), .ZN(n723) );
  OR2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n736) );
  AND2_X1 U814 ( .A1(n741), .A2(n736), .ZN(n735) );
  NOR2_X1 U815 ( .A1(G1966), .A2(n772), .ZN(n744) );
  NOR2_X1 U816 ( .A1(G2084), .A2(n725), .ZN(n745) );
  NOR2_X1 U817 ( .A1(n744), .A2(n745), .ZN(n726) );
  AND2_X1 U818 ( .A1(n726), .A2(G8), .ZN(n728) );
  XNOR2_X1 U819 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U820 ( .A1(G168), .A2(n729), .ZN(n730) );
  XNOR2_X1 U821 ( .A(n730), .B(KEYINPUT97), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n731), .A2(G301), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U824 ( .A1(n735), .A2(n742), .ZN(n739) );
  INV_X1 U825 ( .A(n736), .ZN(n737) );
  OR2_X1 U826 ( .A1(n737), .A2(G286), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U828 ( .A(n740), .B(KEYINPUT32), .ZN(n749) );
  AND2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U831 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n763) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U836 ( .A1(n756), .A2(n750), .ZN(n971) );
  XOR2_X1 U837 ( .A(n971), .B(KEYINPUT99), .Z(n751) );
  NAND2_X1 U838 ( .A1(n763), .A2(n751), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT100), .ZN(n754) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n970) );
  INV_X1 U841 ( .A(n970), .ZN(n753) );
  AND2_X1 U842 ( .A1(n754), .A2(n515), .ZN(n755) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n755), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n772), .A2(n757), .ZN(n758) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n964) );
  NAND2_X1 U847 ( .A1(n760), .A2(n964), .ZN(n767) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n761) );
  XOR2_X1 U849 ( .A(KEYINPUT101), .B(n761), .Z(n762) );
  NAND2_X1 U850 ( .A1(G8), .A2(n762), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U852 ( .A1(n765), .A2(n772), .ZN(n766) );
  NAND2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U854 ( .A(n768), .B(KEYINPUT102), .ZN(n774) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U856 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  XNOR2_X1 U857 ( .A(KEYINPUT92), .B(n770), .ZN(n771) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n807) );
  NOR2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U861 ( .A(KEYINPUT87), .B(n777), .Z(n823) );
  XNOR2_X1 U862 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NAND2_X1 U863 ( .A1(G128), .A2(n889), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G116), .A2(n890), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n781) );
  XOR2_X1 U866 ( .A(KEYINPUT35), .B(KEYINPUT90), .Z(n780) );
  XNOR2_X1 U867 ( .A(n781), .B(n780), .ZN(n788) );
  XNOR2_X1 U868 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(KEYINPUT34), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G140), .A2(n549), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G104), .A2(n528), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U873 ( .A(n786), .B(n785), .Z(n787) );
  NOR2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U875 ( .A(KEYINPUT36), .B(n789), .ZN(n900) );
  NOR2_X1 U876 ( .A1(n820), .A2(n900), .ZN(n929) );
  NAND2_X1 U877 ( .A1(n823), .A2(n929), .ZN(n818) );
  NAND2_X1 U878 ( .A1(G141), .A2(n549), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G117), .A2(n890), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n528), .A2(G105), .ZN(n792) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n792), .Z(n793) );
  NOR2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n889), .A2(G129), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n901) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n901), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G119), .A2(n889), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G107), .A2(n890), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G131), .A2(n549), .ZN(n800) );
  NAND2_X1 U891 ( .A1(G95), .A2(n528), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n875) );
  NAND2_X1 U894 ( .A1(G1991), .A2(n875), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n921) );
  NAND2_X1 U896 ( .A1(n823), .A2(n921), .ZN(n805) );
  XOR2_X1 U897 ( .A(KEYINPUT91), .B(n805), .Z(n811) );
  NAND2_X1 U898 ( .A1(n818), .A2(n811), .ZN(n806) );
  NOR2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n810) );
  XNOR2_X1 U900 ( .A(G1986), .B(KEYINPUT86), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(G290), .ZN(n969) );
  NAND2_X1 U902 ( .A1(n969), .A2(n823), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n826) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n901), .ZN(n919) );
  INV_X1 U905 ( .A(n811), .ZN(n815) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n875), .ZN(n812) );
  XOR2_X1 U907 ( .A(KEYINPUT103), .B(n812), .Z(n925) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n925), .A2(n813), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n919), .A2(n816), .ZN(n817) );
  XNOR2_X1 U912 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n820), .A2(n900), .ZN(n922) );
  NAND2_X1 U915 ( .A1(n821), .A2(n922), .ZN(n822) );
  XNOR2_X1 U916 ( .A(KEYINPUT104), .B(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n827) );
  XNOR2_X1 U920 ( .A(n828), .B(n827), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U922 ( .A(n829), .ZN(G223) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U927 ( .A(KEYINPUT107), .B(n833), .Z(G188) );
  XOR2_X1 U928 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n836), .B(KEYINPUT108), .Z(G261) );
  INV_X1 U935 ( .A(G261), .ZN(G325) );
  XOR2_X1 U936 ( .A(KEYINPUT116), .B(G171), .Z(n837) );
  XNOR2_X1 U937 ( .A(n837), .B(n967), .ZN(n839) );
  XOR2_X1 U938 ( .A(n839), .B(n838), .Z(n842) );
  XOR2_X1 U939 ( .A(n840), .B(G286), .Z(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  NOR2_X1 U941 ( .A1(G37), .A2(n843), .ZN(G397) );
  XOR2_X1 U942 ( .A(G2474), .B(G1956), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1981), .B(G1966), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n846), .B(KEYINPUT112), .Z(n849) );
  XOR2_X1 U946 ( .A(n847), .B(G1991), .Z(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U948 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1961), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U952 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(G229) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2084), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n856), .B(KEYINPUT109), .ZN(n866) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2678), .Z(n858) );
  XNOR2_X1 U957 ( .A(KEYINPUT110), .B(G2096), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U959 ( .A(G2100), .B(G2072), .Z(n860) );
  XNOR2_X1 U960 ( .A(G2090), .B(G2078), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n889), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n867), .B(KEYINPUT114), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G112), .A2(n890), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G136), .A2(n549), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G100), .A2(n528), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(G162) );
  XNOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n875), .B(KEYINPUT46), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U978 ( .A(G160), .B(n878), .ZN(n899) );
  NAND2_X1 U979 ( .A1(G130), .A2(n889), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G118), .A2(n890), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G142), .A2(n549), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G106), .A2(n528), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U985 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U987 ( .A(G162), .B(n886), .ZN(n897) );
  NAND2_X1 U988 ( .A1(G139), .A2(n549), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G103), .A2(n528), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G127), .A2(n889), .ZN(n892) );
  NAND2_X1 U992 ( .A1(G115), .A2(n890), .ZN(n891) );
  NAND2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n913) );
  XNOR2_X1 U996 ( .A(n926), .B(n913), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n904) );
  XNOR2_X1 U999 ( .A(G164), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G395) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G397), .A2(n907), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n912), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT117), .B(n908), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G395), .A2(n909), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(n912), .ZN(G319) );
  XNOR2_X1 U1012 ( .A(G164), .B(G2078), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(G2072), .B(n913), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(KEYINPUT120), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n917), .B(KEYINPUT50), .ZN(n936) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n920), .Z(n934) );
  INV_X1 U1020 ( .A(n921), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n932) );
  XOR2_X1 U1022 ( .A(G160), .B(G2084), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(KEYINPUT119), .B(n930), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n937), .ZN(n939) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(G29), .ZN(n1019) );
  XOR2_X1 U1034 ( .A(G32), .B(G1996), .Z(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1036 ( .A(G1991), .B(G25), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G2072), .B(G33), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(n944), .B(G27), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1044 ( .A(n951), .B(KEYINPUT121), .Z(n952) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G35), .B(G2090), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT122), .B(n955), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(KEYINPUT54), .B(G34), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(n956), .B(KEYINPUT123), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G2084), .B(n957), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1053 ( .A(KEYINPUT55), .B(n960), .Z(n962) );
  INV_X1 U1054 ( .A(G29), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n963), .ZN(n1017) );
  INV_X1 U1057 ( .A(G16), .ZN(n1013) );
  XOR2_X1 U1058 ( .A(n1013), .B(KEYINPUT56), .Z(n988) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT57), .ZN(n986) );
  XNOR2_X1 U1062 ( .A(G1341), .B(n967), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n978) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n975) );
  XOR2_X1 U1065 ( .A(G1956), .B(G299), .Z(n973) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT125), .B(n976), .Z(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n984) );
  XOR2_X1 U1071 ( .A(G171), .B(G1961), .Z(n981) );
  XOR2_X1 U1072 ( .A(n979), .B(G1348), .Z(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(KEYINPUT124), .B(n982), .Z(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n1015) );
  XOR2_X1 U1078 ( .A(G1971), .B(KEYINPUT126), .Z(n989) );
  XNOR2_X1 U1079 ( .A(G22), .B(n989), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(G23), .B(G1976), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT58), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(KEYINPUT127), .B(n995), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G21), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n996), .B(G5), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1010) );
  XOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .Z(n1001) );
  XNOR2_X1 U1091 ( .A(G4), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G20), .B(G1956), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1020), .ZN(G150) );
  INV_X1 U1106 ( .A(G150), .ZN(G311) );
endmodule

