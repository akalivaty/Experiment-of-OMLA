//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1052, new_n1053, new_n1054;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT26), .ZN(new_n204));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n203), .A2(KEYINPUT26), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT28), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(KEYINPUT28), .A3(new_n211), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n220), .A2(new_n222), .A3(new_n207), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n223), .A2(new_n228), .A3(KEYINPUT65), .A4(KEYINPUT25), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT25), .A4(new_n207), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n226), .B(new_n227), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n223), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n234), .A2(new_n235), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n235), .B1(new_n234), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n217), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(G113gat), .B2(G120gat), .ZN(new_n248));
  AND2_X1   g047(.A1(G113gat), .A2(G120gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G127gat), .B(G134gat), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(new_n246), .C1(new_n249), .C2(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G227gat), .ZN(new_n257));
  INV_X1    g056(.A(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n252), .A2(new_n254), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n260), .B(new_n217), .C1(new_n243), .C2(new_n244), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n256), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT33), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G15gat), .B(G43gat), .Z(new_n265));
  XNOR2_X1  g064(.A(G71gat), .B(G99gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n256), .A2(new_n261), .ZN(new_n269));
  INV_X1    g068(.A(new_n259), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT34), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT34), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n262), .A2(KEYINPUT32), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n267), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(new_n262), .B2(new_n263), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n273), .B1(new_n269), .B2(new_n270), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT34), .B(new_n259), .C1(new_n256), .C2(new_n261), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n275), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(G211gat), .A2(G218gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(G211gat), .A2(G218gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g087(.A1(G197gat), .A2(G204gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G197gat), .A2(G204gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n292), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT3), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT71), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G148gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n304), .A3(G141gat), .ZN(new_n305));
  INV_X1    g104(.A(G141gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n301), .A2(G141gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n310), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n312), .A2(new_n309), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n308), .A2(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n285), .B1(new_n300), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321));
  XNOR2_X1  g120(.A(G141gat), .B(G148gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n318), .B1(new_n322), .B2(KEYINPUT2), .ZN(new_n323));
  INV_X1    g122(.A(new_n307), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT71), .B(G148gat), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n324), .B1(new_n325), .B2(G141gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n312), .B1(new_n310), .B2(new_n309), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n321), .B(new_n323), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n298), .B1(new_n328), .B2(new_n299), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT77), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n294), .A2(new_n295), .A3(new_n332), .A4(new_n296), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n299), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT78), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n293), .A2(new_n297), .A3(KEYINPUT77), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n299), .A4(new_n333), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n321), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n329), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n330), .B1(new_n343), .B2(new_n284), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT79), .ZN(new_n345));
  INV_X1    g144(.A(G22gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n330), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n329), .B1(new_n339), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n285), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT31), .B(G50gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  AOI21_X1  g153(.A(new_n346), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n354), .ZN(new_n356));
  AOI211_X1 g155(.A(G22gat), .B(new_n356), .C1(new_n349), .C2(new_n350), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n345), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n299), .A3(new_n333), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n359), .B2(KEYINPUT78), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n319), .B1(new_n360), .B2(new_n338), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n284), .B1(new_n361), .B2(new_n329), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT79), .B1(new_n362), .B2(new_n347), .ZN(new_n363));
  OAI21_X1  g162(.A(G22gat), .B1(new_n363), .B2(new_n356), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n351), .A2(new_n346), .A3(new_n354), .ZN(new_n365));
  INV_X1    g164(.A(new_n345), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n358), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n277), .B1(new_n275), .B2(new_n282), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n283), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n371));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(new_n217), .C1(new_n243), .C2(new_n244), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n234), .A2(new_n242), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n299), .B(new_n372), .C1(new_n375), .C2(new_n216), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n298), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT69), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n298), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n373), .B1(new_n245), .B2(new_n299), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT68), .B(new_n373), .C1(new_n375), .C2(new_n216), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT68), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n216), .B1(new_n234), .B2(new_n242), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n372), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n381), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n381), .B1(new_n374), .B2(new_n376), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT69), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND4_X1  g192(.A1(new_n380), .A2(new_n388), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n234), .A2(new_n242), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT66), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n234), .A2(new_n235), .A3(new_n242), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n216), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n372), .B1(new_n400), .B2(KEYINPUT29), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n383), .A2(new_n386), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n403), .A2(new_n381), .B1(KEYINPUT69), .B2(new_n389), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n393), .B1(new_n404), .B2(new_n380), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n404), .A2(KEYINPUT70), .A3(new_n380), .A4(new_n393), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n394), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n409), .A3(new_n395), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT35), .ZN(new_n412));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT0), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT76), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT4), .B1(new_n319), .B2(new_n255), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT73), .B1(new_n260), .B2(new_n340), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT73), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n319), .A2(new_n255), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n423), .B2(KEYINPUT4), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n305), .A2(new_n307), .B1(new_n313), .B2(new_n311), .ZN(new_n425));
  XNOR2_X1  g224(.A(G155gat), .B(G162gat), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n310), .B2(new_n316), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n260), .A3(new_n328), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n430), .B(KEYINPUT72), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n418), .B1(new_n424), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n420), .B2(new_n422), .ZN(new_n438));
  NOR4_X1   g237(.A1(new_n438), .A2(new_n434), .A3(KEYINPUT76), .A4(new_n419), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n433), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n319), .A2(new_n421), .A3(new_n255), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n421), .B1(new_n319), .B2(new_n255), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n319), .A2(new_n255), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n445), .B2(new_n432), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n420), .A2(new_n437), .A3(new_n422), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n319), .A2(new_n255), .A3(KEYINPUT4), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n432), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n447), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT74), .A3(new_n448), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n446), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n417), .B1(new_n440), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n420), .B(new_n422), .C1(new_n255), .C2(new_n319), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n433), .B1(new_n458), .B2(new_n431), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n449), .A2(new_n447), .A3(new_n451), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT74), .B1(new_n453), .B2(new_n448), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT4), .B1(new_n442), .B2(new_n443), .ZN(new_n463));
  INV_X1    g262(.A(new_n419), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT76), .B1(new_n465), .B2(new_n434), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n424), .A2(new_n435), .A3(new_n418), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(new_n468), .A3(new_n416), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n456), .A2(new_n457), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT6), .B(new_n417), .C1(new_n440), .C2(new_n455), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n412), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n370), .A2(new_n371), .A3(new_n411), .A4(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n366), .B1(new_n364), .B2(new_n365), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n282), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n276), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n275), .A2(new_n277), .A3(new_n282), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n476), .A2(new_n479), .A3(new_n472), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n406), .A2(new_n410), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT81), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n470), .A2(new_n471), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n283), .A2(new_n369), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n411), .A2(new_n484), .A3(new_n485), .A4(new_n476), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n473), .A2(new_n483), .B1(new_n486), .B2(KEYINPUT35), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n283), .B2(new_n369), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(KEYINPUT36), .A3(new_n480), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n406), .A2(new_n410), .A3(new_n484), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n489), .A2(new_n490), .B1(new_n491), .B2(new_n368), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT39), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n458), .A2(new_n431), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n424), .A2(new_n429), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n494), .B(new_n495), .C1(new_n496), .C2(new_n431), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n494), .A3(new_n431), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n416), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n456), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n497), .A2(new_n499), .A3(new_n493), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n482), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n393), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n380), .A2(new_n388), .A3(new_n390), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(KEYINPUT37), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n404), .B2(new_n380), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT38), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n407), .A2(new_n409), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n470), .A2(new_n471), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n403), .A2(new_n298), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n377), .B2(new_n381), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT38), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(new_n505), .C1(KEYINPUT37), .C2(new_n506), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n504), .A2(new_n517), .A3(new_n476), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n492), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n202), .B1(new_n487), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n485), .A2(new_n476), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT35), .B1(new_n521), .B2(new_n491), .ZN(new_n522));
  AND4_X1   g321(.A1(new_n476), .A2(new_n479), .A3(new_n472), .A4(new_n480), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n371), .B1(new_n523), .B2(new_n411), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n481), .A2(KEYINPUT81), .A3(new_n482), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n492), .A2(new_n518), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT82), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n346), .A2(G15gat), .ZN(new_n532));
  INV_X1    g331(.A(G15gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G22gat), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT85), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT85), .B1(new_n532), .B2(new_n534), .ZN(new_n536));
  OAI221_X1 g335(.A(KEYINPUT87), .B1(new_n531), .B2(G1gat), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G8gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT85), .ZN(new_n540));
  INV_X1    g339(.A(G1gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  OAI22_X1  g342(.A1(new_n535), .A2(new_n536), .B1(new_n531), .B2(G1gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n530), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n542), .A2(new_n538), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n545), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n549), .A4(new_n537), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n542), .A2(KEYINPUT86), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n538), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT86), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT14), .B(G29gat), .ZN(new_n556));
  INV_X1    g355(.A(G36gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G29gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G43gat), .B(G50gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G43gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT83), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G43gat), .ZN(new_n569));
  INV_X1    g368(.A(G50gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n558), .A2(new_n560), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n565), .B(KEYINPUT84), .C1(new_n564), .C2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n558), .A2(new_n560), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n571), .A2(new_n572), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n563), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n579), .A2(KEYINPUT84), .A3(KEYINPUT17), .A4(new_n565), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n551), .A2(new_n555), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n565), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n547), .A2(new_n550), .B1(new_n554), .B2(new_n553), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT18), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n583), .B(KEYINPUT13), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n551), .A2(new_n555), .ZN(new_n590));
  INV_X1    g389(.A(new_n584), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n585), .A2(new_n584), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n591), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(KEYINPUT18), .A3(new_n583), .A4(new_n582), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G197gat), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT11), .B(G169gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n588), .A2(new_n594), .A3(new_n602), .A4(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G57gat), .B(G64gat), .Z(new_n607));
  INV_X1    g406(.A(G71gat), .ZN(new_n608));
  INV_X1    g407(.A(G78gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT9), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n607), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G57gat), .B(G64gat), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n611), .B(new_n610), .C1(new_n616), .C2(new_n613), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G127gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n590), .B1(KEYINPUT21), .B2(new_n618), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  INV_X1    g424(.A(G155gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G183gat), .B(G211gat), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n624), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT8), .ZN(new_n636));
  NAND2_X1  g435(.A1(G99gat), .A2(G106gat), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(KEYINPUT92), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(KEYINPUT92), .B2(new_n637), .ZN(new_n639));
  XNOR2_X1  g438(.A(G99gat), .B(G106gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n641), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(G85gat), .A3(G92gat), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n639), .A2(new_n640), .A3(new_n642), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT93), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n645), .A2(new_n642), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n648), .B2(new_n639), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AOI211_X1 g449(.A(KEYINPUT93), .B(new_n640), .C1(new_n648), .C2(new_n639), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n635), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n639), .A2(new_n642), .A3(new_n645), .ZN(new_n653));
  INV_X1    g452(.A(new_n640), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(KEYINPUT93), .A3(new_n646), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n647), .A2(new_n649), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT94), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n581), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n652), .A2(new_n591), .A3(new_n658), .ZN(new_n661));
  XNOR2_X1  g460(.A(G190gat), .B(G218gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G232gat), .A2(G233gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT89), .Z(new_n665));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n660), .A2(new_n661), .A3(new_n663), .A4(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT95), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(G134gat), .B(G162gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT90), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n666), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n660), .A2(new_n661), .A3(new_n667), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n662), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n670), .A2(new_n674), .B1(new_n676), .B2(new_n668), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n676), .A2(KEYINPUT95), .A3(new_n668), .A4(new_n674), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n652), .A2(KEYINPUT10), .A3(new_n658), .A4(new_n618), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n615), .A2(new_n617), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n656), .A2(new_n657), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT10), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n649), .A2(new_n682), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n646), .ZN(new_n687));
  AND4_X1   g486(.A1(new_n685), .A2(new_n655), .A3(new_n618), .A4(new_n646), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n683), .B(new_n684), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(G230gat), .A2(G233gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n693));
  INV_X1    g492(.A(new_n691), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(G120gat), .B(G148gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(G176gat), .B(G204gat), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n697), .B(new_n698), .Z(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n692), .A2(new_n695), .A3(new_n699), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n634), .A2(new_n680), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n529), .A2(new_n606), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n484), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT97), .B(G1gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1324gat));
  INV_X1    g507(.A(new_n705), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT98), .B(KEYINPUT16), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n538), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n709), .A2(new_n482), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n538), .B1(new_n709), .B2(new_n482), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT42), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(KEYINPUT42), .B2(new_n712), .ZN(G1325gat));
  INV_X1    g514(.A(new_n489), .ZN(new_n716));
  INV_X1    g515(.A(new_n490), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G15gat), .B1(new_n705), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n485), .A2(new_n533), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n720), .B1(new_n705), .B2(new_n721), .ZN(G1326gat));
  NOR2_X1   g521(.A1(new_n705), .A2(new_n476), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT43), .B(G22gat), .Z(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1327gat));
  INV_X1    g524(.A(new_n680), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n633), .A2(new_n726), .A3(new_n703), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n520), .A2(new_n528), .A3(new_n606), .A4(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(G29gat), .A3(new_n484), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT45), .Z(new_n730));
  NAND3_X1  g529(.A1(new_n520), .A2(new_n528), .A3(new_n680), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n473), .A2(new_n483), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n733), .A2(KEYINPUT101), .A3(new_n522), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT101), .B1(new_n733), .B2(new_n522), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n527), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n678), .A2(KEYINPUT102), .A3(new_n679), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n738));
  INV_X1    g537(.A(new_n679), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n677), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n732), .A2(new_n744), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n604), .A2(KEYINPUT99), .A3(new_n605), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT99), .B1(new_n604), .B2(new_n605), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n703), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n634), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT100), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n745), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT103), .B1(new_n754), .B2(new_n484), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G29gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n754), .A2(KEYINPUT103), .A3(new_n484), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n730), .B1(new_n756), .B2(new_n757), .ZN(G1328gat));
  NOR3_X1   g557(.A1(new_n728), .A2(G36gat), .A3(new_n411), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n752), .B1(new_n732), .B2(new_n744), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n557), .B1(new_n762), .B2(new_n482), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT104), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n759), .B(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g564(.A(G36gat), .B1(new_n754), .B2(new_n411), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(G1329gat));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n770));
  AOI211_X1 g569(.A(new_n719), .B(new_n752), .C1(new_n732), .C2(new_n744), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n567), .A2(new_n569), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n485), .A2(new_n772), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n728), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n771), .B2(new_n772), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n773), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI221_X1 g577(.A(new_n775), .B1(new_n770), .B2(KEYINPUT47), .C1(new_n771), .C2(new_n772), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1330gat));
  AOI21_X1  g579(.A(new_n570), .B1(new_n762), .B2(new_n368), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT48), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n368), .A2(new_n570), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT106), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n728), .A2(new_n784), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n781), .A2(new_n782), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n782), .B1(new_n781), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1331gat));
  NAND4_X1  g587(.A1(new_n748), .A2(new_n726), .A3(new_n633), .A4(new_n703), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT107), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n736), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n512), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n411), .ZN(new_n795));
  NOR2_X1   g594(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n796));
  AND2_X1   g595(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n795), .B2(new_n796), .ZN(G1333gat));
  INV_X1    g598(.A(new_n485), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n791), .A2(KEYINPUT108), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT108), .B1(new_n791), .B2(new_n800), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n608), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n792), .A2(G71gat), .A3(new_n718), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT50), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1334gat));
  NOR2_X1   g608(.A1(new_n791), .A2(new_n476), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(new_n609), .ZN(G1335gat));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT101), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n526), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n487), .A2(KEYINPUT101), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n519), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n748), .A2(new_n634), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n726), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n812), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n736), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(G85gat), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n512), .A4(new_n703), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n817), .A2(new_n750), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n732), .B2(new_n744), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n512), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n824), .B1(new_n828), .B2(new_n823), .ZN(G1336gat));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n482), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n411), .A2(G92gat), .A3(new_n750), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n832), .B(KEYINPUT109), .Z(new_n833));
  AOI22_X1  g632(.A1(new_n831), .A2(G92gat), .B1(new_n822), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n831), .A2(G92gat), .ZN(new_n835));
  INV_X1    g634(.A(new_n822), .ZN(new_n836));
  INV_X1    g635(.A(new_n832), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n830), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n830), .A2(new_n834), .B1(new_n835), .B2(new_n838), .ZN(G1337gat));
  AND2_X1   g638(.A1(new_n827), .A2(new_n718), .ZN(new_n840));
  INV_X1    g639(.A(G99gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n485), .A2(new_n841), .A3(new_n703), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n840), .A2(new_n841), .B1(new_n836), .B2(new_n842), .ZN(G1338gat));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n476), .A2(new_n750), .ZN(new_n845));
  AOI21_X1  g644(.A(G106gat), .B1(new_n822), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n368), .A2(G106gat), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n826), .B(new_n847), .C1(new_n732), .C2(new_n744), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n844), .B(KEYINPUT53), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n816), .A2(new_n812), .A3(new_n819), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT51), .B1(new_n736), .B2(new_n818), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(G106gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n827), .A2(G106gat), .A3(new_n368), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n844), .A2(KEYINPUT53), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n844), .A2(KEYINPUT53), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n849), .A2(new_n858), .ZN(G1339gat));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n681), .A2(new_n689), .A3(new_n694), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n692), .A2(KEYINPUT54), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n694), .B1(new_n681), .B2(new_n689), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n699), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(KEYINPUT55), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n702), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT55), .B1(new_n862), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n868), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(KEYINPUT111), .A3(new_n702), .A4(new_n866), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n869), .B(new_n871), .C1(new_n746), .C2(new_n747), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n592), .A2(new_n593), .A3(new_n589), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n583), .B1(new_n595), .B2(new_n582), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n601), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n703), .A2(new_n605), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n741), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n605), .A2(new_n875), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n741), .A2(new_n878), .A3(new_n869), .A4(new_n871), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n634), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n704), .A2(new_n748), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n368), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n411), .A2(new_n512), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n800), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n604), .A2(new_n605), .ZN(new_n888));
  OAI21_X1  g687(.A(G113gat), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT112), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n484), .B1(new_n881), .B2(new_n882), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n521), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n411), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(G113gat), .A3(new_n748), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n890), .A2(new_n895), .ZN(G1340gat));
  INV_X1    g695(.A(new_n894), .ZN(new_n897));
  AOI21_X1  g696(.A(G120gat), .B1(new_n897), .B2(new_n703), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n703), .A2(G120gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n886), .B2(new_n899), .ZN(G1341gat));
  OAI21_X1  g699(.A(G127gat), .B1(new_n887), .B2(new_n634), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n634), .A2(G127gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n894), .B2(new_n902), .ZN(G1342gat));
  NAND2_X1  g702(.A1(new_n411), .A2(new_n680), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(G134gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n893), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n907));
  OAI21_X1  g706(.A(G134gat), .B1(new_n887), .B2(new_n726), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(KEYINPUT56), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(G1343gat));
  NOR2_X1   g709(.A1(new_n718), .A2(new_n884), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n881), .A2(new_n882), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n912), .B2(new_n368), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT57), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n476), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n870), .A2(new_n702), .A3(new_n866), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n876), .B1(new_n888), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT113), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n920), .B(new_n876), .C1(new_n888), .C2(new_n917), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n680), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n634), .B1(new_n922), .B2(new_n880), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n916), .B1(new_n923), .B2(new_n882), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n606), .B(new_n911), .C1(new_n913), .C2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n921), .ZN(new_n928));
  INV_X1    g727(.A(new_n867), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n606), .A3(new_n870), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n920), .B1(new_n930), .B2(new_n876), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n726), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n633), .B1(new_n932), .B2(new_n879), .ZN(new_n933));
  INV_X1    g732(.A(new_n882), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n915), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n476), .B1(new_n881), .B2(new_n882), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(KEYINPUT57), .B2(new_n936), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n937), .A2(KEYINPUT116), .A3(new_n606), .A4(new_n911), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n938), .A3(G141gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT117), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n892), .A2(KEYINPUT115), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n719), .A2(new_n368), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n891), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n888), .A2(G141gat), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n941), .A2(new_n944), .A3(new_n411), .A4(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT58), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n939), .A2(new_n940), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n940), .B1(new_n939), .B2(new_n948), .ZN(new_n950));
  INV_X1    g749(.A(new_n946), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n911), .B1(new_n913), .B2(new_n924), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT114), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n937), .A2(KEYINPUT114), .A3(new_n911), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n749), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n951), .B1(new_n956), .B2(G141gat), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n949), .A2(new_n950), .B1(new_n947), .B2(new_n957), .ZN(G1344gat));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n944), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(new_n482), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n325), .A3(new_n703), .ZN(new_n961));
  XNOR2_X1  g760(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n680), .A2(new_n870), .A3(new_n929), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT119), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n680), .A2(new_n929), .A3(KEYINPUT119), .A4(new_n870), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n878), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n633), .B1(new_n932), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n704), .A2(new_n888), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n963), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n966), .A2(new_n878), .A3(new_n967), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n922), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g773(.A(KEYINPUT120), .B(new_n970), .C1(new_n974), .C2(new_n633), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n975), .A3(new_n368), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n914), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n916), .B1(new_n881), .B2(new_n882), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n703), .A3(new_n911), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n962), .B1(new_n981), .B2(G148gat), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n325), .A2(KEYINPUT59), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n954), .A2(new_n955), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n984), .B2(new_n703), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n961), .B1(new_n982), .B2(new_n985), .ZN(G1345gat));
  NAND2_X1  g785(.A1(new_n954), .A2(new_n955), .ZN(new_n987));
  OAI21_X1  g786(.A(G155gat), .B1(new_n987), .B2(new_n634), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n960), .A2(new_n626), .A3(new_n633), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1346gat));
  OAI21_X1  g789(.A(G162gat), .B1(new_n987), .B2(new_n742), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n904), .A2(G162gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n959), .B2(new_n992), .ZN(G1347gat));
  NOR2_X1   g792(.A1(new_n411), .A2(new_n512), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n995), .A2(new_n800), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n883), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n998), .A2(new_n218), .A3(new_n749), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT121), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n996), .B(KEYINPUT122), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(new_n883), .ZN(new_n1002));
  OAI21_X1  g801(.A(G169gat), .B1(new_n1002), .B2(new_n888), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1000), .A2(new_n1003), .ZN(G1348gat));
  OAI21_X1  g803(.A(G176gat), .B1(new_n1002), .B2(new_n750), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n998), .A2(new_n219), .A3(new_n703), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1349gat));
  OAI21_X1  g806(.A(G183gat), .B1(new_n1002), .B2(new_n634), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n998), .A2(new_n210), .A3(new_n633), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g810(.A1(new_n998), .A2(new_n211), .A3(new_n741), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1001), .A2(new_n680), .A3(new_n883), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1013), .A2(new_n1014), .A3(G190gat), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1014), .B1(new_n1013), .B2(G190gat), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g816(.A(new_n1017), .B(KEYINPUT123), .Z(G1351gat));
  NOR2_X1   g817(.A1(new_n995), .A2(new_n718), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n936), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(G197gat), .B1(new_n1020), .B2(new_n749), .ZN(new_n1021));
  INV_X1    g820(.A(new_n980), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1019), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g823(.A1(new_n606), .A2(G197gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(G1352gat));
  OAI21_X1  g825(.A(new_n970), .B1(new_n974), .B2(new_n633), .ZN(new_n1027));
  AOI21_X1  g826(.A(new_n476), .B1(new_n1027), .B2(new_n963), .ZN(new_n1028));
  AOI21_X1  g827(.A(KEYINPUT57), .B1(new_n1028), .B2(new_n975), .ZN(new_n1029));
  OAI211_X1 g828(.A(new_n703), .B(new_n1019), .C1(new_n1029), .C2(new_n978), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1030), .A2(KEYINPUT126), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT126), .ZN(new_n1032));
  NAND4_X1  g831(.A1(new_n980), .A2(new_n1032), .A3(new_n703), .A4(new_n1019), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1031), .A2(G204gat), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g833(.A1(new_n750), .A2(G204gat), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g835(.A(KEYINPUT124), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g837(.A1(new_n1020), .A2(KEYINPUT124), .A3(new_n1035), .ZN(new_n1039));
  INV_X1    g838(.A(KEYINPUT125), .ZN(new_n1040));
  AOI22_X1  g839(.A1(new_n1038), .A2(new_n1039), .B1(new_n1040), .B2(KEYINPUT62), .ZN(new_n1041));
  AND2_X1   g840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1042));
  XOR2_X1   g841(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1043));
  AOI21_X1  g842(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g843(.A1(new_n1034), .A2(new_n1044), .ZN(G1353gat));
  INV_X1    g844(.A(G211gat), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n1020), .A2(new_n1046), .A3(new_n633), .ZN(new_n1047));
  OAI211_X1 g846(.A(new_n633), .B(new_n1019), .C1(new_n1029), .C2(new_n978), .ZN(new_n1048));
  AND3_X1   g847(.A1(new_n1048), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1049));
  AOI21_X1  g848(.A(KEYINPUT63), .B1(new_n1048), .B2(G211gat), .ZN(new_n1050));
  OAI21_X1  g849(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(G1354gat));
  INV_X1    g850(.A(G218gat), .ZN(new_n1052));
  NAND3_X1  g851(.A1(new_n1020), .A2(new_n1052), .A3(new_n741), .ZN(new_n1053));
  NOR3_X1   g852(.A1(new_n1022), .A2(new_n726), .A3(new_n1023), .ZN(new_n1054));
  OAI21_X1  g853(.A(new_n1053), .B1(new_n1054), .B2(new_n1052), .ZN(G1355gat));
endmodule


