//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  XOR2_X1   g000(.A(KEYINPUT70), .B(G217), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(G146), .ZN(new_n196));
  INV_X1    g010(.A(G110), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT23), .B1(new_n200), .B2(G119), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n197), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT24), .B(G110), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(G119), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT71), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n198), .A2(new_n207), .A3(G119), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n205), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n196), .A2(new_n204), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT73), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n205), .A3(new_n210), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n199), .A2(new_n203), .A3(new_n197), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT72), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(KEYINPUT72), .A3(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n192), .A2(G146), .A3(new_n194), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT64), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n191), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n214), .B1(new_n221), .B2(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n215), .A2(KEYINPUT72), .A3(new_n216), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT72), .B1(new_n215), .B2(new_n216), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n230), .B(new_n214), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n213), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT22), .B(G137), .Z(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(G221), .A3(G234), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n237), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT73), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n212), .B1(new_n245), .B2(new_n234), .ZN(new_n246));
  INV_X1    g060(.A(new_n242), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n243), .A2(new_n188), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n243), .A2(new_n248), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n190), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n243), .A2(new_n248), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n189), .A2(G902), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(G472), .A2(G902), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT31), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n225), .A2(G143), .A3(new_n226), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n198), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n265), .A2(G146), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n227), .B2(new_n265), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT11), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(G137), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT11), .A3(G134), .ZN(new_n277));
  INV_X1    g091(.A(G131), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(G137), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n275), .A2(new_n277), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n274), .A2(G137), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n276), .A2(G134), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n283), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n272), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n275), .A2(new_n277), .A3(new_n279), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G131), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n280), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n264), .A2(KEYINPUT0), .A3(G128), .A4(new_n266), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT0), .B(G128), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n291), .B(new_n292), .C1(new_n271), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT30), .B1(new_n288), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n271), .A2(new_n293), .ZN(new_n296));
  INV_X1    g110(.A(new_n292), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n286), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n298), .A2(new_n291), .B1(new_n299), .B2(new_n272), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n295), .A2(KEYINPUT67), .B1(new_n300), .B2(KEYINPUT30), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n288), .A2(new_n294), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT30), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G116), .B(G119), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT2), .B(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n309), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n307), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n301), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n300), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(new_n313), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n317));
  NOR2_X1   g131(.A1(G237), .A2(G953), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G210), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G101), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n320), .B(new_n321), .Z(new_n322));
  NOR2_X1   g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n263), .B1(new_n314), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n300), .A2(new_n310), .A3(new_n312), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT28), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n302), .A2(new_n313), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n314), .A2(new_n323), .A3(new_n263), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT69), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n314), .A2(new_n323), .A3(new_n332), .A4(new_n263), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n262), .B1(new_n329), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n337));
  AOI211_X1 g151(.A(KEYINPUT32), .B(new_n262), .C1(new_n329), .C2(new_n334), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n315), .A2(new_n313), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n326), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(KEYINPUT29), .ZN(new_n343));
  INV_X1    g157(.A(new_n322), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n328), .B2(KEYINPUT29), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n188), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n316), .A2(new_n344), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n314), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(KEYINPUT29), .ZN(new_n349));
  OAI21_X1  g163(.A(G472), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n260), .B1(new_n340), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G214), .B1(G237), .B2(G902), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G104), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G107), .ZN(new_n355));
  INV_X1    g169(.A(G107), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G101), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n355), .B2(new_n357), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(new_n354), .B2(G107), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n356), .A3(G104), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G101), .B1(new_n354), .B2(G107), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n361), .A2(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n307), .A2(KEYINPUT5), .ZN(new_n371));
  INV_X1    g185(.A(G116), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n372), .A2(KEYINPUT5), .A3(G119), .ZN(new_n373));
  INV_X1    g187(.A(G113), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n371), .A2(new_n375), .B1(new_n311), .B2(new_n307), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n370), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT8), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n380), .B(KEYINPUT90), .Z(new_n381));
  NAND2_X1  g195(.A1(new_n238), .A2(G224), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT7), .ZN(new_n383));
  OAI21_X1  g197(.A(G125), .B1(new_n296), .B2(new_n297), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT87), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n269), .A2(new_n271), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n193), .A3(new_n268), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n383), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n389), .A2(KEYINPUT91), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(KEYINPUT91), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n381), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n365), .A2(new_n367), .A3(new_n355), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT77), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n396), .A2(new_n398), .B1(new_n310), .B2(new_n312), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(G101), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n365), .A2(new_n369), .A3(new_n367), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT76), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT76), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n400), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n399), .B(KEYINPUT83), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n370), .A2(new_n376), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n402), .A2(KEYINPUT76), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(new_n404), .A3(new_n400), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT83), .B1(new_n412), .B2(new_n399), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n378), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n385), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n384), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT88), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n420), .A3(new_n387), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n415), .B1(new_n421), .B2(new_n383), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n188), .B1(new_n392), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n409), .B2(new_n413), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n399), .B1(new_n403), .B2(new_n406), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n429), .A2(KEYINPUT84), .A3(new_n408), .A4(new_n407), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n378), .B(KEYINPUT85), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n426), .A2(KEYINPUT86), .A3(new_n430), .A4(new_n433), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n426), .A2(new_n430), .A3(new_n431), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n432), .B1(new_n414), .B2(new_n378), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n421), .A2(G224), .A3(new_n238), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n417), .A2(new_n420), .A3(new_n382), .A4(new_n387), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND4_X1   g258(.A1(KEYINPUT89), .A2(new_n438), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n436), .A2(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT89), .B1(new_n446), .B2(new_n444), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n424), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n438), .A2(new_n441), .A3(new_n444), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(KEYINPUT89), .A3(new_n444), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n449), .A3(new_n424), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n353), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT9), .B(G234), .ZN(new_n459));
  OAI21_X1  g273(.A(G221), .B1(new_n459), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n396), .A2(new_n398), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n412), .A2(new_n298), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n370), .A2(KEYINPUT10), .A3(new_n272), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n264), .A2(new_n266), .ZN(new_n465));
  INV_X1    g279(.A(new_n270), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n200), .B1(new_n466), .B2(KEYINPUT1), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n268), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n370), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n291), .B(KEYINPUT80), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n463), .A2(new_n464), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G140), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n238), .A2(G227), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n364), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n401), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n386), .A3(new_n268), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n469), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT12), .B1(new_n483), .B2(new_n291), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n485));
  INV_X1    g299(.A(new_n291), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n485), .B(new_n486), .C1(new_n482), .C2(new_n469), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT81), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n370), .A2(new_n468), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n370), .A2(new_n272), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n291), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n485), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT81), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n483), .A2(KEYINPUT12), .A3(new_n291), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n478), .A2(new_n488), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n478), .A2(new_n488), .A3(new_n495), .A4(KEYINPUT82), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n463), .A2(new_n464), .A3(new_n471), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n291), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n473), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n476), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G469), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n188), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n473), .B1(new_n484), .B2(new_n487), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n478), .A2(new_n501), .B1(new_n507), .B2(new_n476), .ZN(new_n508));
  OAI21_X1  g322(.A(G469), .B1(new_n508), .B2(G902), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n461), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(G234), .A2(G237), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n512), .A2(G952), .A3(new_n238), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n512), .A2(G902), .A3(G953), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n198), .A2(G143), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n265), .A2(G128), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT13), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n265), .A2(KEYINPUT13), .A3(G128), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G134), .ZN(new_n523));
  XNOR2_X1  g337(.A(G116), .B(G122), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G107), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n356), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n518), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n523), .B(new_n528), .C1(G134), .C2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n274), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n527), .A2(KEYINPUT95), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n372), .A2(KEYINPUT14), .A3(G122), .ZN(new_n533));
  OAI211_X1 g347(.A(G107), .B(new_n533), .C1(new_n525), .C2(KEYINPUT14), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(KEYINPUT95), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n530), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n187), .A2(G953), .A3(new_n459), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n530), .B(new_n538), .C1(new_n531), .C2(new_n536), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(KEYINPUT96), .A3(new_n539), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n188), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT97), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(KEYINPUT97), .A3(new_n188), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G478), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(KEYINPUT15), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(new_n552), .A3(G478), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n229), .B1(new_n224), .B2(new_n191), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n318), .A2(G143), .A3(G214), .ZN(new_n558));
  AOI21_X1  g372(.A(G143), .B1(new_n318), .B2(G214), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(new_n278), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT18), .B(G131), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT92), .Z(new_n565));
  OAI211_X1 g379(.A(KEYINPUT17), .B(G131), .C1(new_n558), .C2(new_n559), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n560), .B(new_n278), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n196), .B(new_n566), .C1(new_n567), .C2(KEYINPUT17), .ZN(new_n568));
  XNOR2_X1  g382(.A(G113), .B(G122), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n354), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n191), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT19), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n575), .A2(KEYINPUT94), .A3(new_n228), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT94), .B1(new_n575), .B2(new_n228), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n222), .B(new_n567), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n570), .B1(new_n565), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n556), .B1(new_n571), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT20), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(KEYINPUT20), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n570), .B1(new_n565), .B2(new_n568), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n188), .B1(new_n571), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n582), .A2(new_n583), .B1(G475), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n555), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n511), .A2(new_n516), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n351), .A2(new_n458), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  AOI21_X1  g404(.A(G902), .B1(new_n329), .B2(new_n334), .ZN(new_n591));
  INV_X1    g405(.A(G472), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n336), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n594), .A2(new_n511), .A3(new_n260), .ZN(new_n595));
  INV_X1    g409(.A(new_n516), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n545), .A2(new_n550), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT100), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n542), .A2(KEYINPUT33), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n537), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n530), .B(KEYINPUT98), .C1(new_n531), .C2(new_n536), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n539), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT99), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n601), .A2(new_n605), .A3(new_n539), .A4(new_n602), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n599), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n543), .A2(new_n544), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(KEYINPUT33), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n550), .A2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n598), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n585), .A2(G475), .ZN(new_n614));
  INV_X1    g428(.A(new_n583), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(new_n581), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n595), .A2(new_n458), .A3(new_n596), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NAND2_X1  g435(.A1(new_n586), .A2(new_n554), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n458), .A2(new_n596), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n595), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT101), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT35), .B(G107), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n242), .A2(KEYINPUT36), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n246), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n246), .A2(new_n630), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n256), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n253), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT102), .B1(new_n594), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n591), .A2(new_n592), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n335), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT102), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n251), .A2(new_n252), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n189), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n634), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n639), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n637), .A2(new_n458), .A3(new_n588), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  INV_X1    g461(.A(KEYINPUT32), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n335), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n350), .B1(new_n649), .B2(new_n338), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n650), .A2(new_n510), .A3(new_n643), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n514), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n513), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n586), .A2(new_n554), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n651), .A2(new_n458), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT103), .B(G128), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G30));
  NAND2_X1  g474(.A1(new_n451), .A2(new_n457), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT38), .Z(new_n662));
  AOI21_X1  g476(.A(new_n322), .B1(new_n314), .B2(new_n325), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(G902), .B1(new_n347), .B2(new_n341), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n592), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n337), .B2(new_n339), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n655), .B(KEYINPUT39), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n510), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n667), .B1(KEYINPUT40), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n616), .A2(new_n554), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n643), .A2(new_n671), .A3(new_n353), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n670), .B(new_n672), .C1(KEYINPUT40), .C2(new_n669), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n662), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  INV_X1    g489(.A(new_n655), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n617), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n449), .B1(new_n456), .B2(new_n424), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n450), .B(new_n423), .C1(new_n454), .C2(new_n455), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n352), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n661), .A2(KEYINPUT104), .A3(new_n352), .A4(new_n677), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n651), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  AND3_X1   g499(.A1(new_n504), .A2(new_n505), .A3(new_n188), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n505), .B1(new_n504), .B2(new_n188), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n687), .A3(new_n461), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n650), .A2(new_n259), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n458), .A3(new_n596), .A4(new_n618), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT41), .B(G113), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G15));
  NAND4_X1  g506(.A1(new_n689), .A2(new_n458), .A3(new_n596), .A4(new_n623), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  NOR2_X1   g508(.A1(new_n616), .A2(new_n554), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n650), .A2(new_n596), .A3(new_n695), .A4(new_n643), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n458), .A3(new_n688), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  AOI21_X1  g512(.A(new_n324), .B1(new_n322), .B2(new_n342), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n262), .B1(new_n699), .B2(new_n334), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n700), .A2(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(KEYINPUT105), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n701), .A2(new_n593), .A3(new_n259), .A4(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n688), .A2(new_n596), .ZN(new_n705));
  INV_X1    g519(.A(new_n671), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n458), .A2(new_n704), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  OAI22_X1  g522(.A1(KEYINPUT105), .A2(new_n700), .B1(new_n591), .B2(new_n592), .ZN(new_n709));
  INV_X1    g523(.A(new_n702), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n709), .A2(new_n710), .A3(new_n636), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n458), .A2(new_n677), .A3(new_n688), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  NAND4_X1  g527(.A1(new_n451), .A2(new_n352), .A3(new_n457), .A4(new_n510), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n650), .A2(new_n259), .ZN(new_n715));
  INV_X1    g529(.A(new_n677), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  NOR2_X1   g536(.A1(new_n714), .A2(new_n715), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n656), .B(KEYINPUT107), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(KEYINPUT108), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  INV_X1    g544(.A(new_n613), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n616), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT43), .B1(new_n731), .B2(new_n616), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n643), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n737));
  OR3_X1    g551(.A1(new_n736), .A2(new_n737), .A3(new_n639), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n508), .A2(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n508), .A2(KEYINPUT45), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(G469), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(G469), .A2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n506), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n744), .B1(KEYINPUT46), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT109), .B1(new_n743), .B2(new_n506), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n460), .B(new_n668), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n451), .A2(new_n352), .A3(new_n457), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n737), .B1(new_n736), .B2(new_n639), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n738), .A2(new_n749), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT110), .B(G137), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G39));
  OAI21_X1  g569(.A(new_n460), .B1(new_n746), .B2(new_n747), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n750), .A2(new_n716), .A3(new_n650), .A4(new_n259), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  NAND2_X1  g579(.A1(new_n734), .A2(new_n735), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(new_n703), .A3(new_n654), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n458), .A3(new_n688), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(G952), .A3(new_n238), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n751), .A2(new_n688), .ZN(new_n770));
  INV_X1    g584(.A(new_n667), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n770), .A2(new_n260), .A3(new_n654), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n769), .B1(new_n618), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT48), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n766), .A2(new_n654), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n751), .A3(new_n688), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT118), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n751), .A3(new_n778), .A4(new_n688), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n774), .B1(new_n780), .B2(new_n351), .ZN(new_n781));
  AOI211_X1 g595(.A(KEYINPUT48), .B(new_n715), .C1(new_n777), .C2(new_n779), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n773), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT120), .Z(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n780), .A2(new_n786), .A3(new_n711), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n780), .B2(new_n711), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n688), .A2(new_n353), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT117), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n662), .A2(new_n767), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n686), .A2(new_n687), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n758), .B(new_n759), .C1(new_n460), .C2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n767), .A2(new_n751), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n613), .A2(new_n616), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n798), .A2(new_n799), .B1(new_n772), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n785), .B1(new_n790), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n789), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n787), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(KEYINPUT51), .A3(new_n795), .A4(new_n801), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n784), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n619), .A2(new_n645), .A3(new_n589), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n352), .B(new_n596), .C1(new_n678), .C2(new_n679), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n622), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n458), .A2(KEYINPUT113), .A3(new_n596), .A4(new_n623), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n595), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n697), .A2(new_n707), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT112), .A3(new_n690), .A4(new_n693), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n690), .A2(new_n697), .A3(new_n693), .A4(new_n707), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n814), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n711), .A2(new_n677), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n587), .A2(new_n676), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n352), .A3(new_n451), .A4(new_n457), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n650), .A2(new_n510), .A3(new_n643), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n821), .A2(new_n714), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n729), .A2(new_n721), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n643), .B2(new_n676), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n636), .A2(KEYINPUT114), .A3(new_n655), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n511), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n458), .A3(new_n706), .A4(new_n771), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n684), .A2(new_n658), .A3(new_n712), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n658), .A2(new_n712), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT114), .B1(new_n636), .B2(new_n655), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n253), .A2(new_n635), .A3(new_n828), .A4(new_n676), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n510), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n667), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n353), .B(new_n671), .C1(new_n451), .C2(new_n457), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n834), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n836), .A2(new_n684), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n820), .A2(new_n827), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n832), .A2(new_n658), .A3(KEYINPUT52), .A4(new_n712), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n682), .A2(new_n651), .A3(new_n683), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT115), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n836), .A2(new_n850), .A3(new_n842), .A4(new_n684), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n835), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n820), .A2(new_n852), .A3(new_n853), .A4(new_n827), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n845), .A2(new_n853), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n835), .A2(new_n849), .A3(new_n851), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n645), .A2(new_n589), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n858), .A2(new_n619), .A3(new_n813), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n817), .A2(new_n853), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n723), .A2(new_n677), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n719), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n825), .B1(new_n862), .B2(new_n718), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n859), .A2(new_n860), .A3(new_n863), .A4(new_n729), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT116), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n690), .A2(new_n697), .A3(new_n693), .A4(new_n707), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(KEYINPUT53), .A3(new_n813), .A4(new_n808), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n729), .A2(new_n721), .A3(new_n826), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n870), .B2(new_n852), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n856), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n855), .B1(new_n872), .B2(KEYINPUT54), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n807), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n732), .A2(new_n259), .A3(new_n352), .A4(new_n460), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n662), .A2(new_n667), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n874), .A2(new_n879), .ZN(G75));
  NAND3_X1  g694(.A1(new_n872), .A2(G210), .A3(G902), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n446), .B(new_n444), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT55), .Z(new_n884));
  AND3_X1   g698(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n881), .B2(new_n882), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n238), .A2(G952), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(G51));
  XOR2_X1   g702(.A(new_n742), .B(KEYINPUT57), .Z(new_n889));
  OAI21_X1  g703(.A(KEYINPUT116), .B1(new_n857), .B2(new_n864), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n870), .A2(new_n866), .A3(new_n852), .ZN(new_n891));
  AOI221_X4 g705(.A(KEYINPUT54), .B1(new_n845), .B2(new_n853), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n856), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n889), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n504), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n890), .A2(new_n891), .B1(new_n853), .B2(new_n845), .ZN(new_n898));
  OR3_X1    g712(.A1(new_n898), .A2(new_n188), .A3(new_n741), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n887), .B1(new_n897), .B2(new_n899), .ZN(G54));
  AND2_X1   g714(.A1(KEYINPUT58), .A2(G475), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n872), .A2(G902), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n571), .A2(new_n579), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n902), .A2(KEYINPUT121), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT121), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  INV_X1    g719(.A(new_n903), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n872), .A2(G902), .A3(new_n906), .A4(new_n901), .ZN(new_n907));
  INV_X1    g721(.A(new_n887), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n904), .A2(new_n905), .A3(new_n909), .ZN(G60));
  NAND2_X1  g724(.A1(G478), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT59), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n610), .B1(new_n873), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n610), .A2(new_n912), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n898), .A2(new_n893), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n913), .A2(new_n887), .A3(new_n917), .ZN(G63));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT60), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n255), .B1(new_n898), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n920), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n872), .A2(new_n633), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n923), .A3(new_n908), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT61), .A4(new_n908), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G66));
  INV_X1    g742(.A(new_n515), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n238), .B1(new_n929), .B2(G224), .ZN(new_n930));
  INV_X1    g744(.A(new_n820), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(new_n238), .ZN(new_n932));
  INV_X1    g746(.A(new_n446), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(G898), .B2(new_n238), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT122), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n932), .B(new_n935), .ZN(G69));
  AND2_X1   g750(.A1(new_n836), .A2(new_n684), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n674), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n938), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT124), .B1(new_n938), .B2(KEYINPUT62), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n669), .B1(new_n617), .B2(new_n622), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n751), .A2(new_n351), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n764), .A2(new_n753), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(G953), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n301), .A2(new_n306), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n575), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT123), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n937), .A2(new_n753), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n749), .A2(new_n351), .A3(new_n841), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n721), .A2(new_n764), .A3(new_n729), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(G953), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n949), .B1(G900), .B2(G953), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI22_X1  g773(.A1(new_n947), .A2(new_n950), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n238), .B1(G227), .B2(G900), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n960), .B(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n956), .B2(new_n931), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n314), .A3(new_n347), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n846), .A2(new_n854), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n664), .A2(new_n348), .A3(new_n967), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n969), .B(new_n908), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n946), .B(new_n820), .C1(new_n939), .C2(new_n940), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n973), .A2(KEYINPUT127), .A3(new_n967), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT127), .B1(new_n973), .B2(new_n967), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n974), .A2(new_n975), .A3(new_n664), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n972), .A2(new_n976), .ZN(G57));
endmodule


