//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g0014(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT65), .B(G238), .Z(new_n227));
  OAI211_X1 g0027(.A(new_n224), .B(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(new_n230));
  OAI21_X1  g0030(.A(new_n208), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n211), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT67), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G150), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n206), .A2(G33), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n252), .B1(new_n201), .B2(new_n206), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n214), .A2(new_n215), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n214), .A2(new_n259), .A3(new_n215), .A4(new_n256), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n205), .A2(G20), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT69), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(new_n265), .A3(G50), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT9), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(G226), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n287), .A2(G223), .B1(new_n290), .B2(G77), .ZN(new_n291));
  AOI21_X1  g0091(.A(G1698), .B1(new_n285), .B2(new_n286), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G222), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n216), .A2(new_n275), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n281), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n261), .A2(KEYINPUT9), .A3(new_n266), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n297), .B(new_n298), .C1(new_n299), .C2(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT10), .B1(new_n271), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n269), .B(KEYINPUT71), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n267), .C1(G179), .C2(new_n296), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g0110(.A(new_n264), .B(KEYINPUT69), .Z(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(new_n253), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(new_n263), .B1(new_n260), .B2(new_n253), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n285), .A2(new_n206), .A3(new_n286), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n286), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(KEYINPUT77), .A3(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(KEYINPUT77), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(G68), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G58), .A2(G68), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT76), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n324), .B(new_n325), .C1(G58), .C2(G68), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n214), .A2(new_n215), .A3(new_n256), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n326), .A2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n251), .A2(G159), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n226), .B1(new_n317), .B2(new_n318), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n336), .B2(KEYINPUT16), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n314), .B1(new_n330), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G226), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G1698), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G223), .B2(G1698), .ZN(new_n341));
  INV_X1    g0141(.A(G87), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n341), .A2(new_n290), .B1(new_n284), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n216), .A2(new_n275), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT78), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT78), .B1(new_n343), .B2(new_n344), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT79), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n276), .A2(new_n279), .A3(new_n348), .A4(G232), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n349), .A2(new_n277), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n276), .A2(G232), .A3(new_n279), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT79), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G223), .A2(G1698), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n339), .B2(G1698), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT3), .B(G33), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n357), .A2(new_n358), .B1(G33), .B2(G87), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n350), .B(new_n352), .C1(new_n295), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n307), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT18), .B1(new_n338), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n353), .A2(G190), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G200), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n338), .A2(KEYINPUT17), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT17), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT16), .B1(new_n321), .B2(new_n327), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT7), .B1(new_n290), .B2(new_n206), .ZN(new_n372));
  INV_X1    g0172(.A(new_n318), .ZN(new_n373));
  OAI21_X1  g0173(.A(G68), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n257), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n313), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n347), .A2(new_n364), .B1(new_n360), .B2(new_n366), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n370), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n347), .A2(new_n354), .B1(new_n360), .B2(new_n307), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n377), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n363), .A2(new_n369), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n311), .A2(new_n202), .A3(new_n262), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n202), .B2(new_n260), .ZN(new_n385));
  INV_X1    g0185(.A(new_n251), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n253), .A2(new_n386), .B1(new_n206), .B2(new_n202), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT70), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT15), .B(G87), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n387), .A2(new_n388), .B1(new_n254), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n387), .A2(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n257), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n292), .A2(G232), .B1(new_n290), .B2(G107), .ZN(new_n394));
  INV_X1    g0194(.A(new_n287), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n227), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n344), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n278), .B1(G244), .B2(new_n280), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n393), .B1(new_n400), .B2(G190), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n366), .B2(new_n400), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n392), .A2(new_n385), .B1(new_n399), .B2(new_n307), .ZN(new_n403));
  INV_X1    g0203(.A(G179), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n310), .A2(new_n383), .A3(new_n407), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n254), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n409), .A2(KEYINPUT75), .B1(new_n258), .B2(new_n386), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(KEYINPUT75), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n257), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT11), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n311), .A2(new_n226), .A3(new_n262), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT12), .B1(new_n259), .B2(G68), .ZN(new_n416));
  OR3_X1    g0216(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n413), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n414), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n278), .B1(G238), .B2(new_n280), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT73), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(G33), .A3(G97), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n292), .B2(G226), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT72), .B1(new_n287), .B2(G232), .ZN(new_n429));
  OAI211_X1 g0229(.A(G232), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT72), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n422), .B(new_n428), .C1(new_n429), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n344), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n430), .B(new_n431), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n422), .B1(new_n435), .B2(new_n428), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n421), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(new_n421), .C1(new_n434), .C2(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n420), .B1(new_n441), .B2(new_n299), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n366), .B1(new_n438), .B2(new_n440), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n440), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n428), .B1(new_n429), .B2(new_n432), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT74), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n344), .A3(new_n433), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n439), .B1(new_n448), .B2(new_n421), .ZN(new_n449));
  OAI21_X1  g0249(.A(G169), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n438), .A2(G179), .A3(new_n440), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT14), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(G169), .C1(new_n445), .C2(new_n449), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n420), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n444), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n408), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(G244), .B(new_n282), .C1(new_n288), .C2(new_n289), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n461), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n358), .A2(G244), .A3(new_n282), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n358), .A2(G250), .A3(G1698), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G283), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n462), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n344), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n273), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G257), .A3(new_n276), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n469), .A2(new_n276), .A3(G274), .A4(new_n470), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n468), .A2(G179), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n344), .B2(new_n467), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n307), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n319), .A2(G107), .A3(new_n320), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G97), .A2(G107), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(KEYINPUT6), .A3(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n257), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n259), .A2(G97), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n284), .A2(G1), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n262), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(G97), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT81), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n331), .B1(new_n479), .B2(new_n488), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT81), .ZN(new_n497));
  INV_X1    g0297(.A(new_n494), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n478), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n468), .A2(new_n474), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n299), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n477), .A2(new_n366), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n496), .A2(new_n498), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n358), .A2(KEYINPUT82), .A3(G244), .A4(G1698), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(G238), .B(new_n282), .C1(new_n288), .C2(new_n289), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n295), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n470), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n517), .A2(G250), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n276), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n276), .A2(G274), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n517), .ZN(new_n521));
  OAI21_X1  g0321(.A(G200), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n484), .A2(new_n342), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT19), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n424), .B2(new_n426), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n525), .B2(G20), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n206), .B(G68), .C1(new_n288), .C2(new_n289), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n254), .B2(new_n481), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n331), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n389), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n259), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n262), .A2(new_n342), .A3(new_n492), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n520), .A2(new_n517), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n276), .B2(new_n518), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n514), .B1(new_n509), .B2(new_n510), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(G190), .C1(new_n537), .C2(new_n295), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n522), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n307), .B1(new_n516), .B2(new_n521), .ZN(new_n540));
  INV_X1    g0340(.A(new_n532), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n493), .A2(new_n531), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n527), .A2(new_n528), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n425), .B1(G33), .B2(G97), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n423), .A2(KEYINPUT73), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT19), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n206), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n523), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n541), .B(new_n542), .C1(new_n548), .C2(new_n331), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n536), .B(new_n404), .C1(new_n537), .C2(new_n295), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n540), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n539), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n500), .A2(new_n506), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n500), .A2(new_n506), .A3(new_n552), .A4(KEYINPUT83), .ZN(new_n556));
  INV_X1    g0356(.A(new_n473), .ZN(new_n557));
  INV_X1    g0357(.A(new_n212), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n469), .A2(new_n470), .B1(new_n558), .B2(new_n275), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(G270), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G264), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n561));
  OAI211_X1 g0361(.A(G257), .B(new_n282), .C1(new_n288), .C2(new_n289), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n285), .A2(G303), .A3(new_n286), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT84), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n562), .A3(new_n567), .A4(new_n563), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n344), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n560), .B(G190), .C1(new_n566), .C2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n492), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n331), .A2(G116), .A3(new_n259), .A4(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n260), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(G33), .B2(G283), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n284), .A2(G97), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(G20), .B2(new_n573), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n577), .A2(new_n257), .A3(KEYINPUT20), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT20), .B1(new_n577), .B2(new_n257), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n572), .B(new_n574), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n559), .A2(G270), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n473), .ZN(new_n583));
  INV_X1    g0383(.A(new_n569), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n565), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n570), .B(new_n581), .C1(new_n585), .C2(new_n366), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n580), .A2(G169), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(G179), .A3(new_n580), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n560), .B1(new_n566), .B2(new_n569), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(KEYINPUT21), .A3(G169), .A4(new_n580), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n586), .A2(new_n589), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n594));
  OAI211_X1 g0394(.A(G250), .B(new_n282), .C1(new_n288), .C2(new_n289), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G294), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n344), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n559), .A2(G264), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n473), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(new_n299), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n597), .A2(new_n344), .B1(new_n559), .B2(G264), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n366), .B1(new_n602), .B2(new_n473), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT85), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n206), .B(G87), .C1(new_n288), .C2(new_n289), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT22), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT22), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n358), .A2(new_n609), .A3(new_n206), .A4(G87), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n482), .A2(KEYINPUT23), .A3(G20), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT23), .B1(new_n482), .B2(G20), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(G20), .B2(new_n513), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n605), .B(new_n606), .C1(new_n611), .C2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n608), .B2(new_n610), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT24), .B1(new_n616), .B2(KEYINPUT85), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n605), .B(new_n614), .C1(new_n608), .C2(new_n610), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n615), .B(new_n257), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT86), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT25), .ZN(new_n621));
  INV_X1    g0421(.A(G13), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G1), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n206), .A2(G107), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n620), .A2(KEYINPUT25), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n623), .A2(new_n626), .A3(new_n624), .A4(new_n621), .ZN(new_n627));
  AOI211_X1 g0427(.A(new_n625), .B(new_n627), .C1(G107), .C2(new_n493), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n604), .A2(new_n619), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n600), .A2(new_n307), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n602), .A2(new_n404), .A3(new_n473), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n619), .B2(new_n628), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n593), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n459), .A2(new_n555), .A3(new_n556), .A4(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n454), .A2(new_n452), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n453), .B1(new_n441), .B2(G169), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n456), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n444), .B2(new_n406), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n369), .A2(new_n379), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n363), .A2(new_n382), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n306), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n309), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n619), .A2(new_n628), .ZN(new_n648));
  INV_X1    g0448(.A(new_n633), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n592), .A2(new_n590), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n589), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n490), .A2(KEYINPUT81), .A3(new_n494), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n497), .B1(new_n496), .B2(new_n498), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n655), .A2(new_n478), .B1(new_n504), .B2(new_n505), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n652), .A2(new_n656), .A3(new_n552), .A4(new_n629), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n490), .A2(new_n494), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n551), .A2(new_n539), .A3(new_n659), .A4(new_n478), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n501), .A2(G169), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n653), .A2(new_n654), .B1(new_n663), .B2(new_n475), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(new_n552), .A3(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n664), .A2(new_n552), .A3(new_n658), .A4(KEYINPUT26), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n657), .A2(new_n666), .A3(new_n551), .A4(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n647), .B1(new_n458), .B2(new_n669), .ZN(G369));
  NAND2_X1  g0470(.A1(new_n623), .A2(new_n206), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT27), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT88), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n623), .A2(new_n674), .A3(new_n206), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G213), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n673), .B1(new_n672), .B2(new_n675), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G343), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT89), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n648), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT90), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(KEYINPUT90), .A3(new_n648), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n650), .A3(new_n629), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n634), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n681), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n589), .A2(new_n592), .A3(new_n590), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n688), .A2(new_n692), .B1(new_n634), .B2(new_n689), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n689), .A2(new_n581), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n690), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n593), .B2(new_n694), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n688), .A2(new_n696), .A3(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(G399));
  INV_X1    g0498(.A(new_n209), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(G41), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n523), .A2(G116), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT92), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n219), .B2(new_n701), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n666), .A2(new_n667), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n629), .B1(new_n690), .B2(new_n634), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n551), .B1(new_n553), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n689), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT94), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT94), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT26), .B1(new_n664), .B2(new_n552), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n660), .A2(new_n661), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n551), .B1(new_n553), .B2(new_n708), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT95), .B1(new_n719), .B2(new_n689), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n717), .A2(new_n718), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT95), .B(new_n689), .C1(new_n709), .C2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT29), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n555), .A2(new_n635), .A3(new_n556), .A4(new_n689), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n516), .A2(new_n521), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n477), .A3(new_n602), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n585), .A2(G179), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n477), .A2(new_n602), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n591), .A2(new_n404), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT30), .A4(new_n728), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n728), .A2(new_n477), .ZN(new_n735));
  AOI21_X1  g0535(.A(G179), .B1(new_n602), .B2(new_n473), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n591), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n731), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT93), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n735), .A2(KEYINPUT93), .A3(new_n591), .A4(new_n736), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(new_n734), .A3(new_n731), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n681), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n726), .A2(new_n739), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n725), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n706), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(new_n622), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n205), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OR3_X1    g0554(.A1(new_n700), .A2(KEYINPUT96), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT96), .B1(new_n700), .B2(new_n754), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n696), .B2(G330), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G330), .B2(new_n696), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n209), .A2(new_n358), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n209), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n699), .A2(new_n358), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n273), .B2(new_n220), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n249), .A2(G45), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n217), .B1(G20), .B2(new_n307), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n758), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n773), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n696), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n206), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n299), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n482), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n206), .A2(new_n404), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n783), .A2(new_n299), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n785), .A2(new_n226), .B1(new_n787), .B2(new_n258), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n299), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n206), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n781), .B(new_n788), .C1(G97), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n779), .A2(G190), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT98), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G87), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G190), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n779), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G159), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT32), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n782), .A2(G190), .A3(new_n366), .ZN(new_n805));
  INV_X1    g0605(.A(G58), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n358), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n782), .A2(new_n800), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(G77), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n792), .A2(new_n799), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n797), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G326), .ZN(new_n814));
  INV_X1    g0614(.A(G294), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n787), .A2(new_n814), .B1(new_n815), .B2(new_n790), .ZN(new_n816));
  INV_X1    g0616(.A(new_n780), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(G283), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT33), .B(G317), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n820), .A2(new_n784), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G322), .ZN(new_n823));
  INV_X1    g0623(.A(G329), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n805), .A2(new_n823), .B1(new_n801), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n358), .B(new_n825), .C1(G311), .C2(new_n809), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n818), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n811), .B1(new_n813), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n776), .B(new_n778), .C1(new_n770), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n761), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n681), .A2(new_n393), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n402), .A2(new_n832), .B1(new_n405), .B2(new_n403), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n406), .A2(new_n681), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n710), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n668), .A2(new_n689), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n758), .B1(new_n839), .B2(new_n748), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n748), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n770), .A2(new_n771), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n805), .ZN(new_n844));
  INV_X1    g0644(.A(new_n801), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n844), .A2(G294), .B1(new_n845), .B2(G311), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n290), .C1(new_n573), .C2(new_n808), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n784), .A2(G283), .B1(new_n817), .B2(G87), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n848), .B1(new_n481), .B2(new_n790), .C1(new_n812), .C2(new_n787), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(G107), .C2(new_n798), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n358), .B1(new_n801), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G68), .B2(new_n817), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n806), .B2(new_n790), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n844), .A2(G143), .B1(new_n809), .B2(G159), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  INV_X1    g0656(.A(G150), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n855), .B1(new_n787), .B2(new_n856), .C1(new_n857), .C2(new_n785), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n854), .B(new_n860), .C1(G50), .C2(new_n798), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n850), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n770), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n758), .B1(G77), .B2(new_n843), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n771), .B2(new_n835), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT100), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n841), .A2(new_n867), .ZN(G384));
  NOR2_X1   g0668(.A1(new_n752), .A2(new_n205), .ZN(new_n869));
  INV_X1    g0669(.A(G330), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n456), .B(new_n681), .C1(new_n455), .C2(new_n444), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n442), .A2(new_n443), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n681), .A2(new_n456), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n639), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n835), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n375), .A3(new_n257), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n313), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(KEYINPUT102), .A3(new_n313), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n880), .A2(new_n679), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n383), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n338), .A2(new_n368), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n377), .A2(new_n380), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n377), .A2(new_n679), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n679), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n362), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n880), .A3(new_n881), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n885), .B1(new_n892), .B2(new_n884), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n883), .B(KEYINPUT38), .C1(new_n889), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  INV_X1    g0696(.A(new_n887), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n896), .A2(new_n888), .B1(new_n383), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(KEYINPUT38), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n726), .A2(new_n746), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n875), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n892), .A2(new_n884), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n888), .B1(new_n904), .B2(new_n885), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n883), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n894), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(new_n910), .A3(new_n875), .A4(new_n901), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT104), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n459), .A2(new_n901), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n870), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n913), .ZN(new_n916));
  AOI211_X1 g0716(.A(KEYINPUT94), .B(KEYINPUT29), .C1(new_n668), .C2(new_n689), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n714), .B1(new_n710), .B2(new_n711), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n459), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n689), .B1(new_n709), .B2(new_n721), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT95), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n711), .B1(new_n922), .B2(new_n722), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT103), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n716), .A2(new_n925), .A3(new_n459), .A4(new_n724), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n646), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n899), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n455), .A2(new_n456), .A3(new_n689), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n931), .C1(new_n909), .C2(new_n928), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n834), .B(KEYINPUT101), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n838), .A2(new_n934), .B1(new_n874), .B2(new_n871), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n909), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n644), .A2(new_n890), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n932), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n927), .B(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n869), .B1(new_n916), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n939), .B2(new_n916), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n942), .A2(G116), .A3(new_n218), .A4(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT36), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n220), .A2(G77), .A3(new_n324), .A4(new_n325), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(G50), .B2(new_n226), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(G1), .A3(new_n622), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n941), .A2(new_n945), .A3(new_n948), .ZN(G367));
  AOI21_X1  g0749(.A(new_n775), .B1(new_n699), .B2(new_n531), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n765), .A2(new_n241), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n757), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n358), .B1(new_n801), .B2(new_n856), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n785), .A2(new_n802), .B1(new_n202), .B2(new_n780), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(G50), .C2(new_n809), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n805), .A2(new_n857), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n790), .A2(new_n226), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(G143), .C2(new_n786), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n955), .B(new_n959), .C1(new_n806), .C2(new_n797), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n958), .A2(KEYINPUT109), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT46), .B1(new_n798), .B2(G116), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n785), .A2(new_n815), .B1(new_n481), .B2(new_n780), .ZN(new_n963));
  XOR2_X1   g0763(.A(KEYINPUT107), .B(G311), .Z(new_n964));
  OAI22_X1  g0764(.A1(new_n787), .A2(new_n964), .B1(new_n482), .B2(new_n790), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(G283), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n805), .A2(new_n812), .B1(new_n808), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT108), .B(G317), .Z(new_n969));
  AOI211_X1 g0769(.A(new_n358), .B(new_n968), .C1(new_n845), .C2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n798), .A2(KEYINPUT46), .A3(G116), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n966), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n960), .A2(new_n961), .B1(new_n962), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT47), .Z(new_n974));
  OR2_X1    g0774(.A1(new_n689), .A2(new_n534), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(new_n552), .Z(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n952), .B1(new_n864), .B2(new_n974), .C1(new_n977), .C2(new_n777), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n696), .A2(G330), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n686), .A3(new_n687), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n980), .A2(new_n697), .A3(new_n692), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n692), .B1(new_n980), .B2(new_n697), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n750), .A2(KEYINPUT106), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n693), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n681), .A2(new_n659), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n656), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n681), .A2(new_n478), .A3(new_n659), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(KEYINPUT44), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  INV_X1    g0791(.A(new_n989), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n693), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n693), .A2(new_n992), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n994), .A2(new_n999), .A3(new_n697), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n697), .B1(new_n994), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n983), .A2(new_n725), .A3(new_n748), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n984), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n750), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n700), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n754), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT43), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n976), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n989), .B(KEYINPUT105), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n500), .B1(new_n1013), .B2(new_n650), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n689), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n992), .A2(new_n688), .A3(new_n692), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT42), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1012), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(KEYINPUT43), .B2(new_n977), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1015), .A2(new_n1018), .A3(new_n1011), .A4(new_n976), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1013), .A2(new_n697), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1022), .B(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n978), .B1(new_n1010), .B2(new_n1025), .ZN(G387));
  NAND3_X1  g0826(.A1(new_n686), .A2(new_n687), .A3(new_n773), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n238), .A2(G45), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1028), .A2(new_n766), .B1(new_n703), .B2(new_n762), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n253), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT50), .B1(new_n253), .B2(G50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n703), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1029), .A2(new_n1033), .B1(new_n482), .B2(new_n699), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n758), .B1(new_n1034), .B2(new_n775), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n805), .A2(new_n258), .B1(new_n801), .B2(new_n857), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n290), .B(new_n1036), .C1(G68), .C2(new_n809), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n798), .A2(G77), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n791), .A2(new_n531), .B1(new_n817), .B2(G97), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n253), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G159), .A2(new_n786), .B1(new_n784), .B2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n844), .A2(new_n969), .B1(new_n809), .B2(G303), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n787), .B2(new_n823), .C1(new_n785), .C2(new_n964), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n798), .A2(G294), .B1(G283), .B2(new_n791), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n290), .B1(new_n801), .B2(new_n814), .C1(new_n573), .C2(new_n780), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1042), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1035), .B1(new_n1055), .B2(new_n770), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n983), .A2(new_n754), .B1(new_n1027), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1003), .A2(KEYINPUT110), .A3(new_n700), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n750), .B2(new_n983), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT110), .B1(new_n1003), .B2(new_n700), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(G393));
  INV_X1    g0861(.A(new_n1003), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1006), .B(new_n700), .C1(new_n1062), .C2(new_n1002), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1002), .A2(new_n754), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1013), .A2(new_n773), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n246), .A2(new_n765), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n775), .B1(G97), .B2(new_n699), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n757), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n787), .A2(new_n857), .B1(new_n802), .B2(new_n805), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT111), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  INV_X1    g0871(.A(G143), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n358), .B1(new_n801), .B2(new_n1072), .C1(new_n253), .C2(new_n808), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n791), .A2(G77), .B1(new_n817), .B2(G87), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n258), .B2(new_n785), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(G68), .C2(new_n798), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G317), .A2(new_n786), .B1(new_n844), .B2(G311), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT52), .Z(new_n1078));
  OAI221_X1 g0878(.A(new_n290), .B1(new_n801), .B2(new_n823), .C1(new_n815), .C2(new_n808), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n781), .B1(G116), .B2(new_n791), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n812), .B2(new_n785), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(G283), .C2(new_n798), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1071), .A2(new_n1076), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1065), .B(new_n1068), .C1(new_n864), .C2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1064), .A2(KEYINPUT112), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT112), .B1(new_n1064), .B2(new_n1084), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1063), .B1(new_n1086), .B2(new_n1087), .ZN(G390));
  OAI21_X1  g0888(.A(new_n929), .B1(new_n909), .B2(new_n928), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n771), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n757), .B1(new_n253), .B2(new_n842), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n799), .A2(new_n290), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT114), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G97), .A2(new_n809), .B1(new_n845), .B2(G294), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n573), .B2(new_n805), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n790), .A2(new_n202), .B1(new_n780), .B2(new_n226), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n785), .A2(new_n482), .B1(new_n787), .B2(new_n967), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n797), .A2(new_n857), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n290), .B1(new_n845), .B2(G125), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1102), .B1(new_n851), .B2(new_n805), .C1(new_n808), .C2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n786), .A2(G128), .B1(new_n817), .B2(G50), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n856), .B2(new_n785), .C1(new_n802), .C2(new_n790), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1101), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1098), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1090), .B(new_n1091), .C1(new_n864), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n871), .A2(new_n874), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n835), .B1(new_n922), .B2(new_n722), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n933), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n898), .A2(KEYINPUT38), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n931), .B1(new_n1113), .B2(new_n894), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n908), .A2(KEYINPUT39), .A3(new_n894), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT39), .B1(new_n1113), .B2(new_n894), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1116), .A2(new_n1117), .B1(new_n935), .B2(new_n931), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1110), .A2(G330), .A3(new_n747), .A4(new_n837), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n838), .A2(new_n934), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1110), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n930), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1089), .A2(new_n1123), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n901), .A2(G330), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n875), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1120), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1109), .B1(new_n1127), .B2(new_n753), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n924), .A2(new_n926), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n459), .A2(new_n1125), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n901), .A2(G330), .A3(new_n837), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1122), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n837), .B1(new_n720), .B2(new_n723), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n934), .A4(new_n1119), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n747), .A2(G330), .A3(new_n837), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1125), .A2(new_n875), .B1(new_n1135), .B2(new_n1122), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1121), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1129), .A2(new_n647), .A3(new_n1130), .A4(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1138), .A2(new_n1127), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n701), .B1(new_n1138), .B2(new_n1127), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1128), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(new_n1130), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n646), .B(new_n1143), .C1(new_n924), .C2(new_n926), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1137), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1127), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n938), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n267), .A2(new_n679), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n306), .A2(new_n309), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n306), .B2(new_n309), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1153), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n1151), .A3(new_n1148), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n875), .A2(new_n901), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT40), .B1(new_n908), .B2(new_n894), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1159), .A2(new_n1160), .B1(new_n902), .B2(KEYINPUT40), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1158), .B1(new_n1161), .B2(new_n870), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n912), .A2(G330), .A3(new_n1157), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1147), .B1(new_n1164), .B2(KEYINPUT118), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT118), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1166), .B(new_n938), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1146), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1157), .B1(new_n912), .B2(G330), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n870), .B(new_n1158), .C1(new_n903), .C2(new_n911), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1147), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1162), .A2(new_n938), .A3(new_n1163), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1169), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n701), .B1(new_n1175), .B2(new_n1146), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1170), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1158), .A2(new_n771), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n758), .B1(G50), .B2(new_n843), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n358), .A2(G41), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G50), .B(new_n1180), .C1(new_n284), .C2(new_n272), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n817), .A2(G58), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n845), .A2(G283), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1038), .A2(new_n1182), .A3(new_n1180), .A4(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT115), .Z(new_n1185));
  NOR2_X1   g0985(.A1(new_n805), .A2(new_n482), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT116), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1186), .A2(new_n1187), .B1(new_n784), .B2(G97), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n1187), .B2(new_n1186), .C1(new_n573), .C2(new_n787), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n957), .B(new_n1189), .C1(new_n531), .C2(new_n809), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1181), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n808), .A2(new_n856), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n785), .A2(new_n851), .B1(new_n857), .B2(new_n790), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(G125), .C2(new_n786), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1103), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n798), .A2(new_n1197), .B1(G128), .B2(new_n844), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT117), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1196), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n817), .A2(G159), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G33), .B(G41), .C1(new_n845), .C2(G124), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1193), .B(new_n1207), .C1(new_n1192), .C2(new_n1191), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1179), .B1(new_n1208), .B2(new_n770), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1178), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n754), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1177), .A2(new_n1213), .ZN(G375));
  NAND2_X1  g1014(.A1(new_n1137), .A2(new_n754), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1110), .A2(new_n772), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT119), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n757), .B1(new_n226), .B2(new_n842), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n805), .A2(new_n856), .B1(new_n808), .B2(new_n857), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n290), .B(new_n1219), .C1(G128), .C2(new_n845), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n798), .A2(G159), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n791), .A2(G50), .B1(new_n817), .B2(G58), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G132), .A2(new_n786), .B1(new_n784), .B2(new_n1197), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n805), .A2(new_n967), .B1(new_n801), .B2(new_n812), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n358), .B(new_n1225), .C1(G107), .C2(new_n809), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n798), .A2(G97), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n791), .A2(new_n531), .B1(new_n817), .B2(G77), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G116), .A2(new_n784), .B1(new_n786), .B2(G294), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1217), .B(new_n1218), .C1(new_n864), .C2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1215), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1008), .B1(new_n1144), .B2(new_n1137), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n458), .B1(new_n713), .B2(new_n715), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n925), .B1(new_n1235), .B2(new_n724), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n919), .A2(KEYINPUT103), .A3(new_n923), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n647), .B(new_n1130), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1145), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1233), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G381));
  INV_X1    g1041(.A(new_n1087), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1002), .A2(new_n1062), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(new_n701), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1242), .A2(new_n1085), .B1(new_n1244), .B2(new_n1006), .ZN(new_n1245));
  INV_X1    g1045(.A(G384), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G393), .A2(G396), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(new_n1247), .A2(G387), .A3(G381), .A4(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT120), .Z(new_n1250));
  NAND3_X1  g1050(.A1(new_n1177), .A2(new_n1141), .A3(new_n1213), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(G407));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G343), .C2(new_n1251), .ZN(G409));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G387), .B2(new_n1245), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(G393), .B(new_n830), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G387), .A2(new_n1245), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1022), .B(new_n1023), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1008), .B1(new_n1006), .B2(new_n750), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n754), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G390), .B1(new_n1262), .B2(new_n978), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n1256), .A2(new_n1258), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G387), .A2(new_n1245), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n978), .A3(G390), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1233), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT122), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT60), .B1(new_n1238), .B2(new_n1145), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1138), .A2(new_n700), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1238), .A2(new_n1145), .A3(KEYINPUT60), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1270), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1144), .B2(new_n1137), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n701), .B1(new_n1144), .B2(new_n1137), .ZN(new_n1278));
  AND4_X1   g1078(.A1(new_n1270), .A2(new_n1277), .A3(new_n1278), .A4(new_n1274), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1269), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1274), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT122), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1273), .A2(new_n1270), .A3(new_n1274), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1288), .A2(KEYINPUT123), .A3(new_n1246), .A4(new_n1269), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1141), .B1(new_n1177), .B2(new_n1213), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n754), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT121), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1210), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n753), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT121), .B1(new_n1296), .B2(new_n1211), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1146), .B(new_n1009), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1295), .A2(new_n1141), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G343), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(G213), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1291), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1290), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT124), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT124), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1290), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT62), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT61), .B1(new_n1304), .B2(KEYINPUT62), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1300), .A2(G213), .A3(G2897), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1290), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1303), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1310), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1283), .A2(new_n1289), .A3(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1311), .A2(new_n1312), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1309), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1268), .B1(new_n1308), .B2(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1303), .B(KEYINPUT125), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1305), .A2(new_n1320), .A3(new_n1307), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1304), .A2(new_n1320), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1264), .A2(new_n1323), .A3(new_n1267), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1319), .A2(new_n1321), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1317), .A2(new_n1326), .ZN(G405));
  NAND3_X1  g1127(.A1(new_n1268), .A2(new_n1289), .A3(new_n1283), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1264), .A2(new_n1267), .A3(new_n1290), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1330), .B1(new_n1252), .B2(new_n1291), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1291), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1328), .A2(new_n1251), .A3(new_n1332), .A4(new_n1329), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(G402));
endmodule


