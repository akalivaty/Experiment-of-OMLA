

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U551 ( .A1(G160), .A2(G40), .ZN(n780) );
  XOR2_X2 U552 ( .A(KEYINPUT17), .B(n520), .Z(n893) );
  XNOR2_X1 U553 ( .A(n733), .B(KEYINPUT102), .ZN(n748) );
  AND2_X1 U554 ( .A1(n782), .A2(n780), .ZN(n713) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n782) );
  XNOR2_X1 U556 ( .A(n687), .B(KEYINPUT97), .ZN(n688) );
  XNOR2_X1 U557 ( .A(n689), .B(n688), .ZN(n691) );
  NOR2_X1 U558 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X2 U559 ( .A1(G2105), .A2(n517), .ZN(n892) );
  NOR2_X1 U560 ( .A1(G651), .A2(n651), .ZN(n656) );
  NOR2_X1 U561 ( .A1(n526), .A2(n525), .ZN(G164) );
  INV_X1 U562 ( .A(G2104), .ZN(n517) );
  INV_X1 U563 ( .A(G2105), .ZN(n521) );
  NOR2_X2 U564 ( .A1(n517), .A2(n521), .ZN(n888) );
  NAND2_X1 U565 ( .A1(n888), .A2(G114), .ZN(n516) );
  XNOR2_X1 U566 ( .A(n516), .B(KEYINPUT88), .ZN(n519) );
  NAND2_X1 U567 ( .A1(G102), .A2(n892), .ZN(n518) );
  NAND2_X1 U568 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  NAND2_X1 U570 ( .A1(G138), .A2(n893), .ZN(n524) );
  NOR2_X1 U571 ( .A1(n521), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U572 ( .A(n522), .B(KEYINPUT64), .ZN(n889) );
  NAND2_X1 U573 ( .A1(G126), .A2(n889), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U575 ( .A1(G101), .A2(n892), .ZN(n527) );
  XNOR2_X1 U576 ( .A(n527), .B(KEYINPUT65), .ZN(n528) );
  XNOR2_X1 U577 ( .A(n528), .B(KEYINPUT23), .ZN(n530) );
  NAND2_X1 U578 ( .A1(G113), .A2(n888), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U580 ( .A1(G137), .A2(n893), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G125), .A2(n889), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X2 U583 ( .A1(n534), .A2(n533), .ZN(G160) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U585 ( .A1(n642), .A2(G85), .ZN(n536) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n651) );
  XOR2_X1 U587 ( .A(G651), .B(KEYINPUT66), .Z(n537) );
  NOR2_X1 U588 ( .A1(n651), .A2(n537), .ZN(n645) );
  NAND2_X1 U589 ( .A1(G72), .A2(n645), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n543) );
  NAND2_X1 U591 ( .A1(n656), .A2(G47), .ZN(n541) );
  NOR2_X1 U592 ( .A1(G543), .A2(n537), .ZN(n538) );
  XNOR2_X1 U593 ( .A(n538), .B(KEYINPUT1), .ZN(n539) );
  XNOR2_X1 U594 ( .A(KEYINPUT67), .B(n539), .ZN(n655) );
  NAND2_X1 U595 ( .A1(G60), .A2(n655), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U597 ( .A1(n543), .A2(n542), .ZN(G290) );
  XOR2_X1 U598 ( .A(KEYINPUT109), .B(G2435), .Z(n545) );
  XNOR2_X1 U599 ( .A(G2430), .B(G2438), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n545), .B(n544), .ZN(n552) );
  XOR2_X1 U601 ( .A(G2446), .B(G2454), .Z(n547) );
  XNOR2_X1 U602 ( .A(G2451), .B(G2443), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U604 ( .A(n548), .B(G2427), .Z(n550) );
  XNOR2_X1 U605 ( .A(G1341), .B(G1348), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n552), .B(n551), .ZN(n553) );
  AND2_X1 U608 ( .A1(n553), .A2(G14), .ZN(G401) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G120), .ZN(G236) );
  INV_X1 U613 ( .A(G69), .ZN(G235) );
  NAND2_X1 U614 ( .A1(G64), .A2(n655), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n554), .B(KEYINPUT68), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G52), .A2(n656), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT69), .B(n557), .Z(n563) );
  NAND2_X1 U619 ( .A1(n642), .A2(G90), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT70), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G77), .A2(n645), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U624 ( .A1(n563), .A2(n562), .ZN(G171) );
  NAND2_X1 U625 ( .A1(n656), .A2(G51), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT75), .B(n564), .Z(n566) );
  NAND2_X1 U627 ( .A1(G63), .A2(n655), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT6), .B(n567), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G89), .A2(n642), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(KEYINPUT74), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT4), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G76), .A2(n645), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U635 ( .A(n572), .B(KEYINPUT5), .Z(n573) );
  NOR2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT76), .B(n575), .Z(n576) );
  XNOR2_X1 U638 ( .A(KEYINPUT7), .B(n576), .ZN(G168) );
  XOR2_X1 U639 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U640 ( .A1(G94), .A2(G452), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT71), .ZN(G173) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U644 ( .A(G223), .ZN(n835) );
  NAND2_X1 U645 ( .A1(n835), .A2(G567), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(n579), .Z(G234) );
  NAND2_X1 U647 ( .A1(n642), .A2(G81), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT12), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G68), .A2(n645), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n583), .Z(n587) );
  NAND2_X1 U652 ( .A1(n655), .A2(G56), .ZN(n584) );
  XNOR2_X1 U653 ( .A(n584), .B(KEYINPUT14), .ZN(n585) );
  XNOR2_X1 U654 ( .A(n585), .B(KEYINPUT73), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n656), .A2(G43), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n942) );
  INV_X1 U658 ( .A(G860), .ZN(n609) );
  OR2_X1 U659 ( .A1(n942), .A2(n609), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n642), .A2(G92), .ZN(n591) );
  NAND2_X1 U663 ( .A1(G79), .A2(n645), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n656), .A2(G54), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G66), .A2(n655), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT15), .B(n596), .Z(n941) );
  OR2_X1 U670 ( .A1(n941), .A2(G868), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G78), .A2(n645), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G65), .A2(n655), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n642), .A2(G91), .ZN(n601) );
  XOR2_X1 U676 ( .A(KEYINPUT72), .B(n601), .Z(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n656), .A2(G53), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G299) );
  INV_X1 U680 ( .A(G868), .ZN(n668) );
  NOR2_X1 U681 ( .A1(G286), .A2(n668), .ZN(n606) );
  XOR2_X1 U682 ( .A(KEYINPUT77), .B(n606), .Z(n608) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n610), .A2(n941), .ZN(n611) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n942), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G868), .A2(n941), .ZN(n612) );
  NOR2_X1 U690 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U692 ( .A(KEYINPUT78), .B(n615), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G111), .A2(n888), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G99), .A2(n892), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n889), .A2(G123), .ZN(n618) );
  XOR2_X1 U697 ( .A(KEYINPUT18), .B(n618), .Z(n619) );
  NOR2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n893), .A2(G135), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n999) );
  XOR2_X1 U701 ( .A(n999), .B(G2096), .Z(n624) );
  XNOR2_X1 U702 ( .A(G2100), .B(KEYINPUT79), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G559), .A2(n941), .ZN(n625) );
  XOR2_X1 U705 ( .A(n942), .B(n625), .Z(n666) );
  XOR2_X1 U706 ( .A(n666), .B(KEYINPUT80), .Z(n626) );
  NOR2_X1 U707 ( .A1(G860), .A2(n626), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT82), .B(n627), .Z(n635) );
  NAND2_X1 U709 ( .A1(n642), .A2(G93), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G80), .A2(n645), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G55), .A2(n656), .ZN(n630) );
  XNOR2_X1 U713 ( .A(KEYINPUT81), .B(n630), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G67), .A2(n655), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n669) );
  XNOR2_X1 U717 ( .A(n635), .B(n669), .ZN(G145) );
  NAND2_X1 U718 ( .A1(n642), .A2(G88), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G75), .A2(n645), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n656), .A2(G50), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G62), .A2(n655), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U724 ( .A1(n641), .A2(n640), .ZN(G166) );
  NAND2_X1 U725 ( .A1(G86), .A2(n642), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G48), .A2(n656), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n645), .A2(G73), .ZN(n646) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G61), .A2(n655), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G87), .A2(n651), .ZN(n653) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U737 ( .A1(G49), .A2(n656), .ZN(n657) );
  XOR2_X1 U738 ( .A(KEYINPUT83), .B(n657), .Z(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(G288) );
  INV_X1 U740 ( .A(G299), .ZN(n694) );
  XNOR2_X1 U741 ( .A(G166), .B(n694), .ZN(n665) );
  XOR2_X1 U742 ( .A(G290), .B(G305), .Z(n660) );
  XNOR2_X1 U743 ( .A(n669), .B(n660), .ZN(n661) );
  XNOR2_X1 U744 ( .A(KEYINPUT84), .B(n661), .ZN(n663) );
  XNOR2_X1 U745 ( .A(G288), .B(KEYINPUT19), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n665), .B(n664), .ZN(n841) );
  XOR2_X1 U748 ( .A(n841), .B(n666), .Z(n667) );
  NOR2_X1 U749 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U750 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U751 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XNOR2_X1 U753 ( .A(n672), .B(KEYINPUT20), .ZN(n673) );
  XNOR2_X1 U754 ( .A(n673), .B(KEYINPUT85), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G235), .A2(G236), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G108), .A2(n677), .ZN(n678) );
  NOR2_X1 U761 ( .A1(n678), .A2(G237), .ZN(n679) );
  XNOR2_X1 U762 ( .A(n679), .B(KEYINPUT87), .ZN(n839) );
  NAND2_X1 U763 ( .A1(n839), .A2(G567), .ZN(n685) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U766 ( .A1(G218), .A2(n681), .ZN(n682) );
  XNOR2_X1 U767 ( .A(KEYINPUT86), .B(n682), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n683), .A2(G96), .ZN(n840) );
  NAND2_X1 U769 ( .A1(n840), .A2(G2106), .ZN(n684) );
  NAND2_X1 U770 ( .A1(n685), .A2(n684), .ZN(n913) );
  NAND2_X1 U771 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U772 ( .A1(n913), .A2(n686), .ZN(n838) );
  NAND2_X1 U773 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U775 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n834) );
  XNOR2_X1 U776 ( .A(n713), .B(KEYINPUT96), .ZN(n711) );
  NAND2_X1 U777 ( .A1(G2072), .A2(n711), .ZN(n689) );
  XOR2_X1 U778 ( .A(KEYINPUT98), .B(KEYINPUT27), .Z(n687) );
  XNOR2_X1 U779 ( .A(G1956), .B(KEYINPUT99), .ZN(n962) );
  NOR2_X1 U780 ( .A1(n711), .A2(n962), .ZN(n690) );
  NOR2_X1 U781 ( .A1(n691), .A2(n690), .ZN(n693) );
  NOR2_X1 U782 ( .A1(n694), .A2(n693), .ZN(n692) );
  XOR2_X1 U783 ( .A(n692), .B(KEYINPUT28), .Z(n709) );
  NAND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n707) );
  XNOR2_X1 U785 ( .A(G1996), .B(KEYINPUT100), .ZN(n917) );
  NAND2_X1 U786 ( .A1(n917), .A2(n713), .ZN(n695) );
  XNOR2_X1 U787 ( .A(n695), .B(KEYINPUT26), .ZN(n697) );
  NAND2_X1 U788 ( .A1(n782), .A2(n780), .ZN(n737) );
  NAND2_X1 U789 ( .A1(n737), .A2(G1341), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n942), .A2(n698), .ZN(n699) );
  OR2_X1 U792 ( .A1(n941), .A2(n699), .ZN(n705) );
  NAND2_X1 U793 ( .A1(n941), .A2(n699), .ZN(n703) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n711), .ZN(n701) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n737), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U801 ( .A(n710), .B(KEYINPUT29), .ZN(n717) );
  XOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .Z(n918) );
  INV_X1 U803 ( .A(n711), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n918), .A2(n712), .ZN(n715) );
  NOR2_X1 U805 ( .A1(n713), .A2(G1961), .ZN(n714) );
  NOR2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n722) );
  NOR2_X1 U807 ( .A1(G301), .A2(n722), .ZN(n716) );
  NOR2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n727) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n737), .ZN(n730) );
  NAND2_X1 U810 ( .A1(G8), .A2(n737), .ZN(n736) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n736), .ZN(n718) );
  XNOR2_X1 U812 ( .A(KEYINPUT95), .B(n718), .ZN(n729) );
  NAND2_X1 U813 ( .A1(G8), .A2(n729), .ZN(n719) );
  NOR2_X1 U814 ( .A1(n730), .A2(n719), .ZN(n720) );
  XOR2_X1 U815 ( .A(KEYINPUT30), .B(n720), .Z(n721) );
  NOR2_X1 U816 ( .A1(G168), .A2(n721), .ZN(n724) );
  AND2_X1 U817 ( .A1(G301), .A2(n722), .ZN(n723) );
  NOR2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U819 ( .A(n725), .B(KEYINPUT31), .ZN(n726) );
  NOR2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U821 ( .A(n728), .B(KEYINPUT101), .ZN(n735) );
  AND2_X1 U822 ( .A1(n735), .A2(n729), .ZN(n732) );
  NAND2_X1 U823 ( .A1(G8), .A2(n730), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n733) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n744) );
  INV_X1 U827 ( .A(G8), .ZN(n742) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n736), .ZN(n739) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n737), .ZN(n738) );
  NOR2_X1 U830 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  AND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n746) );
  XOR2_X1 U834 ( .A(KEYINPUT103), .B(KEYINPUT32), .Z(n745) );
  XNOR2_X1 U835 ( .A(n746), .B(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n808) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n756), .A2(n749), .ZN(n950) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n750) );
  AND2_X1 U841 ( .A1(n950), .A2(n750), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n808), .A2(n751), .ZN(n755) );
  INV_X1 U843 ( .A(n736), .ZN(n752) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n949) );
  AND2_X1 U845 ( .A1(n752), .A2(n949), .ZN(n753) );
  OR2_X1 U846 ( .A1(KEYINPUT33), .A2(n753), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n760) );
  NAND2_X1 U848 ( .A1(KEYINPUT33), .A2(n756), .ZN(n757) );
  NOR2_X1 U849 ( .A1(n736), .A2(n757), .ZN(n758) );
  XNOR2_X1 U850 ( .A(n758), .B(KEYINPUT104), .ZN(n759) );
  XOR2_X1 U851 ( .A(KEYINPUT105), .B(n761), .Z(n799) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n937) );
  NAND2_X1 U853 ( .A1(G107), .A2(n888), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G119), .A2(n889), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n768) );
  NAND2_X1 U856 ( .A1(G95), .A2(n892), .ZN(n765) );
  NAND2_X1 U857 ( .A1(G131), .A2(n893), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U859 ( .A(KEYINPUT91), .B(n766), .Z(n767) );
  OR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n884) );
  AND2_X1 U861 ( .A1(n884), .A2(G1991), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G117), .A2(n888), .ZN(n770) );
  NAND2_X1 U863 ( .A1(G129), .A2(n889), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n775) );
  XOR2_X1 U865 ( .A(KEYINPUT38), .B(KEYINPUT93), .Z(n772) );
  NAND2_X1 U866 ( .A1(G105), .A2(n892), .ZN(n771) );
  XNOR2_X1 U867 ( .A(n772), .B(n771), .ZN(n773) );
  XOR2_X1 U868 ( .A(KEYINPUT92), .B(n773), .Z(n774) );
  NOR2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n893), .A2(G141), .ZN(n776) );
  NAND2_X1 U871 ( .A1(n777), .A2(n776), .ZN(n880) );
  AND2_X1 U872 ( .A1(n880), .A2(G1996), .ZN(n778) );
  NOR2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n995) );
  INV_X1 U874 ( .A(n780), .ZN(n781) );
  NOR2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n829) );
  INV_X1 U876 ( .A(n829), .ZN(n783) );
  NOR2_X1 U877 ( .A1(n995), .A2(n783), .ZN(n821) );
  INV_X1 U878 ( .A(n821), .ZN(n795) );
  XNOR2_X1 U879 ( .A(KEYINPUT37), .B(G2067), .ZN(n827) );
  NAND2_X1 U880 ( .A1(n893), .A2(G140), .ZN(n784) );
  XOR2_X1 U881 ( .A(KEYINPUT89), .B(n784), .Z(n786) );
  NAND2_X1 U882 ( .A1(n892), .A2(G104), .ZN(n785) );
  NAND2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n788) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(KEYINPUT90), .ZN(n787) );
  XNOR2_X1 U885 ( .A(n788), .B(n787), .ZN(n793) );
  NAND2_X1 U886 ( .A1(G116), .A2(n888), .ZN(n790) );
  NAND2_X1 U887 ( .A1(G128), .A2(n889), .ZN(n789) );
  NAND2_X1 U888 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U889 ( .A(KEYINPUT35), .B(n791), .Z(n792) );
  NOR2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U891 ( .A(KEYINPUT36), .B(n794), .ZN(n885) );
  NOR2_X1 U892 ( .A1(n827), .A2(n885), .ZN(n998) );
  NAND2_X1 U893 ( .A1(n829), .A2(n998), .ZN(n825) );
  NAND2_X1 U894 ( .A1(n795), .A2(n825), .ZN(n813) );
  INV_X1 U895 ( .A(n813), .ZN(n796) );
  AND2_X1 U896 ( .A1(n937), .A2(n796), .ZN(n797) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n948) );
  NAND2_X1 U898 ( .A1(n948), .A2(n829), .ZN(n800) );
  AND2_X1 U899 ( .A1(n797), .A2(n800), .ZN(n798) );
  NAND2_X1 U900 ( .A1(n799), .A2(n798), .ZN(n817) );
  INV_X1 U901 ( .A(n800), .ZN(n815) );
  NOR2_X1 U902 ( .A1(G2090), .A2(G303), .ZN(n801) );
  NAND2_X1 U903 ( .A1(G8), .A2(n801), .ZN(n806) );
  NOR2_X1 U904 ( .A1(G1981), .A2(G305), .ZN(n802) );
  XOR2_X1 U905 ( .A(n802), .B(KEYINPUT94), .Z(n803) );
  XNOR2_X1 U906 ( .A(KEYINPUT24), .B(n803), .ZN(n804) );
  NOR2_X1 U907 ( .A1(n736), .A2(n804), .ZN(n809) );
  INV_X1 U908 ( .A(n809), .ZN(n805) );
  AND2_X1 U909 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U910 ( .A1(n808), .A2(n807), .ZN(n811) );
  OR2_X1 U911 ( .A1(n809), .A2(n736), .ZN(n810) );
  NAND2_X1 U912 ( .A1(n811), .A2(n810), .ZN(n812) );
  OR2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n814) );
  OR2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  AND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n832) );
  XOR2_X1 U916 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n824) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n880), .ZN(n992) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n884), .ZN(n1002) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n818) );
  XNOR2_X1 U920 ( .A(KEYINPUT106), .B(n818), .ZN(n819) );
  NOR2_X1 U921 ( .A1(n1002), .A2(n819), .ZN(n820) );
  NOR2_X1 U922 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U923 ( .A1(n992), .A2(n822), .ZN(n823) );
  XNOR2_X1 U924 ( .A(n824), .B(n823), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n827), .A2(n885), .ZN(n1006) );
  NAND2_X1 U927 ( .A1(n828), .A2(n1006), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U933 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G188) );
  XOR2_X1 U936 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  NOR2_X1 U939 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U941 ( .A(n942), .B(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(G171), .B(n941), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U944 ( .A(n844), .B(G286), .Z(n845) );
  NOR2_X1 U945 ( .A1(G37), .A2(n845), .ZN(G397) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2072), .B(G2678), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n848), .B(KEYINPUT110), .Z(n850) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2100), .Z(n852) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1976), .B(G1966), .Z(n856) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1971), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U959 ( .A(G1981), .B(G1956), .Z(n858) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U962 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U963 ( .A(G2474), .B(KEYINPUT41), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n864) );
  XOR2_X1 U965 ( .A(G1961), .B(KEYINPUT111), .Z(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G112), .A2(n888), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G136), .A2(n893), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n889), .A2(G124), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n867), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G100), .A2(n892), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n868), .B(KEYINPUT112), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G103), .A2(n892), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G139), .A2(n893), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G115), .A2(n888), .ZN(n876) );
  NAND2_X1 U980 ( .A1(G127), .A2(n889), .ZN(n875) );
  NAND2_X1 U981 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U983 ( .A1(n879), .A2(n878), .ZN(n1009) );
  XNOR2_X1 U984 ( .A(n999), .B(G162), .ZN(n882) );
  XOR2_X1 U985 ( .A(G164), .B(n880), .Z(n881) );
  XNOR2_X1 U986 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U987 ( .A(n1009), .B(n883), .ZN(n887) );
  XOR2_X1 U988 ( .A(n885), .B(n884), .Z(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n905) );
  XOR2_X1 U990 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n902) );
  NAND2_X1 U991 ( .A1(G118), .A2(n888), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G106), .A2(n892), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G142), .A2(n893), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U997 ( .A(KEYINPUT45), .B(n896), .ZN(n897) );
  XNOR2_X1 U998 ( .A(KEYINPUT113), .B(n897), .ZN(n898) );
  NOR2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n900), .B(KEYINPUT48), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(G160), .B(n903), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n906), .ZN(G395) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n913), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1008 ( .A1(G397), .A2(n908), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n911) );
  NOR2_X1 U1010 ( .A1(n911), .A2(G395), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n912), .B(KEYINPUT115), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n913), .ZN(G319) );
  XOR2_X1 U1014 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n932) );
  XNOR2_X1 U1015 ( .A(G2090), .B(G35), .ZN(n927) );
  XOR2_X1 U1016 ( .A(G25), .B(G1991), .Z(n914) );
  NAND2_X1 U1017 ( .A1(n914), .A2(G28), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(G2067), .B(G26), .ZN(n916) );
  XNOR2_X1 U1019 ( .A(G33), .B(G2072), .ZN(n915) );
  NOR2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n917), .B(G32), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(G27), .B(n918), .ZN(n919) );
  NOR2_X1 U1023 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(KEYINPUT53), .B(n925), .ZN(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1028 ( .A(G2084), .B(G34), .Z(n928) );
  XNOR2_X1 U1029 ( .A(KEYINPUT54), .B(n928), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(n932), .B(n931), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(n933), .B(KEYINPUT55), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(G29), .A2(n934), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT123), .B(n935), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n936), .A2(G11), .ZN(n990) );
  XNOR2_X1 U1036 ( .A(G16), .B(KEYINPUT56), .ZN(n961) );
  XNOR2_X1 U1037 ( .A(G168), .B(G1966), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(n939), .B(KEYINPUT124), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT57), .B(n940), .ZN(n959) );
  XNOR2_X1 U1041 ( .A(n941), .B(G1348), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(n942), .B(G1341), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(G299), .B(G1956), .ZN(n943) );
  NOR2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n952) );
  AND2_X1 U1048 ( .A1(G303), .A2(G1971), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1050 ( .A(KEYINPUT125), .B(n953), .Z(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(G1961), .B(G301), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n988) );
  INV_X1 U1056 ( .A(G16), .ZN(n986) );
  XNOR2_X1 U1057 ( .A(G20), .B(n962), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G1341), .B(G19), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G1981), .B(G6), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1062 ( .A(KEYINPUT59), .B(G1348), .Z(n967) );
  XNOR2_X1 U1063 ( .A(G4), .B(n967), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1065 ( .A(KEYINPUT60), .B(n970), .Z(n972) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G21), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(KEYINPUT126), .B(n973), .ZN(n982) );
  XNOR2_X1 U1069 ( .A(G1961), .B(G5), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G1971), .B(G22), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G23), .B(G1976), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n977) );
  XOR2_X1 U1073 ( .A(G1986), .B(G24), .Z(n976) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(KEYINPUT58), .B(n978), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n983), .B(KEYINPUT61), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT127), .B(n984), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n1021) );
  XOR2_X1 U1083 ( .A(G2090), .B(G162), .Z(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1085 ( .A(KEYINPUT51), .B(n993), .Z(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT118), .B(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(G160), .B(G2084), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(KEYINPUT117), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1015) );
  XNOR2_X1 U1095 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1008), .B(KEYINPUT50), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(G2072), .B(n1009), .Z(n1011) );
  XOR2_X1 U1098 ( .A(G164), .B(G2078), .Z(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1016), .ZN(n1018) );
  INV_X1 U1103 ( .A(KEYINPUT55), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(G29), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

