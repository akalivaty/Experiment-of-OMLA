//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1039, new_n1040, new_n1041;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT73), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT73), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n208), .B(new_n202), .C1(new_n203), .C2(new_n204), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n206), .A2(new_n211), .A3(new_n207), .A4(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G226gat), .A2(G233gat), .ZN(new_n216));
  OR2_X1    g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT26), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n217), .A2(KEYINPUT26), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  OAI22_X1  g022(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(KEYINPUT27), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  AOI21_X1  g025(.A(G190gat), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n227), .B(KEYINPUT69), .C1(new_n226), .C2(new_n228), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n228), .A2(KEYINPUT28), .A3(new_n223), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n224), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT24), .ZN(new_n237));
  XOR2_X1   g036(.A(G183gat), .B(G190gat), .Z(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(KEYINPUT24), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT66), .B(KEYINPUT23), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n217), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n219), .B1(new_n217), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(KEYINPUT67), .B(new_n219), .C1(new_n217), .C2(new_n242), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n239), .A2(new_n241), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT25), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT65), .B(G176gat), .Z(new_n249));
  INV_X1    g048(.A(G169gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(KEYINPUT23), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n239), .A2(new_n251), .A3(new_n241), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n236), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT74), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT74), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n236), .B2(new_n254), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n216), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n216), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n255), .A2(KEYINPUT29), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n215), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n260), .A2(KEYINPUT29), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n256), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n215), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n255), .A2(new_n260), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G8gat), .B(G36gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n262), .A2(new_n271), .A3(new_n267), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(KEYINPUT30), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n262), .A2(new_n276), .A3(new_n271), .A4(new_n267), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT75), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(G155gat), .A3(G162gat), .ZN(new_n282));
  INV_X1    g081(.A(G155gat), .ZN(new_n283));
  INV_X1    g082(.A(G162gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n280), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G141gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(G148gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n281), .A2(KEYINPUT2), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n289), .B2(G141gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n287), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n290), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n279), .B1(new_n285), .B2(KEYINPUT2), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n286), .A2(new_n293), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G127gat), .B(G134gat), .Z(new_n300));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301));
  INV_X1    g100(.A(G127gat), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n302), .A2(G134gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304));
  OAI221_X1 g103(.A(new_n300), .B1(new_n301), .B2(new_n303), .C1(KEYINPUT1), .C2(new_n304), .ZN(new_n305));
  OAI22_X1  g104(.A1(new_n304), .A2(KEYINPUT1), .B1(new_n303), .B2(new_n301), .ZN(new_n306));
  INV_X1    g105(.A(new_n300), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  OR3_X1    g108(.A1(new_n309), .A2(KEYINPUT80), .A3(KEYINPUT4), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT80), .B1(new_n309), .B2(KEYINPUT4), .ZN(new_n311));
  INV_X1    g110(.A(new_n299), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT71), .B1(new_n305), .B2(new_n308), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n308), .A3(KEYINPUT71), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n310), .B(new_n311), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G225gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n308), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n308), .A3(KEYINPUT77), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(KEYINPUT3), .B2(new_n312), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n299), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n299), .A2(new_n329), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n320), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n299), .B1(new_n323), .B2(new_n324), .ZN(new_n335));
  INV_X1    g134(.A(new_n309), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n320), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n337), .B2(KEYINPUT5), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n305), .A2(new_n308), .A3(KEYINPUT77), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT77), .B1(new_n305), .B2(new_n308), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n312), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n319), .B1(new_n341), .B2(new_n309), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n342), .A2(KEYINPUT81), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n333), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT0), .ZN(new_n347));
  XNOR2_X1  g146(.A(G57gat), .B(G85gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n316), .A2(new_n317), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n309), .A2(KEYINPUT4), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n351), .A2(KEYINPUT82), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(KEYINPUT82), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n343), .A3(new_n332), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n345), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT6), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n345), .A2(new_n355), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n349), .B1(new_n359), .B2(KEYINPUT90), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT81), .B1(new_n342), .B2(new_n343), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n334), .A3(KEYINPUT5), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n361), .A2(new_n362), .B1(new_n332), .B2(new_n318), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n354), .A2(new_n343), .A3(new_n332), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT90), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n358), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n349), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT6), .B(new_n369), .C1(new_n363), .C2(new_n364), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT84), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n359), .A2(new_n372), .A3(KEYINPUT6), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n278), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT93), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n254), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n234), .A2(new_n235), .ZN(new_n379));
  INV_X1    g178(.A(new_n224), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n315), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n313), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n236), .A2(new_n254), .B1(new_n382), .B2(new_n313), .ZN(new_n385));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT64), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT32), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G15gat), .B(G43gat), .Z(new_n392));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n388), .B(KEYINPUT32), .C1(new_n390), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n384), .A2(new_n385), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n386), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT34), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n387), .A2(KEYINPUT34), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n404), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n331), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(KEYINPUT86), .A3(new_n265), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n214), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n409), .B(new_n413), .C1(new_n215), .C2(KEYINPUT85), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n299), .B1(new_n414), .B2(new_n326), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT29), .B1(new_n328), .B2(new_n330), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n215), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n411), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G228gat), .ZN(new_n421));
  INV_X1    g220(.A(G233gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n215), .B1(new_n410), .B2(KEYINPUT87), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n418), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n424), .B1(new_n430), .B2(new_n312), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n420), .A2(new_n424), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(G22gat), .B1(new_n432), .B2(KEYINPUT88), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n424), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n431), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT88), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n408), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n410), .A2(new_n265), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n415), .B1(new_n440), .B2(new_n417), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n423), .B1(new_n441), .B2(new_n411), .ZN(new_n442));
  INV_X1    g241(.A(new_n431), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n425), .B2(new_n427), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n439), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n445), .A2(KEYINPUT89), .A3(G22gat), .A4(new_n436), .ZN(new_n446));
  XOR2_X1   g245(.A(G78gat), .B(G106gat), .Z(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G22gat), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n449), .B1(new_n432), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n438), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n435), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(G22gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n432), .A2(new_n450), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n449), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n407), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n278), .B(KEYINPUT93), .C1(new_n368), .C2(new_n374), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n377), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT35), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n451), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n450), .B1(new_n453), .B2(new_n439), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT89), .B1(new_n463), .B2(new_n436), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n456), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n398), .A2(new_n466), .A3(new_n404), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n404), .B1(new_n398), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(KEYINPUT35), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT36), .B1(new_n405), .B2(new_n406), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n452), .B(new_n456), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n278), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT6), .B1(new_n365), .B2(new_n349), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n477), .A2(KEYINPUT83), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n359), .A2(new_n369), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(KEYINPUT83), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n371), .A2(new_n373), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n360), .A2(new_n367), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n325), .A2(new_n331), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n319), .B1(new_n354), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n335), .A2(new_n320), .A3(new_n336), .ZN(new_n489));
  OR3_X1    g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n369), .B1(new_n487), .B2(new_n488), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n490), .A2(KEYINPUT40), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT40), .B1(new_n490), .B2(new_n491), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n485), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n485), .A2(new_n477), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n268), .A2(KEYINPUT37), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n271), .B1(new_n262), .B2(new_n267), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n271), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT38), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n496), .A2(new_n502), .A3(new_n482), .A4(new_n274), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n264), .A2(new_n266), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n215), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n259), .A2(new_n261), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n265), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT91), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n499), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n498), .B2(new_n500), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n504), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n500), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT38), .B1(new_n273), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n256), .A2(new_n258), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n260), .ZN(new_n519));
  INV_X1    g318(.A(new_n261), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI22_X1  g320(.A1(new_n521), .A2(new_n215), .B1(new_n510), .B2(KEYINPUT91), .ZN(new_n522));
  INV_X1    g321(.A(new_n511), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT37), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(KEYINPUT92), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n515), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n495), .B1(new_n503), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n472), .ZN(new_n528));
  INV_X1    g327(.A(new_n473), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n528), .A2(new_n529), .B1(new_n452), .B2(new_n456), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n461), .A2(new_n484), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT16), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(G1gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(G1gat), .B2(new_n533), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G8gat), .ZN(new_n537));
  INV_X1    g336(.A(G8gat), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n535), .B(new_n538), .C1(G1gat), .C2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT97), .A2(G71gat), .A3(G78gat), .ZN(new_n546));
  INV_X1    g345(.A(G71gat), .ZN(new_n547));
  INV_X1    g346(.A(G78gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT98), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(G57gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G64gat), .ZN(new_n555));
  INV_X1    g354(.A(G64gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G57gat), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n545), .A2(new_n549), .A3(KEYINPUT98), .A4(new_n546), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n549), .A2(new_n543), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT99), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT99), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n541), .B1(new_n542), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT103), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G127gat), .B(G155gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n573), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT102), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT101), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n577), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n574), .A2(new_n575), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n574), .B2(new_n575), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n587), .A2(KEYINPUT106), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT7), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(G85gat), .A3(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT104), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(KEYINPUT104), .A2(G92gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G99gat), .ZN(new_n600));
  INV_X1    g399(.A(G106gat), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT8), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n593), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G99gat), .B(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n593), .A2(new_n599), .A3(new_n604), .A4(new_n602), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n606), .A2(KEYINPUT105), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT105), .B1(new_n606), .B2(new_n607), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT15), .ZN(new_n611));
  NOR2_X1   g410(.A1(G43gat), .A2(G50gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G43gat), .A2(G50gat), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G29gat), .ZN(new_n616));
  INV_X1    g415(.A(G36gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT14), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT14), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(G29gat), .B2(G36gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(G29gat), .A2(G36gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(G43gat), .A2(G50gat), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT15), .B1(new_n624), .B2(new_n612), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n625), .A2(new_n620), .A3(new_n618), .A4(new_n621), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n614), .A2(new_n611), .ZN(new_n627));
  AND2_X1   g426(.A1(KEYINPUT94), .A2(G43gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(KEYINPUT94), .A2(G43gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G50gat), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n623), .B1(new_n626), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT95), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT17), .ZN(new_n635));
  INV_X1    g434(.A(new_n627), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT94), .B(G43gat), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(G50gat), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n625), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n634), .A2(new_n635), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n640), .B2(new_n623), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n615), .A2(new_n622), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT95), .B1(new_n645), .B2(new_n638), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT17), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n610), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT8), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(G99gat), .B2(G106gat), .ZN(new_n651));
  AND2_X1   g450(.A1(KEYINPUT104), .A2(G92gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(KEYINPUT104), .A2(G92gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n651), .B1(new_n654), .B2(new_n597), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n604), .B1(new_n655), .B2(new_n593), .ZN(new_n656));
  INV_X1    g455(.A(new_n607), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n649), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n606), .A2(KEYINPUT105), .A3(new_n607), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n646), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662));
  AND2_X1   g461(.A1(G232gat), .A2(G233gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n660), .A2(new_n661), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n588), .B1(new_n648), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G134gat), .B(G162gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n588), .B(new_n669), .C1(new_n648), .C2(new_n665), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n587), .A2(KEYINPUT106), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n664), .A2(new_n662), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n668), .B2(new_n670), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n586), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(G113gat), .B(G141gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G197gat), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT11), .B(G169gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT12), .ZN(new_n684));
  NAND2_X1  g483(.A1(G229gat), .A2(G233gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n540), .B1(new_n647), .B2(new_n643), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n540), .B1(new_n644), .B2(new_n646), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  AOI211_X1 g489(.A(new_n688), .B(new_n540), .C1(new_n647), .C2(new_n643), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT18), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT18), .B(new_n685), .C1(new_n690), .C2(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n661), .A2(new_n541), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n687), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n685), .B(KEYINPUT13), .Z(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND4_X1   g498(.A1(new_n684), .A2(new_n694), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n699), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n692), .B2(new_n693), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n684), .B1(new_n702), .B2(new_n695), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(G120gat), .B(G148gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(G176gat), .B(G204gat), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n705), .B(new_n706), .Z(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(G230gat), .A2(G233gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n561), .A2(new_n564), .A3(KEYINPUT10), .A4(new_n566), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT108), .B1(new_n660), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n711), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n659), .A4(new_n658), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n606), .A2(new_n607), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n567), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n555), .A2(new_n557), .ZN(new_n720));
  INV_X1    g519(.A(new_n553), .ZN(new_n721));
  AND4_X1   g520(.A1(new_n565), .A2(new_n720), .A3(new_n562), .A4(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n565), .B1(new_n558), .B2(new_n562), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n724), .A2(new_n561), .B1(new_n607), .B2(new_n606), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT107), .B(KEYINPUT10), .Z(new_n727));
  NAND3_X1  g526(.A1(new_n719), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n710), .B1(new_n716), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n718), .A2(new_n725), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n709), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n708), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n731), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n712), .A2(new_n715), .B1(new_n730), .B2(new_n727), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n733), .B(new_n707), .C1(new_n734), .C2(new_n710), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n732), .A2(KEYINPUT109), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT109), .B1(new_n732), .B2(new_n735), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n679), .A2(new_n704), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n532), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n481), .A2(new_n482), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT110), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g545(.A(KEYINPUT16), .B(G8gat), .Z(new_n747));
  AND3_X1   g546(.A1(new_n742), .A2(new_n476), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT42), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n742), .A2(new_n476), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT42), .B1(new_n751), .B2(new_n538), .ZN(new_n752));
  INV_X1    g551(.A(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n749), .B1(new_n748), .B2(KEYINPUT42), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(G1325gat));
  INV_X1    g555(.A(G15gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n407), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n528), .A2(new_n529), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n742), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n762), .B2(new_n757), .ZN(G1326gat));
  INV_X1    g562(.A(new_n465), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n742), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT43), .B(G22gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1327gat));
  AOI22_X1  g566(.A1(new_n460), .A2(new_n459), .B1(new_n527), .B2(new_n530), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n678), .B1(new_n768), .B2(new_n484), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n586), .A2(new_n740), .A3(new_n704), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n744), .A2(new_n616), .ZN(new_n773));
  OR3_X1    g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n532), .B2(new_n677), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n675), .B2(new_n676), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n668), .A2(new_n670), .ZN(new_n784));
  INV_X1    g583(.A(new_n673), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(KEYINPUT114), .A3(new_n674), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n780), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n768), .B2(new_n484), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n781), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n770), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n743), .B(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G29gat), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n774), .A2(new_n777), .A3(new_n775), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n795), .A3(new_n796), .ZN(G1328gat));
  NOR3_X1   g596(.A1(new_n771), .A2(G36gat), .A3(new_n278), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT46), .ZN(new_n799));
  OAI21_X1  g598(.A(G36gat), .B1(new_n792), .B2(new_n278), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1329gat));
  NOR2_X1   g600(.A1(new_n760), .A2(new_n630), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n791), .A2(new_n770), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n630), .B1(new_n771), .B2(new_n407), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n803), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1330gat));
  OAI211_X1 g608(.A(new_n764), .B(new_n770), .C1(new_n781), .C2(new_n790), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G50gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n769), .A2(new_n631), .A3(new_n764), .A4(new_n770), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT48), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n811), .B(new_n812), .C1(KEYINPUT115), .C2(KEYINPUT48), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1331gat));
  INV_X1    g617(.A(new_n740), .ZN(new_n819));
  INV_X1    g618(.A(new_n684), .ZN(new_n820));
  INV_X1    g619(.A(new_n685), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n644), .A2(new_n646), .A3(KEYINPUT17), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n635), .B1(new_n634), .B2(new_n642), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n541), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n634), .A2(new_n642), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT96), .B1(new_n825), .B2(new_n540), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n686), .A2(KEYINPUT96), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n821), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n699), .B1(new_n829), .B2(KEYINPUT18), .ZN(new_n830));
  INV_X1    g629(.A(new_n695), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n820), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n702), .A2(new_n684), .A3(new_n695), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n679), .A2(new_n819), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n532), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n794), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(new_n554), .ZN(G1332gat));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n278), .ZN(new_n839));
  NOR2_X1   g638(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n840));
  AND2_X1   g639(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n839), .B2(new_n840), .ZN(G1333gat));
  OAI21_X1  g642(.A(G71gat), .B1(new_n836), .B2(new_n760), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n758), .A2(new_n547), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n836), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g646(.A1(new_n836), .A2(new_n465), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n548), .ZN(G1335gat));
  NAND2_X1  g648(.A1(new_n704), .A2(new_n585), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT116), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n819), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n791), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G85gat), .B1(new_n854), .B2(new_n794), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n532), .A2(new_n677), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n852), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n769), .A2(KEYINPUT51), .A3(new_n851), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n819), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n597), .A3(new_n744), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n855), .A2(new_n861), .ZN(G1336gat));
  NOR2_X1   g661(.A1(new_n278), .A2(G92gat), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n819), .B(new_n864), .C1(new_n858), .C2(new_n859), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n476), .B(new_n853), .C1(new_n781), .C2(new_n790), .ZN(new_n866));
  INV_X1    g665(.A(new_n654), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT52), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n860), .A2(new_n863), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n866), .A2(new_n867), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n873), .ZN(G1337gat));
  OAI21_X1  g673(.A(G99gat), .B1(new_n854), .B2(new_n760), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n600), .A3(new_n758), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1338gat));
  XNOR2_X1  g676(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n465), .A2(G106gat), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n819), .B(new_n881), .C1(new_n858), .C2(new_n859), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n764), .B(new_n853), .C1(new_n781), .C2(new_n790), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(G106gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n860), .A2(new_n880), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(G106gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n878), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(G1339gat));
  AOI21_X1  g688(.A(new_n714), .B1(new_n610), .B2(new_n713), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n608), .A2(new_n711), .A3(new_n609), .A4(KEYINPUT108), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n728), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n709), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n716), .A2(new_n710), .A3(new_n728), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(KEYINPUT54), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n707), .B1(new_n729), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT55), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n735), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT55), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT54), .B1(new_n734), .B2(new_n710), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n716), .A2(new_n710), .A3(new_n728), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n892), .A2(new_n896), .A3(new_n709), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n708), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n900), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n834), .A2(new_n899), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n690), .A2(new_n691), .A3(new_n685), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n697), .A2(new_n698), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n683), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n833), .B(new_n910), .C1(new_n736), .C2(new_n738), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n788), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n783), .A2(new_n787), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n906), .A2(new_n735), .A3(new_n898), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n833), .A2(new_n910), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n585), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n819), .A2(new_n704), .A3(new_n586), .A4(new_n678), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n744), .A2(new_n278), .A3(new_n457), .A4(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(G113gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n704), .ZN(new_n922));
  INV_X1    g721(.A(new_n918), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n911), .B1(new_n704), .B2(new_n914), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n913), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n914), .A2(new_n915), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n788), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n923), .B1(new_n928), .B2(new_n585), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n794), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n465), .A2(new_n469), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(new_n278), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(new_n704), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n922), .B1(new_n933), .B2(new_n921), .ZN(G1340gat));
  OAI21_X1  g733(.A(G120gat), .B1(new_n920), .B2(new_n819), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n819), .A2(G120gat), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n935), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT118), .ZN(G1341gat));
  OAI21_X1  g738(.A(G127gat), .B1(new_n920), .B2(new_n585), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n586), .A2(new_n302), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n932), .B2(new_n941), .ZN(G1342gat));
  INV_X1    g741(.A(G134gat), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n476), .A2(new_n678), .ZN(new_n944));
  AND4_X1   g743(.A1(new_n943), .A2(new_n930), .A3(new_n931), .A4(new_n944), .ZN(new_n945));
  XOR2_X1   g744(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n946));
  OR2_X1    g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G134gat), .B1(new_n920), .B2(new_n678), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n946), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G1343gat));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n465), .B1(new_n917), .B2(new_n918), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(KEYINPUT57), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT57), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT120), .B(new_n954), .C1(new_n929), .C2(new_n465), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n465), .A2(new_n954), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n924), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n907), .A2(KEYINPUT121), .A3(new_n911), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(new_n678), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n586), .B1(new_n960), .B2(new_n927), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n956), .B1(new_n961), .B2(new_n923), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n953), .A2(new_n955), .A3(new_n962), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n794), .A2(new_n761), .A3(new_n476), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n834), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT122), .B1(new_n965), .B2(G141gat), .ZN(new_n966));
  INV_X1    g765(.A(new_n474), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n744), .A2(new_n967), .A3(new_n919), .ZN(new_n968));
  NOR4_X1   g767(.A1(new_n968), .A2(G141gat), .A3(new_n476), .A4(new_n704), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n969), .B1(new_n965), .B2(G141gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n966), .A2(new_n970), .A3(KEYINPUT58), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT58), .ZN(new_n972));
  AOI221_X4 g771(.A(new_n969), .B1(KEYINPUT122), .B2(new_n972), .C1(new_n965), .C2(G141gat), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n971), .A2(new_n973), .ZN(G1344gat));
  NOR2_X1   g773(.A1(new_n968), .A2(new_n476), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(new_n289), .A3(new_n740), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n963), .A2(new_n964), .ZN(new_n977));
  AOI211_X1 g776(.A(KEYINPUT59), .B(new_n289), .C1(new_n977), .C2(new_n740), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT59), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n926), .A2(new_n677), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n586), .B1(new_n960), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n764), .B1(new_n981), .B2(new_n923), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(new_n954), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n919), .A2(new_n956), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n740), .B(new_n964), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n979), .B1(new_n985), .B2(G148gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n976), .B1(new_n978), .B2(new_n986), .ZN(G1345gat));
  NAND3_X1  g786(.A1(new_n975), .A2(new_n283), .A3(new_n586), .ZN(new_n988));
  AND2_X1   g787(.A1(new_n977), .A2(new_n586), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n989), .B2(new_n283), .ZN(G1346gat));
  NOR4_X1   g789(.A1(new_n968), .A2(G162gat), .A3(new_n476), .A4(new_n678), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT123), .Z(new_n992));
  AND2_X1   g791(.A1(new_n977), .A2(new_n788), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n992), .B1(new_n993), .B2(new_n284), .ZN(G1347gat));
  NOR2_X1   g793(.A1(new_n744), .A2(new_n929), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n995), .A2(new_n931), .A3(new_n476), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(G169gat), .B1(new_n997), .B2(new_n834), .ZN(new_n998));
  OAI21_X1  g797(.A(KEYINPUT124), .B1(new_n744), .B2(new_n278), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n794), .A2(new_n1000), .A3(new_n476), .ZN(new_n1001));
  AND4_X1   g800(.A1(new_n457), .A2(new_n999), .A3(new_n919), .A4(new_n1001), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n704), .A2(new_n250), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n998), .B1(new_n1002), .B2(new_n1003), .ZN(G1348gat));
  AOI21_X1  g803(.A(G176gat), .B1(new_n997), .B2(new_n740), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n819), .A2(new_n249), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1005), .B1(new_n1002), .B2(new_n1006), .ZN(G1349gat));
  AOI21_X1  g806(.A(new_n222), .B1(new_n1002), .B2(new_n586), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n586), .A2(new_n228), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n996), .A2(new_n1009), .ZN(new_n1010));
  OR3_X1    g809(.A1(new_n1008), .A2(KEYINPUT60), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g810(.A(KEYINPUT60), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1350gat));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n223), .A3(new_n788), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1002), .A2(new_n677), .ZN(new_n1015));
  XNOR2_X1  g814(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1016));
  AND3_X1   g815(.A1(new_n1015), .A2(G190gat), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1016), .B1(new_n1015), .B2(G190gat), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(G1351gat));
  NOR2_X1   g818(.A1(new_n474), .A2(new_n278), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n995), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g821(.A(G197gat), .B1(new_n1022), .B2(new_n834), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n983), .A2(new_n984), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n999), .A2(new_n760), .A3(new_n1001), .ZN(new_n1025));
  AND2_X1   g824(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g825(.A1(new_n834), .A2(G197gat), .ZN(new_n1027));
  AOI21_X1  g826(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(G1352gat));
  NAND3_X1  g827(.A1(new_n1024), .A2(new_n740), .A3(new_n1025), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1029), .A2(G204gat), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n1021), .A2(G204gat), .A3(new_n819), .ZN(new_n1031));
  XNOR2_X1  g830(.A(new_n1031), .B(KEYINPUT62), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1030), .A2(new_n1032), .ZN(G1353gat));
  NAND3_X1  g832(.A1(new_n1022), .A2(new_n203), .A3(new_n586), .ZN(new_n1034));
  OAI211_X1 g833(.A(new_n1025), .B(new_n586), .C1(new_n983), .C2(new_n984), .ZN(new_n1035));
  AND3_X1   g834(.A1(new_n1035), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1036));
  AOI21_X1  g835(.A(KEYINPUT63), .B1(new_n1035), .B2(G211gat), .ZN(new_n1037));
  OAI21_X1  g836(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(G1354gat));
  OAI21_X1  g837(.A(new_n204), .B1(new_n1021), .B2(new_n913), .ZN(new_n1039));
  XNOR2_X1  g838(.A(new_n1039), .B(KEYINPUT126), .ZN(new_n1040));
  NOR2_X1   g839(.A1(new_n678), .A2(new_n204), .ZN(new_n1041));
  AOI21_X1  g840(.A(new_n1040), .B1(new_n1026), .B2(new_n1041), .ZN(G1355gat));
endmodule


