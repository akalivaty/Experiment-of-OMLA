//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT84), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT0), .A4(G128), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n191), .A2(new_n193), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT0), .B(G128), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT72), .B(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(new_n193), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT65), .B(KEYINPUT1), .C1(new_n192), .C2(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(G128), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n204), .B1(new_n209), .B2(new_n201), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n200), .B1(new_n210), .B2(new_n199), .ZN(new_n211));
  INV_X1    g025(.A(G224), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G953), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n211), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G104), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(G101), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n222), .A2(KEYINPUT78), .A3(G101), .A4(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(G116), .B(G119), .Z(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n229), .A2(KEYINPUT66), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT2), .B(G113), .Z(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n231), .A2(new_n235), .B1(new_n234), .B2(new_n233), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT75), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n222), .B2(G101), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G101), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n217), .A2(new_n220), .A3(new_n241), .A4(new_n221), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n222), .A2(new_n238), .A3(G101), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n243), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT76), .B1(new_n247), .B2(new_n239), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n237), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT5), .ZN(new_n250));
  INV_X1    g064(.A(G119), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(G116), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT80), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(G113), .C1(new_n250), .C2(new_n229), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT66), .B1(new_n229), .B2(new_n230), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n233), .A2(new_n232), .A3(new_n234), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n216), .A2(G107), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n219), .A2(G104), .ZN(new_n259));
  OAI21_X1  g073(.A(G101), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n242), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n254), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n215), .B1(new_n249), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n248), .A2(new_n246), .ZN(new_n265));
  OAI211_X1 g079(.A(KEYINPUT81), .B(new_n262), .C1(new_n265), .C2(new_n237), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G122), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n249), .A2(new_n263), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(new_n267), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n267), .A2(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n264), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT82), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n264), .A2(new_n266), .A3(new_n276), .A4(new_n273), .ZN(new_n277));
  AOI221_X4 g091(.A(new_n214), .B1(new_n269), .B2(new_n272), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n261), .B1(new_n254), .B2(new_n257), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n263), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n267), .B(KEYINPUT8), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT7), .B1(new_n212), .B2(G953), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n211), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n211), .A2(new_n282), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n280), .A2(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n285), .A2(KEYINPUT83), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n285), .A2(KEYINPUT83), .B1(new_n271), .B2(new_n267), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n189), .B1(new_n278), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT9), .B(G234), .ZN(new_n292));
  OAI21_X1  g106(.A(G221), .B1(new_n292), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n289), .ZN(new_n296));
  INV_X1    g110(.A(G953), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G227), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(KEYINPUT74), .ZN(new_n299));
  XNOR2_X1  g113(.A(G110), .B(G140), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n228), .A2(new_n198), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(new_n246), .B2(new_n248), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n195), .B1(G128), .B2(new_n205), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n261), .B1(new_n304), .B2(new_n204), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT10), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n242), .A2(new_n260), .A3(KEYINPUT10), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n210), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n208), .A2(G128), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT65), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n201), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n204), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n309), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT79), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n307), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT11), .B1(new_n319), .B2(G137), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT11), .ZN(new_n321));
  INV_X1    g135(.A(G137), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G134), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT64), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n322), .B2(G134), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n319), .A2(KEYINPUT64), .A3(G137), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n324), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n327), .A2(new_n328), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n325), .B1(new_n331), .B2(new_n324), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n303), .A2(new_n318), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n248), .A2(new_n246), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n197), .B1(new_n226), .B2(new_n227), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n308), .B1(new_n210), .B2(new_n309), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT79), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n339), .A2(new_n340), .B1(new_n306), .B2(new_n305), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n333), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n301), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n338), .A2(new_n333), .A3(new_n341), .ZN(new_n344));
  INV_X1    g158(.A(new_n301), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n305), .B1(new_n315), .B2(new_n261), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n334), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT12), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT12), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n349), .A3(new_n334), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n344), .A2(new_n345), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(G902), .B1(new_n343), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n296), .B1(new_n352), .B2(new_n295), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n344), .A2(new_n348), .A3(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n301), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n334), .B1(new_n303), .B2(new_n318), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n344), .A3(new_n345), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(G469), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n294), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G214), .B1(G237), .B2(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n275), .A2(new_n277), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n269), .A2(new_n272), .ZN(new_n362));
  INV_X1    g176(.A(new_n214), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n286), .B2(new_n287), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n188), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n291), .A2(new_n359), .A3(new_n360), .A4(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G475), .ZN(new_n368));
  INV_X1    g182(.A(G237), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n297), .A3(G214), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(G143), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT18), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(new_n325), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n370), .B(new_n192), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT18), .A3(G131), .ZN(new_n375));
  NOR2_X1   g189(.A1(G125), .A2(G140), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n199), .B2(G140), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(G146), .ZN(new_n378));
  XOR2_X1   g192(.A(G125), .B(G140), .Z(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G146), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n373), .B(new_n375), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n374), .A2(G131), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n325), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(KEYINPUT17), .A3(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT16), .ZN(new_n388));
  AND2_X1   g202(.A1(KEYINPUT72), .A2(G125), .ZN(new_n389));
  NOR2_X1   g203(.A1(KEYINPUT72), .A2(G125), .ZN(new_n390));
  OAI21_X1  g204(.A(G140), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n376), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(KEYINPUT16), .A2(G140), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n199), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n190), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n199), .A2(new_n394), .ZN(new_n397));
  OAI211_X1 g211(.A(G146), .B(new_n397), .C1(new_n377), .C2(new_n388), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n381), .B1(new_n387), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n216), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n402), .B(new_n381), .C1(new_n387), .C2(new_n399), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n368), .B1(new_n406), .B2(new_n289), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  INV_X1    g222(.A(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n382), .A2(new_n383), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n379), .A2(KEYINPUT19), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(KEYINPUT19), .B2(new_n377), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n398), .B(new_n410), .C1(new_n413), .C2(G146), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n402), .B1(new_n414), .B2(new_n381), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n408), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n381), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n403), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n416), .B1(new_n420), .B2(KEYINPUT20), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n419), .A2(new_n405), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n417), .A3(new_n423), .A4(new_n408), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n407), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(KEYINPUT87), .A2(G952), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT87), .A2(G952), .ZN(new_n428));
  AOI21_X1  g242(.A(G953), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G234), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(new_n369), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(G902), .B(G953), .C1(new_n430), .C2(new_n369), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT88), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(G898), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n292), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(G217), .A3(new_n297), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n192), .A2(G128), .ZN(new_n441));
  INV_X1    g255(.A(G128), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G143), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(new_n319), .ZN(new_n445));
  XNOR2_X1  g259(.A(G116), .B(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n219), .ZN(new_n447));
  INV_X1    g261(.A(G116), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT14), .A3(G122), .ZN(new_n449));
  INV_X1    g263(.A(new_n446), .ZN(new_n450));
  OAI211_X1 g264(.A(G107), .B(new_n449), .C1(new_n450), .C2(KEYINPUT14), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n453));
  INV_X1    g267(.A(new_n441), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n443), .B1(new_n454), .B2(KEYINPUT13), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT13), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n441), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G134), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n446), .B(new_n219), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n444), .A2(new_n319), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n452), .A2(new_n453), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n453), .B1(new_n452), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n440), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  INV_X1    g280(.A(new_n440), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n467), .A3(new_n462), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n468), .A3(new_n289), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n469), .B(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n425), .A2(new_n438), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n367), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT22), .B(G137), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n297), .A2(G221), .A3(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n442), .A2(G119), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n251), .A2(G128), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT24), .B(G110), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n251), .B2(G128), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n442), .A2(KEYINPUT23), .A3(G119), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n485), .A2(new_n486), .A3(new_n480), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT71), .ZN(new_n488));
  INV_X1    g302(.A(G110), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n486), .A3(new_n480), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT71), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n483), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n489), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n481), .A2(new_n482), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n380), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n399), .A2(new_n493), .B1(new_n398), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n478), .B1(new_n497), .B2(KEYINPUT73), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n399), .A2(new_n493), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n398), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT73), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n502), .A3(new_n478), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT25), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G217), .B1(new_n430), .B2(G902), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT70), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n506), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n504), .A2(new_n505), .ZN(new_n512));
  INV_X1    g326(.A(new_n510), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(G902), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n508), .A2(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n319), .A2(G137), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n322), .A2(G134), .ZN(new_n520));
  OAI21_X1  g334(.A(G131), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n329), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n518), .B1(new_n210), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n315), .A2(KEYINPUT67), .A3(new_n329), .A4(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n198), .B1(new_n330), .B2(new_n332), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n255), .A2(new_n256), .B1(new_n229), .B2(new_n230), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n369), .A2(new_n297), .A3(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT27), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT30), .A4(new_n525), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n210), .A2(new_n522), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n324), .A2(new_n327), .A3(new_n328), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G131), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n197), .B1(new_n539), .B2(new_n329), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n536), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  AND4_X1   g355(.A1(new_n534), .A2(new_n535), .A3(new_n236), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n202), .B1(G143), .B2(new_n190), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n442), .B1(new_n543), .B2(KEYINPUT65), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n195), .B1(new_n544), .B2(new_n207), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n329), .B(new_n521), .C1(new_n545), .C2(new_n204), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n525), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n526), .B1(new_n547), .B2(new_n536), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n534), .B1(new_n548), .B2(new_n535), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n517), .B(new_n533), .C1(new_n542), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n547), .B2(new_n236), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n547), .A2(new_n236), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n552), .B(new_n553), .C1(new_n551), .C2(new_n527), .ZN(new_n554));
  INV_X1    g368(.A(new_n531), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n535), .A2(new_n236), .A3(new_n541), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT68), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n548), .A2(new_n534), .A3(new_n535), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n532), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n561), .A2(KEYINPUT69), .A3(new_n517), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n533), .B1(new_n542), .B2(new_n549), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(KEYINPUT31), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n557), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n552), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n236), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n527), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n571), .B1(new_n574), .B2(KEYINPUT28), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n555), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n559), .A2(new_n560), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n531), .B1(new_n579), .B2(new_n527), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n576), .B1(new_n554), .B2(new_n555), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n566), .A2(new_n570), .B1(G472), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n550), .A2(new_n556), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT69), .B1(new_n561), .B2(new_n517), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n564), .A2(new_n563), .A3(KEYINPUT31), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n569), .B1(new_n587), .B2(new_n568), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n516), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n475), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  OAI21_X1  g405(.A(KEYINPUT89), .B1(new_n587), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT89), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n566), .A2(new_n593), .A3(new_n289), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n594), .A3(G472), .ZN(new_n595));
  AND4_X1   g409(.A1(new_n344), .A2(new_n345), .A3(new_n348), .A4(new_n350), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n345), .B1(new_n356), .B2(new_n344), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n295), .B(new_n289), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n296), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n358), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n515), .A2(new_n600), .A3(new_n293), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n587), .A2(new_n568), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n595), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n604), .B1(new_n595), .B2(new_n603), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT91), .B(KEYINPUT33), .Z(new_n609));
  AND3_X1   g423(.A1(new_n465), .A2(new_n468), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n465), .A2(new_n468), .B1(KEYINPUT91), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n470), .A2(G902), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n613), .A2(new_n614), .B1(new_n470), .B2(new_n469), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n425), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n291), .A2(new_n438), .A3(new_n360), .A4(new_n366), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n608), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  XNOR2_X1  g435(.A(new_n416), .B(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n406), .A2(new_n289), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G475), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT92), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n407), .A2(KEYINPUT92), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n622), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n628), .A2(new_n473), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n608), .A2(new_n618), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  INV_X1    g447(.A(new_n367), .ZN(new_n634));
  INV_X1    g448(.A(new_n602), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n478), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n501), .B(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n514), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n506), .A2(new_n507), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n513), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n506), .A2(new_n507), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n645), .A2(new_n425), .A3(new_n438), .A4(new_n473), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n634), .A2(new_n635), .A3(new_n595), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT93), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  NAND3_X1  g465(.A1(new_n645), .A2(new_n600), .A3(new_n293), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n583), .B2(new_n588), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n364), .A2(new_n365), .A3(new_n188), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n188), .B1(new_n364), .B2(new_n365), .ZN(new_n655));
  INV_X1    g469(.A(new_n360), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n431), .B(KEYINPUT94), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n659), .B1(new_n660), .B2(new_n435), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n629), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n653), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NOR2_X1   g478(.A1(new_n654), .A2(new_n655), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT38), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n291), .A2(new_n366), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT38), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n661), .B(KEYINPUT39), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n359), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT40), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n527), .B1(new_n542), .B2(new_n549), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n531), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n574), .A2(new_n531), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(G902), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n566), .A2(new_n570), .B1(G472), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n588), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n425), .A2(new_n473), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n640), .B1(new_n508), .B2(new_n511), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n360), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT95), .ZN(new_n685));
  OR4_X1    g499(.A1(new_n670), .A2(new_n673), .A3(new_n681), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT96), .B(G143), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G45));
  NOR3_X1   g502(.A1(new_n615), .A2(new_n425), .A3(new_n661), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n653), .A2(new_n657), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  OAI21_X1  g505(.A(new_n289), .B1(new_n596), .B2(new_n597), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n693), .A2(new_n293), .A3(new_n598), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n618), .A2(new_n589), .A3(new_n616), .A4(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT41), .B(G113), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT97), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n695), .B(new_n697), .ZN(G15));
  NAND4_X1  g512(.A1(new_n618), .A2(new_n589), .A3(new_n630), .A4(new_n694), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  AND4_X1   g514(.A1(new_n360), .A2(new_n291), .A3(new_n366), .A4(new_n694), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n646), .B1(new_n583), .B2(new_n588), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  INV_X1    g518(.A(KEYINPUT99), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n694), .A2(new_n438), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n657), .A2(new_n707), .A3(new_n682), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n587), .B2(G902), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n567), .B(KEYINPUT98), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n550), .B1(new_n531), .B2(new_n575), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n561), .A2(new_n517), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n709), .A2(new_n515), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n705), .B1(new_n708), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n291), .A2(new_n682), .A3(new_n360), .A4(new_n366), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n706), .ZN(new_n717));
  INV_X1    g531(.A(new_n714), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(KEYINPUT99), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  AND4_X1   g535(.A1(new_n645), .A2(new_n709), .A3(new_n689), .A4(new_n713), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n701), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(KEYINPUT101), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT32), .B1(new_n566), .B2(new_n567), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n581), .B1(new_n555), .B2(new_n674), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n575), .A2(new_n577), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n289), .ZN(new_n732));
  OAI21_X1  g546(.A(G472), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n570), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n733), .B1(new_n587), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n515), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n355), .A2(KEYINPUT100), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT100), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n354), .A2(new_n738), .A3(new_n301), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(G469), .A3(new_n357), .A4(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n294), .B1(new_n353), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n360), .B(new_n741), .C1(new_n654), .C2(new_n655), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n725), .A2(new_n726), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n689), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n728), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n736), .A2(new_n742), .A3(new_n745), .A4(new_n727), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  NAND2_X1  g564(.A1(new_n743), .A2(new_n662), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  AOI21_X1  g566(.A(KEYINPUT45), .B1(new_n355), .B2(new_n357), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n295), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n737), .A2(KEYINPUT45), .A3(new_n357), .A4(new_n739), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n296), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n756), .A2(KEYINPUT103), .A3(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT103), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n598), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n293), .A3(new_n671), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n613), .A2(new_n614), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n469), .A2(new_n470), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT105), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n765), .B(new_n425), .C1(new_n766), .C2(KEYINPUT43), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n421), .A2(new_n424), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n624), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n771));
  OAI22_X1  g585(.A1(new_n769), .A2(new_n615), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n767), .A2(new_n772), .A3(KEYINPUT106), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n683), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n595), .A2(new_n635), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT44), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n656), .B1(new_n291), .B2(new_n366), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n777), .A2(KEYINPUT44), .A3(new_n778), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n762), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(KEYINPUT107), .B(G137), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G39));
  NAND2_X1  g601(.A1(new_n760), .A2(new_n293), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n760), .A2(KEYINPUT47), .A3(new_n293), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n588), .A2(new_n583), .A3(new_n516), .A4(new_n689), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n780), .A3(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT108), .B(G140), .Z(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G42));
  NAND2_X1  g610(.A1(new_n693), .A2(new_n598), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(KEYINPUT49), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n294), .A2(new_n656), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n515), .A2(new_n765), .A3(new_n425), .A4(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n670), .A2(new_n681), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n661), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n473), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n628), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n780), .A2(KEYINPUT109), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n360), .B(new_n806), .C1(new_n654), .C2(new_n655), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT109), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n653), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(KEYINPUT110), .A3(new_n653), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n589), .A2(new_n741), .A3(new_n780), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n727), .B1(new_n817), .B2(new_n745), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n743), .A2(new_n746), .A3(new_n728), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n722), .A2(new_n741), .A3(new_n780), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n751), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n473), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n616), .B1(new_n425), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n617), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n608), .A2(new_n824), .B1(new_n715), .B2(new_n719), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n648), .A2(new_n695), .A3(new_n699), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n590), .A2(new_n703), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n816), .A2(new_n821), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n653), .B(new_n657), .C1(new_n662), .C2(new_n689), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n640), .B(new_n661), .C1(new_n508), .C2(new_n511), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n741), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n657), .A2(new_n835), .A3(new_n680), .A4(new_n682), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n723), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n832), .B(KEYINPUT52), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT112), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n837), .B2(new_n832), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n837), .B(new_n842), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n595), .A2(new_n603), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT90), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n605), .A3(new_n824), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT99), .B1(new_n717), .B2(new_n718), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n716), .A2(new_n714), .A3(new_n705), .A4(new_n706), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n475), .A2(new_n589), .B1(new_n701), .B2(new_n702), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n648), .A3(new_n695), .A4(new_n699), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n846), .A2(new_n855), .A3(new_n816), .A4(new_n821), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n830), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n845), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n694), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n781), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n658), .B1(new_n767), .B2(new_n772), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n589), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT48), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n718), .A2(new_n862), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n701), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n680), .A2(new_n516), .A3(new_n431), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n616), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n864), .A2(new_n429), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n866), .A2(KEYINPUT114), .A3(new_n780), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n865), .B2(new_n781), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n797), .A2(new_n293), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n792), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n709), .A2(new_n713), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n645), .A2(new_n861), .A3(new_n878), .A4(new_n862), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n765), .A2(new_n769), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n861), .A2(new_n868), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(KEYINPUT117), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(KEYINPUT117), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n860), .A2(new_n360), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n666), .A2(new_n669), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n666), .A2(new_n669), .A3(KEYINPUT115), .A4(new_n885), .ZN(new_n889));
  OR2_X1    g703(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n888), .A2(new_n866), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n888), .A2(new_n866), .A3(new_n889), .ZN(new_n892));
  XOR2_X1   g706(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n877), .A2(new_n884), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT51), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT51), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n877), .A2(new_n884), .A3(new_n897), .A4(new_n894), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n871), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n837), .B(KEYINPUT52), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n829), .A2(new_n830), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n751), .A2(new_n820), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT110), .B1(new_n811), .B2(new_n653), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n359), .B(new_n645), .C1(new_n729), .C2(new_n735), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n813), .B(new_n904), .C1(new_n807), .C2(new_n810), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n749), .B(new_n902), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n648), .A2(new_n695), .A3(new_n699), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(new_n720), .A3(new_n853), .A4(new_n849), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT111), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT111), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n855), .A2(new_n910), .A3(new_n816), .A4(new_n821), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n844), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n901), .B1(new_n912), .B2(new_n830), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n859), .B(new_n899), .C1(new_n913), .C2(new_n858), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT119), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n914), .B2(new_n915), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n803), .B1(new_n916), .B2(new_n919), .ZN(G75));
  NAND2_X1  g734(.A1(new_n845), .A2(new_n857), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(G902), .A3(new_n188), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n361), .A2(new_n362), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n363), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n297), .A2(G952), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G51));
  XNOR2_X1  g744(.A(new_n296), .B(KEYINPUT57), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n831), .A2(new_n844), .B1(new_n830), .B2(new_n856), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n858), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n845), .A2(new_n858), .A3(new_n857), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n343), .A2(new_n351), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n921), .A2(G902), .A3(new_n755), .A4(new_n754), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n929), .B1(new_n937), .B2(new_n938), .ZN(G54));
  NAND4_X1  g753(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n940));
  INV_X1    g754(.A(new_n422), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n929), .ZN(G60));
  XOR2_X1   g758(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n945));
  NOR2_X1   g759(.A1(new_n470), .A2(new_n289), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n613), .B(new_n948), .C1(new_n933), .C2(new_n934), .ZN(new_n949));
  INV_X1    g763(.A(new_n929), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n859), .B1(new_n913), .B2(new_n858), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n613), .B1(new_n952), .B2(new_n948), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(G63));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(KEYINPUT61), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n950), .B1(new_n955), .B2(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n932), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n638), .B(KEYINPUT121), .Z(new_n961));
  AOI21_X1  g775(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n505), .B(new_n504), .C1(new_n932), .C2(new_n959), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n956), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n959), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n921), .A2(new_n965), .A3(new_n961), .ZN(new_n966));
  INV_X1    g780(.A(new_n957), .ZN(new_n967));
  AND4_X1   g781(.A1(new_n956), .A2(new_n963), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n964), .A2(new_n968), .ZN(G66));
  OAI21_X1  g783(.A(G953), .B1(new_n436), .B2(new_n212), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n855), .B2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n924), .B1(G898), .B2(new_n297), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  INV_X1    g787(.A(KEYINPUT62), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n833), .A2(new_n723), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n686), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT124), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n686), .A2(new_n974), .A3(new_n975), .ZN(new_n978));
  NOR4_X1   g792(.A1(new_n781), .A2(new_n736), .A3(new_n823), .A4(new_n672), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT125), .Z(new_n980));
  NAND4_X1  g794(.A1(new_n785), .A2(new_n978), .A3(new_n794), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n297), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n535), .A2(new_n541), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT123), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(new_n413), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n736), .A2(new_n716), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n762), .A2(new_n783), .A3(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n749), .A2(new_n751), .A3(new_n975), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n785), .A2(new_n988), .A3(new_n794), .A4(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(G953), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n985), .B1(G900), .B2(G953), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n297), .B1(G227), .B2(G900), .ZN(new_n994));
  AOI22_X1  g808(.A1(new_n991), .A2(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n986), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n994), .A2(new_n993), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n990), .B2(new_n908), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n674), .A2(new_n531), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n929), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n675), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n977), .A2(new_n908), .A3(new_n981), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1000), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OR3_X1    g823(.A1(new_n1006), .A2(new_n1002), .A3(new_n1008), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n913), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1005), .A2(new_n1011), .ZN(G57));
endmodule


