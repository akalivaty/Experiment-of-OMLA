

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U551 ( .A1(G2105), .A2(n559), .ZN(n890) );
  XOR2_X1 U552 ( .A(KEYINPUT23), .B(n570), .Z(n518) );
  OR2_X1 U553 ( .A1(n784), .A2(n783), .ZN(n519) );
  XOR2_X1 U554 ( .A(KEYINPUT87), .B(n771), .Z(n520) );
  BUF_X1 U555 ( .A(n699), .Z(n740) );
  OR2_X1 U556 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U557 ( .A1(n760), .A2(G1966), .ZN(n748) );
  AND2_X1 U558 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U559 ( .A1(n689), .A2(n769), .ZN(n699) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n556) );
  NOR2_X1 U561 ( .A1(G651), .A2(n626), .ZN(n652) );
  OR2_X1 U562 ( .A1(n573), .A2(n572), .ZN(n574) );
  INV_X1 U563 ( .A(G651), .ZN(n526) );
  NOR2_X1 U564 ( .A1(G543), .A2(n526), .ZN(n522) );
  XNOR2_X1 U565 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n521) );
  XNOR2_X1 U566 ( .A(n522), .B(n521), .ZN(n645) );
  NAND2_X1 U567 ( .A1(G63), .A2(n645), .ZN(n524) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n626) );
  NAND2_X1 U569 ( .A1(G51), .A2(n652), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U571 ( .A(KEYINPUT6), .B(n525), .ZN(n533) );
  NOR2_X1 U572 ( .A1(n626), .A2(n526), .ZN(n648) );
  NAND2_X1 U573 ( .A1(n648), .A2(G76), .ZN(n527) );
  XNOR2_X1 U574 ( .A(KEYINPUT76), .B(n527), .ZN(n530) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U576 ( .A1(n644), .A2(G89), .ZN(n528) );
  XNOR2_X1 U577 ( .A(KEYINPUT4), .B(n528), .ZN(n529) );
  NAND2_X1 U578 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U579 ( .A(n531), .B(KEYINPUT5), .Z(n532) );
  NOR2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U581 ( .A(KEYINPUT77), .B(n534), .Z(n535) );
  XOR2_X1 U582 ( .A(KEYINPUT7), .B(n535), .Z(G168) );
  XOR2_X1 U583 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U584 ( .A(KEYINPUT109), .B(G2446), .Z(n537) );
  XNOR2_X1 U585 ( .A(G2430), .B(G2451), .ZN(n536) );
  XNOR2_X1 U586 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U587 ( .A(n538), .B(KEYINPUT110), .Z(n540) );
  XNOR2_X1 U588 ( .A(G1348), .B(G1341), .ZN(n539) );
  XNOR2_X1 U589 ( .A(n540), .B(n539), .ZN(n544) );
  XOR2_X1 U590 ( .A(G2435), .B(KEYINPUT111), .Z(n542) );
  XNOR2_X1 U591 ( .A(G2438), .B(G2454), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U593 ( .A(n544), .B(n543), .Z(n546) );
  XNOR2_X1 U594 ( .A(G2443), .B(G2427), .ZN(n545) );
  XNOR2_X1 U595 ( .A(n546), .B(n545), .ZN(n547) );
  AND2_X1 U596 ( .A1(n547), .A2(G14), .ZN(G401) );
  NAND2_X1 U597 ( .A1(G64), .A2(n645), .ZN(n549) );
  NAND2_X1 U598 ( .A1(G52), .A2(n652), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U600 ( .A1(G77), .A2(n648), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G90), .A2(n644), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n552), .Z(n553) );
  XNOR2_X1 U604 ( .A(KEYINPUT9), .B(n553), .ZN(n554) );
  NOR2_X1 U605 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X2 U607 ( .A(KEYINPUT17), .B(n556), .Z(n892) );
  NAND2_X1 U608 ( .A1(G135), .A2(n892), .ZN(n557) );
  XNOR2_X1 U609 ( .A(n557), .B(KEYINPUT78), .ZN(n566) );
  INV_X1 U610 ( .A(G2104), .ZN(n559) );
  AND2_X1 U611 ( .A1(n559), .A2(G2105), .ZN(n886) );
  NAND2_X1 U612 ( .A1(n886), .A2(G123), .ZN(n558) );
  XNOR2_X1 U613 ( .A(n558), .B(KEYINPUT18), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G99), .A2(n890), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n564) );
  AND2_X1 U616 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U617 ( .A1(G111), .A2(n887), .ZN(n562) );
  XNOR2_X1 U618 ( .A(KEYINPUT79), .B(n562), .ZN(n563) );
  NOR2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n566), .A2(n565), .ZN(n1002) );
  XNOR2_X1 U621 ( .A(G2096), .B(n1002), .ZN(n567) );
  OR2_X1 U622 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U623 ( .A(G57), .ZN(G237) );
  NAND2_X1 U624 ( .A1(G125), .A2(n886), .ZN(n569) );
  NAND2_X1 U625 ( .A1(G137), .A2(n892), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G101), .A2(n890), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G113), .A2(n887), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n518), .A2(n571), .ZN(n572) );
  XNOR2_X1 U630 ( .A(n574), .B(KEYINPUT65), .ZN(G160) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U632 ( .A(n575), .B(KEYINPUT70), .ZN(n576) );
  XNOR2_X1 U633 ( .A(KEYINPUT10), .B(n576), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n835) );
  NAND2_X1 U635 ( .A1(n835), .A2(G567), .ZN(n577) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  NAND2_X1 U637 ( .A1(n644), .A2(G81), .ZN(n578) );
  XNOR2_X1 U638 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G68), .A2(n648), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n582) );
  XOR2_X1 U641 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n581) );
  XNOR2_X1 U642 ( .A(n582), .B(n581), .ZN(n586) );
  NAND2_X1 U643 ( .A1(G56), .A2(n645), .ZN(n583) );
  XNOR2_X1 U644 ( .A(n583), .B(KEYINPUT71), .ZN(n584) );
  XNOR2_X1 U645 ( .A(KEYINPUT14), .B(n584), .ZN(n585) );
  NOR2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n652), .A2(G43), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n588), .A2(n587), .ZN(n918) );
  INV_X1 U649 ( .A(G860), .ZN(n609) );
  OR2_X1 U650 ( .A1(n918), .A2(n609), .ZN(G153) );
  XNOR2_X1 U651 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(KEYINPUT74), .ZN(n599) );
  NAND2_X1 U654 ( .A1(G54), .A2(n652), .ZN(n596) );
  NAND2_X1 U655 ( .A1(G79), .A2(n648), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G92), .A2(n644), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G66), .A2(n645), .ZN(n592) );
  XNOR2_X1 U659 ( .A(KEYINPUT75), .B(n592), .ZN(n593) );
  NOR2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n597), .B(KEYINPUT15), .ZN(n923) );
  OR2_X1 U663 ( .A1(G868), .A2(n923), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U665 ( .A1(G78), .A2(n648), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G91), .A2(n644), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U668 ( .A1(G65), .A2(n645), .ZN(n602) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n602), .ZN(n603) );
  NOR2_X1 U670 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U671 ( .A1(n652), .A2(G53), .ZN(n605) );
  NAND2_X1 U672 ( .A1(n606), .A2(n605), .ZN(G299) );
  INV_X1 U673 ( .A(G868), .ZN(n664) );
  NOR2_X1 U674 ( .A1(G286), .A2(n664), .ZN(n608) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n610), .A2(n923), .ZN(n611) );
  XNOR2_X1 U679 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n918), .ZN(n614) );
  NAND2_X1 U681 ( .A1(G868), .A2(n923), .ZN(n612) );
  NOR2_X1 U682 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U683 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G559), .A2(n923), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n918), .B(n615), .ZN(n661) );
  NOR2_X1 U686 ( .A1(n661), .A2(G860), .ZN(n622) );
  NAND2_X1 U687 ( .A1(G67), .A2(n645), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G55), .A2(n652), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G80), .A2(n648), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G93), .A2(n644), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n663) );
  XNOR2_X1 U694 ( .A(n622), .B(n663), .ZN(G145) );
  NAND2_X1 U695 ( .A1(G49), .A2(n652), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G74), .A2(G651), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U698 ( .A1(n645), .A2(n625), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n626), .A2(G87), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U701 ( .A1(G73), .A2(n648), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n629), .B(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U703 ( .A1(G61), .A2(n645), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G48), .A2(n652), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n644), .A2(G86), .ZN(n632) );
  XOR2_X1 U707 ( .A(KEYINPUT80), .B(n632), .Z(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G62), .A2(n645), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G50), .A2(n652), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U713 ( .A1(G75), .A2(n648), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G88), .A2(n644), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(KEYINPUT81), .ZN(G303) );
  NAND2_X1 U718 ( .A1(G85), .A2(n644), .ZN(n647) );
  NAND2_X1 U719 ( .A1(G60), .A2(n645), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U721 ( .A1(G72), .A2(n648), .ZN(n649) );
  XOR2_X1 U722 ( .A(KEYINPUT66), .B(n649), .Z(n650) );
  NOR2_X1 U723 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n652), .A2(G47), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n654), .A2(n653), .ZN(G290) );
  XOR2_X1 U726 ( .A(KEYINPUT19), .B(KEYINPUT82), .Z(n655) );
  XNOR2_X1 U727 ( .A(G288), .B(n655), .ZN(n658) );
  INV_X1 U728 ( .A(G299), .ZN(n715) );
  XNOR2_X1 U729 ( .A(n715), .B(G305), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(G303), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n660) );
  XNOR2_X1 U732 ( .A(G290), .B(n663), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(n907) );
  XOR2_X1 U734 ( .A(n661), .B(n907), .Z(n662) );
  NAND2_X1 U735 ( .A1(n662), .A2(G868), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U738 ( .A(KEYINPUT83), .B(n667), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U745 ( .A1(G132), .A2(G82), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n672), .B(KEYINPUT84), .ZN(n673) );
  XNOR2_X1 U747 ( .A(n673), .B(KEYINPUT22), .ZN(n674) );
  NOR2_X1 U748 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U749 ( .A1(G96), .A2(n675), .ZN(n841) );
  NAND2_X1 U750 ( .A1(n841), .A2(G2106), .ZN(n679) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U752 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U753 ( .A1(G108), .A2(n677), .ZN(n842) );
  NAND2_X1 U754 ( .A1(n842), .A2(G567), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n679), .A2(n678), .ZN(n843) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U757 ( .A1(n843), .A2(n680), .ZN(n840) );
  NAND2_X1 U758 ( .A1(n840), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(n892), .A2(G138), .ZN(n683) );
  NAND2_X1 U760 ( .A1(G114), .A2(n887), .ZN(n681) );
  XOR2_X1 U761 ( .A(KEYINPUT85), .B(n681), .Z(n682) );
  NAND2_X1 U762 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U763 ( .A1(G126), .A2(n886), .ZN(n685) );
  NAND2_X1 U764 ( .A1(G102), .A2(n890), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U766 ( .A1(n687), .A2(n686), .ZN(G164) );
  INV_X1 U767 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U768 ( .A(G1981), .B(G305), .ZN(n935) );
  INV_X1 U769 ( .A(KEYINPUT92), .ZN(n691) );
  NAND2_X1 U770 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U771 ( .A(n770), .ZN(n689) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n688) );
  XNOR2_X1 U773 ( .A(KEYINPUT64), .B(n688), .ZN(n769) );
  NAND2_X1 U774 ( .A1(n699), .A2(G8), .ZN(n690) );
  XNOR2_X1 U775 ( .A(n691), .B(n690), .ZN(n781) );
  INV_X1 U776 ( .A(n781), .ZN(n760) );
  NOR2_X1 U777 ( .A1(n699), .A2(G2084), .ZN(n693) );
  INV_X1 U778 ( .A(KEYINPUT93), .ZN(n692) );
  XNOR2_X1 U779 ( .A(n693), .B(n692), .ZN(n752) );
  INV_X1 U780 ( .A(n752), .ZN(n694) );
  NAND2_X1 U781 ( .A1(G8), .A2(n694), .ZN(n695) );
  NOR2_X1 U782 ( .A1(n748), .A2(n695), .ZN(n696) );
  XOR2_X1 U783 ( .A(KEYINPUT30), .B(n696), .Z(n697) );
  NOR2_X1 U784 ( .A1(G168), .A2(n697), .ZN(n698) );
  XOR2_X1 U785 ( .A(KEYINPUT103), .B(n698), .Z(n706) );
  INV_X1 U786 ( .A(n740), .ZN(n722) );
  XNOR2_X1 U787 ( .A(G2078), .B(KEYINPUT25), .ZN(n700) );
  XNOR2_X1 U788 ( .A(n700), .B(KEYINPUT96), .ZN(n968) );
  NAND2_X1 U789 ( .A1(n722), .A2(n968), .ZN(n701) );
  XNOR2_X1 U790 ( .A(n701), .B(KEYINPUT97), .ZN(n703) );
  XOR2_X1 U791 ( .A(KEYINPUT95), .B(G1961), .Z(n949) );
  NOR2_X1 U792 ( .A1(n722), .A2(n949), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U794 ( .A(KEYINPUT98), .B(n704), .Z(n735) );
  NOR2_X1 U795 ( .A1(G171), .A2(n735), .ZN(n705) );
  XNOR2_X1 U796 ( .A(n707), .B(KEYINPUT31), .ZN(n739) );
  NAND2_X1 U797 ( .A1(n740), .A2(G1956), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n722), .A2(G2072), .ZN(n708) );
  XOR2_X1 U799 ( .A(KEYINPUT27), .B(n708), .Z(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U801 ( .A(n711), .B(KEYINPUT99), .ZN(n716) );
  NOR2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n714) );
  XNOR2_X1 U803 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n712) );
  XNOR2_X1 U804 ( .A(n712), .B(KEYINPUT28), .ZN(n713) );
  XNOR2_X1 U805 ( .A(n714), .B(n713), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n731) );
  INV_X1 U807 ( .A(G1996), .ZN(n974) );
  NOR2_X1 U808 ( .A1(n740), .A2(n974), .ZN(n717) );
  XOR2_X1 U809 ( .A(n717), .B(KEYINPUT26), .Z(n719) );
  NAND2_X1 U810 ( .A1(n740), .A2(G1341), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U812 ( .A1(n918), .A2(n720), .ZN(n721) );
  OR2_X1 U813 ( .A1(n923), .A2(n721), .ZN(n729) );
  NAND2_X1 U814 ( .A1(n923), .A2(n721), .ZN(n727) );
  AND2_X1 U815 ( .A1(n722), .A2(G2067), .ZN(n723) );
  XOR2_X1 U816 ( .A(n723), .B(KEYINPUT102), .Z(n725) );
  NAND2_X1 U817 ( .A1(n740), .A2(G1348), .ZN(n724) );
  NAND2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U823 ( .A(KEYINPUT29), .B(n734), .Z(n737) );
  NAND2_X1 U824 ( .A1(G171), .A2(n735), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n749) );
  NAND2_X1 U827 ( .A1(n749), .A2(G286), .ZN(n745) );
  NOR2_X1 U828 ( .A1(n760), .A2(G1971), .ZN(n742) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n743), .A2(G303), .ZN(n744) );
  NAND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U833 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U834 ( .A(n747), .B(KEYINPUT32), .ZN(n757) );
  INV_X1 U835 ( .A(n748), .ZN(n750) );
  XNOR2_X1 U836 ( .A(n751), .B(KEYINPUT104), .ZN(n755) );
  NAND2_X1 U837 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U838 ( .A(KEYINPUT94), .B(n753), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U840 ( .A1(n757), .A2(n756), .ZN(n780) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U843 ( .A1(n766), .A2(n758), .ZN(n927) );
  NAND2_X1 U844 ( .A1(n780), .A2(n927), .ZN(n763) );
  NAND2_X1 U845 ( .A1(G288), .A2(G1976), .ZN(n759) );
  XOR2_X1 U846 ( .A(KEYINPUT105), .B(n759), .Z(n921) );
  INV_X1 U847 ( .A(n921), .ZN(n761) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U849 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U850 ( .A1(KEYINPUT33), .A2(n764), .ZN(n765) );
  NOR2_X1 U851 ( .A1(n935), .A2(n765), .ZN(n774) );
  AND2_X1 U852 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n767), .A2(n781), .ZN(n772) );
  XNOR2_X1 U854 ( .A(KEYINPUT86), .B(G1986), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(G290), .ZN(n925) );
  NOR2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n830) );
  NAND2_X1 U857 ( .A1(n925), .A2(n830), .ZN(n771) );
  AND2_X1 U858 ( .A1(n772), .A2(n520), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n786) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XNOR2_X1 U861 ( .A(n775), .B(KEYINPUT24), .ZN(n776) );
  AND2_X1 U862 ( .A1(n776), .A2(n781), .ZN(n784) );
  NAND2_X1 U863 ( .A1(G8), .A2(G166), .ZN(n777) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n777), .ZN(n778) );
  XOR2_X1 U865 ( .A(n778), .B(KEYINPUT106), .Z(n779) );
  AND2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n782) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n520), .A2(n519), .ZN(n785) );
  NAND2_X1 U869 ( .A1(n786), .A2(n785), .ZN(n819) );
  XNOR2_X1 U870 ( .A(KEYINPUT88), .B(KEYINPUT34), .ZN(n790) );
  NAND2_X1 U871 ( .A1(G140), .A2(n892), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G104), .A2(n890), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U874 ( .A(n790), .B(n789), .ZN(n795) );
  NAND2_X1 U875 ( .A1(G128), .A2(n886), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G116), .A2(n887), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U878 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  NOR2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U880 ( .A(KEYINPUT36), .B(n796), .ZN(n880) );
  XNOR2_X1 U881 ( .A(KEYINPUT37), .B(G2067), .ZN(n828) );
  NOR2_X1 U882 ( .A1(n880), .A2(n828), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n797), .B(KEYINPUT89), .ZN(n1010) );
  INV_X1 U884 ( .A(n1010), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n798), .A2(n830), .ZN(n827) );
  INV_X1 U886 ( .A(n827), .ZN(n817) );
  NAND2_X1 U887 ( .A1(G141), .A2(n892), .ZN(n805) );
  NAND2_X1 U888 ( .A1(G129), .A2(n886), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G117), .A2(n887), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n890), .A2(G105), .ZN(n801) );
  XOR2_X1 U892 ( .A(KEYINPUT38), .B(n801), .Z(n802) );
  NOR2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n806), .B(KEYINPUT90), .ZN(n883) );
  NAND2_X1 U896 ( .A1(n883), .A2(G1996), .ZN(n814) );
  NAND2_X1 U897 ( .A1(G119), .A2(n886), .ZN(n808) );
  NAND2_X1 U898 ( .A1(G131), .A2(n892), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U900 ( .A1(G107), .A2(n887), .ZN(n810) );
  NAND2_X1 U901 ( .A1(G95), .A2(n890), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n902) );
  NAND2_X1 U904 ( .A1(G1991), .A2(n902), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n990) );
  NAND2_X1 U906 ( .A1(n830), .A2(n990), .ZN(n815) );
  XNOR2_X1 U907 ( .A(KEYINPUT91), .B(n815), .ZN(n816) );
  NOR2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n833) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n883), .ZN(n820) );
  XOR2_X1 U911 ( .A(KEYINPUT107), .B(n820), .Z(n994) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n902), .ZN(n1005) );
  NOR2_X1 U914 ( .A1(n821), .A2(n1005), .ZN(n822) );
  NOR2_X1 U915 ( .A1(n990), .A2(n822), .ZN(n823) );
  NOR2_X1 U916 ( .A1(n994), .A2(n823), .ZN(n824) );
  XNOR2_X1 U917 ( .A(n824), .B(KEYINPUT108), .ZN(n825) );
  XNOR2_X1 U918 ( .A(n825), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n828), .A2(n880), .ZN(n991) );
  NAND2_X1 U921 ( .A1(n829), .A2(n991), .ZN(n831) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U924 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n835), .ZN(G217) );
  INV_X1 U926 ( .A(G661), .ZN(n837) );
  NAND2_X1 U927 ( .A1(G2), .A2(G15), .ZN(n836) );
  NOR2_X1 U928 ( .A1(n837), .A2(n836), .ZN(n838) );
  XOR2_X1 U929 ( .A(KEYINPUT112), .B(n838), .Z(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U933 ( .A(G132), .ZN(G219) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G82), .ZN(G220) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  INV_X1 U939 ( .A(n843), .ZN(G319) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n846), .B(G2100), .Z(n848) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2084), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U947 ( .A(KEYINPUT113), .B(G2678), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n852), .B(n851), .Z(G227) );
  XOR2_X1 U950 ( .A(KEYINPUT115), .B(G1956), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1981), .B(G1961), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n855), .B(KEYINPUT41), .Z(n857) );
  XNOR2_X1 U954 ( .A(G1991), .B(G1996), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1966), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(KEYINPUT114), .B(G2474), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G229) );
  XOR2_X1 U962 ( .A(KEYINPUT44), .B(KEYINPUT117), .Z(n865) );
  NAND2_X1 U963 ( .A1(G124), .A2(n886), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(KEYINPUT116), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n890), .A2(G100), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G112), .A2(n887), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G136), .A2(n892), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G139), .A2(n892), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G103), .A2(n890), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G127), .A2(n886), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G115), .A2(n887), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n996) );
  XNOR2_X1 U980 ( .A(G164), .B(n996), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n880), .B(G160), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(n905) );
  XOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n885) );
  XNOR2_X1 U984 ( .A(n883), .B(KEYINPUT119), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n901) );
  NAND2_X1 U986 ( .A1(G130), .A2(n886), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G118), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n897) );
  NAND2_X1 U989 ( .A1(n890), .A2(G106), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n891), .B(KEYINPUT118), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G142), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U993 ( .A(KEYINPUT45), .B(n895), .Z(n896) );
  NOR2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(G162), .B(n898), .Z(n899) );
  XNOR2_X1 U996 ( .A(n1002), .B(n899), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(n918), .B(n907), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(G171), .B(n923), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1004 ( .A(G286), .B(n910), .Z(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n912) );
  XOR2_X1 U1007 ( .A(KEYINPUT49), .B(n912), .Z(n913) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n913), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n914), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(KEYINPUT120), .B(n915), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G96), .ZN(G221) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1016 ( .A(KEYINPUT56), .B(G16), .ZN(n940) );
  XNOR2_X1 U1017 ( .A(G299), .B(G1956), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n918), .B(G1341), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n933) );
  XOR2_X1 U1021 ( .A(G1348), .B(n923), .Z(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(G1971), .A2(G303), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n929) );
  XOR2_X1 U1025 ( .A(G171), .B(G1961), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G168), .B(G1966), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT57), .B(n936), .Z(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT124), .B(n941), .ZN(n1019) );
  XNOR2_X1 U1035 ( .A(G21), .B(G1966), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n942), .B(KEYINPUT125), .ZN(n953) );
  XNOR2_X1 U1037 ( .A(G1971), .B(G22), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G1976), .B(G23), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1040 ( .A(KEYINPUT126), .B(n945), .Z(n947) );
  XNOR2_X1 U1041 ( .A(G1986), .B(G24), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT58), .B(n948), .Z(n951) );
  XNOR2_X1 U1044 ( .A(n949), .B(G5), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n963) );
  XOR2_X1 U1047 ( .A(G1348), .B(KEYINPUT59), .Z(n954) );
  XNOR2_X1 U1048 ( .A(G4), .B(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G20), .B(G1956), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(G1981), .B(G6), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G1341), .B(G19), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT60), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n964), .Z(n965) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n965), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT127), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(G11), .ZN(n1017) );
  XOR2_X1 U1061 ( .A(n968), .B(G27), .Z(n973) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G26), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G2072), .B(G33), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT121), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(KEYINPUT122), .B(G32), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT123), .B(n978), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n979), .A2(G28), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G25), .B(G1991), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(KEYINPUT53), .B(n982), .Z(n985) );
  XOR2_X1 U1075 ( .A(G34), .B(KEYINPUT54), .Z(n983) );
  XNOR2_X1 U1076 ( .A(G2084), .B(n983), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(G35), .B(G2090), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(G29), .A2(n988), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n989), .B(KEYINPUT55), .ZN(n1015) );
  INV_X1 U1082 ( .A(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1009) );
  XOR2_X1 U1084 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1086 ( .A(KEYINPUT51), .B(n995), .Z(n1007) );
  XOR2_X1 U1087 ( .A(G2072), .B(n996), .Z(n998) );
  XOR2_X1 U1088 ( .A(G164), .B(G2078), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1090 ( .A(KEYINPUT50), .B(n999), .Z(n1001) );
  XOR2_X1 U1091 ( .A(G160), .B(G2084), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(G29), .A2(n1013), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

