

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  NOR2_X1 U324 ( .A1(n537), .A2(n484), .ZN(n428) );
  XNOR2_X1 U325 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U326 ( .A(n300), .B(n299), .ZN(n303) );
  XOR2_X1 U327 ( .A(n313), .B(n312), .Z(n581) );
  XOR2_X1 U328 ( .A(n581), .B(KEYINPUT41), .Z(n557) );
  NOR2_X1 U329 ( .A1(n542), .A2(n454), .ZN(n569) );
  XNOR2_X1 U330 ( .A(n455), .B(KEYINPUT121), .ZN(n456) );
  XOR2_X1 U331 ( .A(n333), .B(n332), .Z(n542) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(n459) );
  INV_X1 U333 ( .A(KEYINPUT107), .ZN(n314) );
  XOR2_X1 U334 ( .A(KEYINPUT72), .B(G78GAT), .Z(n293) );
  XNOR2_X1 U335 ( .A(G148GAT), .B(G106GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n346) );
  INV_X1 U337 ( .A(KEYINPUT33), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n346), .B(n294), .ZN(n296) );
  NAND2_X1 U339 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U341 ( .A(G85GAT), .B(G99GAT), .Z(n380) );
  XNOR2_X1 U342 ( .A(G120GAT), .B(n380), .ZN(n298) );
  INV_X1 U343 ( .A(KEYINPUT31), .ZN(n297) );
  XOR2_X1 U344 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n302) );
  XNOR2_X1 U345 ( .A(KEYINPUT32), .B(KEYINPUT74), .ZN(n301) );
  XOR2_X1 U346 ( .A(n302), .B(n301), .Z(n304) );
  NAND2_X1 U347 ( .A1(n303), .A2(n304), .ZN(n308) );
  INV_X1 U348 ( .A(n303), .ZN(n306) );
  INV_X1 U349 ( .A(n304), .ZN(n305) );
  NAND2_X1 U350 ( .A1(n306), .A2(n305), .ZN(n307) );
  NAND2_X1 U351 ( .A1(n308), .A2(n307), .ZN(n313) );
  XNOR2_X1 U352 ( .A(G57GAT), .B(G71GAT), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n309), .B(KEYINPUT13), .ZN(n398) );
  XOR2_X1 U354 ( .A(G204GAT), .B(G176GAT), .Z(n311) );
  XNOR2_X1 U355 ( .A(G92GAT), .B(G64GAT), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n422) );
  XNOR2_X1 U357 ( .A(n398), .B(n422), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n314), .B(n557), .ZN(n510) );
  XOR2_X1 U359 ( .A(G127GAT), .B(G15GAT), .Z(n400) );
  XOR2_X1 U360 ( .A(KEYINPUT87), .B(G99GAT), .Z(n316) );
  XNOR2_X1 U361 ( .A(G43GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U363 ( .A(n400), .B(n317), .Z(n319) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n333) );
  XOR2_X1 U366 ( .A(G176GAT), .B(G169GAT), .Z(n321) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n323) );
  XNOR2_X1 U370 ( .A(G71GAT), .B(KEYINPUT86), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U372 ( .A(n325), .B(n324), .Z(n331) );
  XOR2_X1 U373 ( .A(G120GAT), .B(KEYINPUT83), .Z(n327) );
  XNOR2_X1 U374 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n435) );
  XOR2_X1 U376 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n329) );
  XNOR2_X1 U377 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n427) );
  XNOR2_X1 U379 ( .A(n435), .B(n427), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U381 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n335) );
  XNOR2_X1 U382 ( .A(KEYINPUT2), .B(G141GAT), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U384 ( .A(KEYINPUT3), .B(n336), .Z(n449) );
  XOR2_X1 U385 ( .A(G197GAT), .B(KEYINPUT21), .Z(n338) );
  XNOR2_X1 U386 ( .A(G218GAT), .B(G211GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n417) );
  XOR2_X1 U388 ( .A(KEYINPUT23), .B(n417), .Z(n340) );
  XOR2_X1 U389 ( .A(G155GAT), .B(G22GAT), .Z(n401) );
  XNOR2_X1 U390 ( .A(n401), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n449), .B(n341), .ZN(n350) );
  XOR2_X1 U393 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n343) );
  NAND2_X1 U394 ( .A1(G228GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U396 ( .A(n344), .B(KEYINPUT88), .Z(n348) );
  XNOR2_X1 U397 ( .A(G162GAT), .B(G50GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n345), .B(KEYINPUT76), .ZN(n382) );
  XNOR2_X1 U399 ( .A(n382), .B(n346), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U401 ( .A(n350), .B(n349), .Z(n465) );
  INV_X1 U402 ( .A(n581), .ZN(n460) );
  XOR2_X1 U403 ( .A(KEYINPUT7), .B(G43GAT), .Z(n352) );
  XNOR2_X1 U404 ( .A(G29GAT), .B(KEYINPUT69), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U406 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n353) );
  XOR2_X1 U407 ( .A(n354), .B(n353), .Z(n385) );
  XOR2_X1 U408 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n356) );
  NAND2_X1 U409 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U411 ( .A(KEYINPUT67), .B(n357), .ZN(n367) );
  XOR2_X1 U412 ( .A(G8GAT), .B(G169GAT), .Z(n420) );
  XOR2_X1 U413 ( .A(n420), .B(G36GAT), .Z(n359) );
  XOR2_X1 U414 ( .A(G113GAT), .B(G1GAT), .Z(n436) );
  XNOR2_X1 U415 ( .A(n436), .B(G50GAT), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U417 ( .A(KEYINPUT66), .B(KEYINPUT68), .Z(n361) );
  XNOR2_X1 U418 ( .A(G15GAT), .B(G197GAT), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U420 ( .A(n363), .B(n362), .Z(n365) );
  XNOR2_X1 U421 ( .A(G141GAT), .B(G22GAT), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n385), .B(n368), .ZN(n578) );
  XOR2_X1 U425 ( .A(G92GAT), .B(G106GAT), .Z(n370) );
  XNOR2_X1 U426 ( .A(G134GAT), .B(G218GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U428 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n372) );
  XNOR2_X1 U429 ( .A(KEYINPUT77), .B(KEYINPUT10), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U431 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U432 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n376) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U435 ( .A(KEYINPUT78), .B(n377), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n384) );
  XOR2_X1 U438 ( .A(G190GAT), .B(G36GAT), .Z(n423) );
  XNOR2_X1 U439 ( .A(n382), .B(n423), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n386) );
  XOR2_X1 U441 ( .A(n386), .B(n385), .Z(n568) );
  XNOR2_X1 U442 ( .A(KEYINPUT36), .B(n568), .ZN(n588) );
  XOR2_X1 U443 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n388) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U446 ( .A(n389), .B(KEYINPUT12), .Z(n397) );
  XOR2_X1 U447 ( .A(G183GAT), .B(G211GAT), .Z(n391) );
  XNOR2_X1 U448 ( .A(G1GAT), .B(G78GAT), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U450 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n393) );
  XNOR2_X1 U451 ( .A(G64GAT), .B(G8GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n399) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n403) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n585) );
  NAND2_X1 U458 ( .A1(n588), .A2(n585), .ZN(n404) );
  XNOR2_X1 U459 ( .A(KEYINPUT45), .B(n404), .ZN(n405) );
  NOR2_X1 U460 ( .A1(n578), .A2(n405), .ZN(n406) );
  NAND2_X1 U461 ( .A1(n460), .A2(n406), .ZN(n415) );
  NAND2_X1 U462 ( .A1(n557), .A2(n578), .ZN(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n411) );
  INV_X1 U465 ( .A(n585), .ZN(n493) );
  INV_X1 U466 ( .A(n568), .ZN(n409) );
  NAND2_X1 U467 ( .A1(n493), .A2(n409), .ZN(n410) );
  NOR2_X1 U468 ( .A1(n411), .A2(n410), .ZN(n413) );
  XNOR2_X1 U469 ( .A(KEYINPUT47), .B(KEYINPUT116), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n414) );
  NAND2_X1 U471 ( .A1(n415), .A2(n414), .ZN(n416) );
  XOR2_X1 U472 ( .A(n416), .B(KEYINPUT48), .Z(n537) );
  XOR2_X1 U473 ( .A(KEYINPUT97), .B(n417), .Z(n419) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n421) );
  XOR2_X1 U476 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U479 ( .A(n427), .B(n426), .Z(n484) );
  XNOR2_X1 U480 ( .A(n428), .B(KEYINPUT54), .ZN(n452) );
  XOR2_X1 U481 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n430) );
  XNOR2_X1 U482 ( .A(KEYINPUT5), .B(KEYINPUT96), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U484 ( .A(KEYINPUT92), .B(n431), .Z(n433) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U487 ( .A(n434), .B(KEYINPUT95), .Z(n441) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n438) );
  XNOR2_X1 U489 ( .A(G162GAT), .B(G85GAT), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n439), .B(KEYINPUT6), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U493 ( .A(G127GAT), .B(G148GAT), .Z(n443) );
  XNOR2_X1 U494 ( .A(G29GAT), .B(G155GAT), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U496 ( .A(n445), .B(n444), .Z(n451) );
  XOR2_X1 U497 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n447) );
  XNOR2_X1 U498 ( .A(G57GAT), .B(KEYINPUT93), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U501 ( .A(n451), .B(n450), .Z(n499) );
  NAND2_X1 U502 ( .A1(n452), .A2(n499), .ZN(n575) );
  NOR2_X1 U503 ( .A1(n465), .A2(n575), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT55), .ZN(n454) );
  AND2_X1 U505 ( .A1(n510), .A2(n569), .ZN(n457) );
  XNOR2_X1 U506 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n455) );
  XOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .Z(n458) );
  XNOR2_X1 U508 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  NAND2_X1 U509 ( .A1(n578), .A2(n460), .ZN(n461) );
  XNOR2_X1 U510 ( .A(n461), .B(KEYINPUT75), .ZN(n497) );
  INV_X1 U511 ( .A(n542), .ZN(n531) );
  INV_X1 U512 ( .A(n484), .ZN(n529) );
  NAND2_X1 U513 ( .A1(n531), .A2(n529), .ZN(n462) );
  XNOR2_X1 U514 ( .A(KEYINPUT98), .B(n462), .ZN(n463) );
  INV_X1 U515 ( .A(n465), .ZN(n471) );
  NAND2_X1 U516 ( .A1(n463), .A2(n471), .ZN(n464) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(n464), .ZN(n468) );
  NAND2_X1 U518 ( .A1(n542), .A2(n465), .ZN(n466) );
  XNOR2_X1 U519 ( .A(KEYINPUT26), .B(n466), .ZN(n576) );
  XOR2_X1 U520 ( .A(n529), .B(KEYINPUT27), .Z(n472) );
  NOR2_X1 U521 ( .A1(n576), .A2(n472), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT99), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n470), .A2(n499), .ZN(n475) );
  XOR2_X1 U525 ( .A(KEYINPUT28), .B(n471), .Z(n540) );
  OR2_X1 U526 ( .A1(n499), .A2(n472), .ZN(n538) );
  NOR2_X1 U527 ( .A1(n540), .A2(n538), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n542), .A2(n473), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n475), .A2(n474), .ZN(n492) );
  XNOR2_X1 U530 ( .A(KEYINPUT16), .B(KEYINPUT82), .ZN(n476) );
  XNOR2_X1 U531 ( .A(n476), .B(KEYINPUT81), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n568), .A2(n493), .ZN(n477) );
  XOR2_X1 U533 ( .A(n478), .B(n477), .Z(n479) );
  NAND2_X1 U534 ( .A1(n492), .A2(n479), .ZN(n480) );
  XOR2_X1 U535 ( .A(KEYINPUT100), .B(n480), .Z(n511) );
  NAND2_X1 U536 ( .A1(n497), .A2(n511), .ZN(n489) );
  NOR2_X1 U537 ( .A1(n499), .A2(n489), .ZN(n482) );
  XNOR2_X1 U538 ( .A(KEYINPUT101), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U541 ( .A1(n484), .A2(n489), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT102), .B(n485), .Z(n486) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n542), .A2(n489), .ZN(n488) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  INV_X1 U547 ( .A(n540), .ZN(n490) );
  NOR2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  NAND2_X1 U550 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U551 ( .A(n494), .B(KEYINPUT103), .ZN(n495) );
  NAND2_X1 U552 ( .A1(n495), .A2(n588), .ZN(n496) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n496), .ZN(n525) );
  NAND2_X1 U554 ( .A1(n497), .A2(n525), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n498), .Z(n507) );
  INV_X1 U556 ( .A(n499), .ZN(n527) );
  NAND2_X1 U557 ( .A1(n507), .A2(n527), .ZN(n502) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT104), .Z(n500) );
  XNOR2_X1 U559 ( .A(KEYINPUT39), .B(n500), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XOR2_X1 U561 ( .A(G36GAT), .B(KEYINPUT105), .Z(n504) );
  NAND2_X1 U562 ( .A1(n507), .A2(n529), .ZN(n503) );
  XNOR2_X1 U563 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n507), .A2(n531), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U567 ( .A1(n507), .A2(n540), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n508), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(n509), .ZN(G1331GAT) );
  INV_X1 U570 ( .A(n510), .ZN(n545) );
  NOR2_X1 U571 ( .A1(n545), .A2(n578), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n511), .A2(n524), .ZN(n512) );
  XOR2_X1 U573 ( .A(KEYINPUT108), .B(n512), .Z(n519) );
  NAND2_X1 U574 ( .A1(n519), .A2(n527), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n513), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  XOR2_X1 U577 ( .A(G64GAT), .B(KEYINPUT109), .Z(n516) );
  NAND2_X1 U578 ( .A1(n519), .A2(n529), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n519), .A2(n531), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U584 ( .A1(n540), .A2(n519), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n523) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT111), .Z(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(KEYINPUT113), .B(n526), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n527), .A2(n533), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n533), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n533), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n535) );
  NAND2_X1 U597 ( .A1(n533), .A2(n540), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  NOR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U601 ( .A(KEYINPUT117), .B(n539), .ZN(n554) );
  OR2_X1 U602 ( .A1(n554), .A2(n540), .ZN(n541) );
  NOR2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n551), .A2(n578), .ZN(n543) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  INV_X1 U606 ( .A(n551), .ZN(n544) );
  NOR2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n549) );
  NAND2_X1 U611 ( .A1(n551), .A2(n585), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U613 ( .A(G127GAT), .B(n550), .Z(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U615 ( .A1(n551), .A2(n568), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  XOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT119), .Z(n556) );
  NOR2_X1 U618 ( .A1(n576), .A2(n554), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n562), .A2(n578), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U622 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n585), .A2(n562), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n568), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n578), .A2(n569), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT120), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT123), .Z(n567) );
  NAND2_X1 U633 ( .A1(n569), .A2(n585), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n571) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G190GAT), .B(n572), .Z(G1351GAT) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(KEYINPUT59), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(n574), .Z(n580) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(n577), .Z(n587) );
  NAND2_X1 U644 ( .A1(n587), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n584), .Z(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

