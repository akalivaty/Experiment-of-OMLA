

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U545 ( .A1(n781), .A2(n779), .ZN(n736) );
  XNOR2_X1 U546 ( .A(n682), .B(n681), .ZN(n779) );
  NAND2_X1 U547 ( .A1(n867), .A2(G137), .ZN(n528) );
  NOR2_X1 U548 ( .A1(n689), .A2(n905), .ZN(n691) );
  XNOR2_X1 U549 ( .A(n712), .B(n711), .ZN(n716) );
  NAND2_X1 U550 ( .A1(n710), .A2(n709), .ZN(n712) );
  XOR2_X1 U551 ( .A(KEYINPUT1), .B(n516), .Z(n645) );
  NOR2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X1 U553 ( .A(KEYINPUT101), .B(n765), .Z(n509) );
  INV_X1 U554 ( .A(n736), .ZN(n700) );
  INV_X1 U555 ( .A(KEYINPUT64), .ZN(n690) );
  XNOR2_X1 U556 ( .A(n691), .B(n690), .ZN(n697) );
  XNOR2_X1 U557 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n719) );
  XNOR2_X1 U558 ( .A(n720), .B(n719), .ZN(n721) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n711) );
  XNOR2_X1 U560 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n725) );
  XNOR2_X1 U561 ( .A(n685), .B(n684), .ZN(n717) );
  AND2_X1 U562 ( .A1(n729), .A2(n735), .ZN(n730) );
  AND2_X1 U563 ( .A1(n743), .A2(n742), .ZN(n745) );
  XNOR2_X1 U564 ( .A(KEYINPUT92), .B(n683), .ZN(n764) );
  AND2_X1 U565 ( .A1(G40), .A2(n680), .ZN(n682) );
  INV_X1 U566 ( .A(KEYINPUT17), .ZN(n526) );
  NOR2_X1 U567 ( .A1(n801), .A2(n800), .ZN(n804) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n640) );
  AND2_X2 U569 ( .A1(n532), .A2(G2104), .ZN(n868) );
  NOR2_X1 U570 ( .A1(G651), .A2(n634), .ZN(n644) );
  NOR2_X1 U571 ( .A1(n536), .A2(n535), .ZN(n680) );
  BUF_X1 U572 ( .A(n680), .Z(G160) );
  NAND2_X1 U573 ( .A1(G89), .A2(n640), .ZN(n510) );
  XOR2_X1 U574 ( .A(KEYINPUT75), .B(n510), .Z(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT4), .ZN(n513) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  XOR2_X1 U577 ( .A(G651), .B(KEYINPUT68), .Z(n515) );
  NOR2_X1 U578 ( .A1(n634), .A2(n515), .ZN(n641) );
  NAND2_X1 U579 ( .A1(G76), .A2(n641), .ZN(n512) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(KEYINPUT5), .B(n514), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n644), .A2(G51), .ZN(n518) );
  NOR2_X1 U583 ( .A1(G543), .A2(n515), .ZN(n516) );
  NAND2_X1 U584 ( .A1(G63), .A2(n645), .ZN(n517) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT76), .B(KEYINPUT6), .Z(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT7), .B(n523), .ZN(G168) );
  INV_X1 U590 ( .A(G2105), .ZN(n532) );
  NAND2_X1 U591 ( .A1(G101), .A2(n868), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n524), .B(KEYINPUT65), .ZN(n525) );
  XNOR2_X1 U593 ( .A(KEYINPUT23), .B(n525), .ZN(n530) );
  XNOR2_X2 U594 ( .A(n527), .B(n526), .ZN(n867) );
  XOR2_X1 U595 ( .A(n528), .B(KEYINPUT67), .Z(n529) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n536) );
  NAND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XOR2_X2 U598 ( .A(KEYINPUT66), .B(n531), .Z(n871) );
  NAND2_X1 U599 ( .A1(G113), .A2(n871), .ZN(n534) );
  NOR2_X1 U600 ( .A1(G2104), .A2(n532), .ZN(n873) );
  NAND2_X1 U601 ( .A1(n873), .A2(G125), .ZN(n533) );
  NAND2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U603 ( .A1(G138), .A2(n867), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(KEYINPUT86), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n868), .A2(G102), .ZN(n538) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U607 ( .A1(n873), .A2(G126), .ZN(n541) );
  NAND2_X1 U608 ( .A1(G114), .A2(n871), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(G164) );
  NAND2_X1 U611 ( .A1(n640), .A2(G91), .ZN(n545) );
  NAND2_X1 U612 ( .A1(G65), .A2(n645), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n644), .A2(G53), .ZN(n547) );
  NAND2_X1 U615 ( .A1(G78), .A2(n641), .ZN(n546) );
  NAND2_X1 U616 ( .A1(n547), .A2(n546), .ZN(n548) );
  OR2_X1 U617 ( .A1(n549), .A2(n548), .ZN(G299) );
  NAND2_X1 U618 ( .A1(n640), .A2(G85), .ZN(n551) );
  NAND2_X1 U619 ( .A1(G60), .A2(n645), .ZN(n550) );
  NAND2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n644), .A2(G47), .ZN(n553) );
  NAND2_X1 U622 ( .A1(G72), .A2(n641), .ZN(n552) );
  NAND2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n554) );
  OR2_X1 U624 ( .A1(n555), .A2(n554), .ZN(G290) );
  XOR2_X1 U625 ( .A(G2430), .B(G2451), .Z(n557) );
  XNOR2_X1 U626 ( .A(KEYINPUT103), .B(G2443), .ZN(n556) );
  XNOR2_X1 U627 ( .A(n557), .B(n556), .ZN(n564) );
  XOR2_X1 U628 ( .A(G2435), .B(G2446), .Z(n559) );
  XNOR2_X1 U629 ( .A(G2427), .B(G2454), .ZN(n558) );
  XNOR2_X1 U630 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U631 ( .A(n560), .B(G2438), .Z(n562) );
  XNOR2_X1 U632 ( .A(G1348), .B(G1341), .ZN(n561) );
  XNOR2_X1 U633 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U634 ( .A(n564), .B(n563), .ZN(n565) );
  AND2_X1 U635 ( .A1(n565), .A2(G14), .ZN(G401) );
  AND2_X1 U636 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U637 ( .A(G132), .ZN(G219) );
  INV_X1 U638 ( .A(G69), .ZN(G235) );
  NAND2_X1 U639 ( .A1(n644), .A2(G52), .ZN(n567) );
  NAND2_X1 U640 ( .A1(G64), .A2(n645), .ZN(n566) );
  NAND2_X1 U641 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U642 ( .A1(G90), .A2(n640), .ZN(n569) );
  NAND2_X1 U643 ( .A1(G77), .A2(n641), .ZN(n568) );
  NAND2_X1 U644 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U645 ( .A(KEYINPUT9), .B(n570), .Z(n571) );
  NOR2_X1 U646 ( .A1(n572), .A2(n571), .ZN(G171) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U649 ( .A(n573), .B(KEYINPUT70), .ZN(n574) );
  XNOR2_X1 U650 ( .A(KEYINPUT10), .B(n574), .ZN(G223) );
  INV_X1 U651 ( .A(G223), .ZN(n821) );
  NAND2_X1 U652 ( .A1(n821), .A2(G567), .ZN(n575) );
  XNOR2_X1 U653 ( .A(n575), .B(KEYINPUT71), .ZN(n576) );
  XNOR2_X1 U654 ( .A(KEYINPUT11), .B(n576), .ZN(G234) );
  XOR2_X1 U655 ( .A(G860), .B(KEYINPUT72), .Z(n599) );
  NAND2_X1 U656 ( .A1(n645), .A2(G56), .ZN(n577) );
  XOR2_X1 U657 ( .A(KEYINPUT14), .B(n577), .Z(n583) );
  NAND2_X1 U658 ( .A1(n640), .A2(G81), .ZN(n578) );
  XNOR2_X1 U659 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U660 ( .A1(G68), .A2(n641), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U662 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U663 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n644), .A2(G43), .ZN(n584) );
  NAND2_X1 U665 ( .A1(n585), .A2(n584), .ZN(n905) );
  OR2_X1 U666 ( .A1(n599), .A2(n905), .ZN(G153) );
  INV_X1 U667 ( .A(G171), .ZN(G301) );
  NAND2_X1 U668 ( .A1(G66), .A2(n645), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G92), .A2(n640), .ZN(n587) );
  NAND2_X1 U670 ( .A1(G54), .A2(n644), .ZN(n586) );
  NAND2_X1 U671 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U672 ( .A1(G79), .A2(n641), .ZN(n588) );
  XNOR2_X1 U673 ( .A(KEYINPUT73), .B(n588), .ZN(n589) );
  NOR2_X1 U674 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U675 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U676 ( .A(KEYINPUT15), .B(n593), .Z(n696) );
  INV_X1 U677 ( .A(G868), .ZN(n658) );
  NAND2_X1 U678 ( .A1(n696), .A2(n658), .ZN(n594) );
  XNOR2_X1 U679 ( .A(n594), .B(KEYINPUT74), .ZN(n596) );
  NAND2_X1 U680 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U681 ( .A1(n596), .A2(n595), .ZN(G284) );
  NOR2_X1 U682 ( .A1(G286), .A2(n658), .ZN(n598) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U684 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n599), .A2(G559), .ZN(n600) );
  INV_X1 U686 ( .A(n696), .ZN(n910) );
  NAND2_X1 U687 ( .A1(n600), .A2(n910), .ZN(n601) );
  XNOR2_X1 U688 ( .A(n601), .B(KEYINPUT77), .ZN(n602) );
  XOR2_X1 U689 ( .A(KEYINPUT16), .B(n602), .Z(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n905), .ZN(n603) );
  XNOR2_X1 U691 ( .A(KEYINPUT78), .B(n603), .ZN(n606) );
  NAND2_X1 U692 ( .A1(G868), .A2(n910), .ZN(n604) );
  NOR2_X1 U693 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U694 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U695 ( .A1(n868), .A2(G99), .ZN(n607) );
  XOR2_X1 U696 ( .A(KEYINPUT79), .B(n607), .Z(n609) );
  NAND2_X1 U697 ( .A1(G111), .A2(n871), .ZN(n608) );
  NAND2_X1 U698 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U699 ( .A(KEYINPUT80), .B(n610), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G123), .A2(n873), .ZN(n611) );
  XNOR2_X1 U701 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U702 ( .A1(n867), .A2(G135), .ZN(n612) );
  NAND2_X1 U703 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U704 ( .A1(n615), .A2(n614), .ZN(n959) );
  XNOR2_X1 U705 ( .A(n959), .B(G2096), .ZN(n617) );
  INV_X1 U706 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U707 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U708 ( .A1(n640), .A2(G93), .ZN(n619) );
  NAND2_X1 U709 ( .A1(G67), .A2(n645), .ZN(n618) );
  NAND2_X1 U710 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U711 ( .A1(G55), .A2(n644), .ZN(n620) );
  XNOR2_X1 U712 ( .A(KEYINPUT81), .B(n620), .ZN(n621) );
  NOR2_X1 U713 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U714 ( .A1(G80), .A2(n641), .ZN(n623) );
  NAND2_X1 U715 ( .A1(n624), .A2(n623), .ZN(n660) );
  NAND2_X1 U716 ( .A1(n910), .A2(G559), .ZN(n656) );
  XNOR2_X1 U717 ( .A(n905), .B(n656), .ZN(n625) );
  NOR2_X1 U718 ( .A1(G860), .A2(n625), .ZN(n626) );
  XOR2_X1 U719 ( .A(n660), .B(n626), .Z(G145) );
  NAND2_X1 U720 ( .A1(G86), .A2(n640), .ZN(n628) );
  NAND2_X1 U721 ( .A1(G48), .A2(n644), .ZN(n627) );
  NAND2_X1 U722 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U723 ( .A1(n641), .A2(G73), .ZN(n629) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U725 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U726 ( .A1(G61), .A2(n645), .ZN(n632) );
  NAND2_X1 U727 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U728 ( .A1(G87), .A2(n634), .ZN(n636) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U730 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U731 ( .A1(n645), .A2(n637), .ZN(n639) );
  NAND2_X1 U732 ( .A1(n644), .A2(G49), .ZN(n638) );
  NAND2_X1 U733 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U734 ( .A1(G88), .A2(n640), .ZN(n643) );
  NAND2_X1 U735 ( .A1(G75), .A2(n641), .ZN(n642) );
  NAND2_X1 U736 ( .A1(n643), .A2(n642), .ZN(n649) );
  NAND2_X1 U737 ( .A1(n644), .A2(G50), .ZN(n647) );
  NAND2_X1 U738 ( .A1(G62), .A2(n645), .ZN(n646) );
  NAND2_X1 U739 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U740 ( .A1(n649), .A2(n648), .ZN(G166) );
  XOR2_X1 U741 ( .A(G305), .B(n905), .Z(n650) );
  XNOR2_X1 U742 ( .A(n660), .B(n650), .ZN(n651) );
  XNOR2_X1 U743 ( .A(KEYINPUT19), .B(n651), .ZN(n653) );
  XNOR2_X1 U744 ( .A(G288), .B(G166), .ZN(n652) );
  XNOR2_X1 U745 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U746 ( .A(n654), .B(G299), .Z(n655) );
  XNOR2_X1 U747 ( .A(G290), .B(n655), .ZN(n892) );
  XNOR2_X1 U748 ( .A(KEYINPUT82), .B(n892), .ZN(n657) );
  XNOR2_X1 U749 ( .A(n657), .B(n656), .ZN(n659) );
  NOR2_X1 U750 ( .A1(n659), .A2(n658), .ZN(n662) );
  NOR2_X1 U751 ( .A1(G868), .A2(n660), .ZN(n661) );
  NOR2_X1 U752 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U757 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U759 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NAND2_X1 U760 ( .A1(G120), .A2(G57), .ZN(n667) );
  NOR2_X1 U761 ( .A1(G235), .A2(n667), .ZN(n668) );
  XNOR2_X1 U762 ( .A(KEYINPUT84), .B(n668), .ZN(n669) );
  NAND2_X1 U763 ( .A1(n669), .A2(G108), .ZN(n826) );
  NAND2_X1 U764 ( .A1(n826), .A2(G567), .ZN(n675) );
  NOR2_X1 U765 ( .A1(G219), .A2(G220), .ZN(n670) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U767 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U768 ( .A1(G96), .A2(n672), .ZN(n827) );
  NAND2_X1 U769 ( .A1(G2106), .A2(n827), .ZN(n673) );
  XOR2_X1 U770 ( .A(KEYINPUT83), .B(n673), .Z(n674) );
  NAND2_X1 U771 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U772 ( .A(n676), .B(KEYINPUT85), .ZN(G319) );
  INV_X1 U773 ( .A(G319), .ZN(n678) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n677) );
  NOR2_X1 U775 ( .A1(n678), .A2(n677), .ZN(n825) );
  NAND2_X1 U776 ( .A1(n825), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U778 ( .A(KEYINPUT100), .B(G1981), .ZN(n679) );
  XNOR2_X1 U779 ( .A(n679), .B(G305), .ZN(n902) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n781) );
  INV_X1 U781 ( .A(KEYINPUT87), .ZN(n681) );
  NAND2_X1 U782 ( .A1(G8), .A2(n736), .ZN(n683) );
  NOR2_X1 U783 ( .A1(n764), .A2(G1966), .ZN(n685) );
  INV_X1 U784 ( .A(KEYINPUT93), .ZN(n684) );
  INV_X1 U785 ( .A(n717), .ZN(n729) );
  XNOR2_X1 U786 ( .A(KEYINPUT94), .B(G1996), .ZN(n931) );
  NAND2_X1 U787 ( .A1(n931), .A2(n700), .ZN(n686) );
  XNOR2_X1 U788 ( .A(n686), .B(KEYINPUT26), .ZN(n688) );
  NAND2_X1 U789 ( .A1(n736), .A2(G1341), .ZN(n687) );
  NAND2_X1 U790 ( .A1(n688), .A2(n687), .ZN(n689) );
  OR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n695) );
  NOR2_X1 U792 ( .A1(G2067), .A2(n736), .ZN(n693) );
  NOR2_X1 U793 ( .A1(n700), .A2(G1348), .ZN(n692) );
  NOR2_X1 U794 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U795 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n700), .A2(G2072), .ZN(n701) );
  XOR2_X1 U799 ( .A(KEYINPUT27), .B(n701), .Z(n703) );
  NAND2_X1 U800 ( .A1(G1956), .A2(n736), .ZN(n702) );
  NAND2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U802 ( .A1(G299), .A2(n707), .ZN(n704) );
  XNOR2_X1 U803 ( .A(n704), .B(KEYINPUT95), .ZN(n705) );
  NAND2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U805 ( .A1(G299), .A2(n707), .ZN(n708) );
  XNOR2_X1 U806 ( .A(n708), .B(KEYINPUT28), .ZN(n709) );
  XNOR2_X1 U807 ( .A(KEYINPUT25), .B(G2078), .ZN(n937) );
  NOR2_X1 U808 ( .A1(n736), .A2(n937), .ZN(n714) );
  AND2_X1 U809 ( .A1(n736), .A2(G1961), .ZN(n713) );
  NOR2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n722) );
  NAND2_X1 U811 ( .A1(G171), .A2(n722), .ZN(n715) );
  NAND2_X1 U812 ( .A1(n716), .A2(n715), .ZN(n728) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n736), .ZN(n731) );
  NOR2_X1 U814 ( .A1(n717), .A2(n731), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n718), .A2(G8), .ZN(n720) );
  NOR2_X1 U816 ( .A1(n721), .A2(G168), .ZN(n724) );
  NOR2_X1 U817 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n726) );
  XNOR2_X1 U819 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n735) );
  XNOR2_X1 U821 ( .A(n730), .B(KEYINPUT98), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n731), .A2(G8), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n747) );
  AND2_X1 U824 ( .A1(G286), .A2(G8), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n743) );
  INV_X1 U826 ( .A(G8), .ZN(n741) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n736), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n764), .A2(G1971), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U830 ( .A1(G303), .A2(n739), .ZN(n740) );
  OR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U832 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n744) );
  XNOR2_X1 U833 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n762) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U836 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n753), .A2(n748), .ZN(n918) );
  NAND2_X1 U838 ( .A1(n762), .A2(n918), .ZN(n749) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n914) );
  NAND2_X1 U840 ( .A1(n749), .A2(n914), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n750), .A2(n764), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n902), .A2(n752), .ZN(n756) );
  AND2_X1 U844 ( .A1(n753), .A2(KEYINPUT33), .ZN(n754) );
  INV_X1 U845 ( .A(n764), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n754), .A2(n758), .ZN(n755) );
  AND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n768) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XNOR2_X1 U849 ( .A(n757), .B(KEYINPUT24), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n766) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U852 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n509), .ZN(n767) );
  NOR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n801) );
  NAND2_X1 U857 ( .A1(G140), .A2(n867), .ZN(n770) );
  NAND2_X1 U858 ( .A1(G104), .A2(n868), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n771), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G116), .A2(n871), .ZN(n772) );
  XOR2_X1 U862 ( .A(KEYINPUT89), .B(n772), .Z(n774) );
  NAND2_X1 U863 ( .A1(n873), .A2(G128), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  NOR2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n778), .ZN(n887) );
  XNOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .ZN(n814) );
  NOR2_X1 U869 ( .A1(n887), .A2(n814), .ZN(n970) );
  INV_X1 U870 ( .A(n779), .ZN(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n816) );
  NAND2_X1 U872 ( .A1(n970), .A2(n816), .ZN(n813) );
  NAND2_X1 U873 ( .A1(G95), .A2(n868), .ZN(n783) );
  NAND2_X1 U874 ( .A1(G107), .A2(n871), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G131), .A2(n867), .ZN(n785) );
  NAND2_X1 U877 ( .A1(G119), .A2(n873), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n864) );
  INV_X1 U880 ( .A(G1991), .ZN(n928) );
  NOR2_X1 U881 ( .A1(n864), .A2(n928), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G105), .A2(n868), .ZN(n788) );
  XNOR2_X1 U883 ( .A(n788), .B(KEYINPUT38), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G129), .A2(n873), .ZN(n789) );
  XNOR2_X1 U885 ( .A(n789), .B(KEYINPUT90), .ZN(n791) );
  NAND2_X1 U886 ( .A1(G117), .A2(n871), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U888 ( .A1(G141), .A2(n867), .ZN(n792) );
  XNOR2_X1 U889 ( .A(KEYINPUT91), .B(n792), .ZN(n793) );
  NOR2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n881) );
  AND2_X1 U892 ( .A1(G1996), .A2(n881), .ZN(n797) );
  NOR2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n963) );
  INV_X1 U894 ( .A(n963), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n799), .A2(n816), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n813), .A2(n805), .ZN(n800) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n920) );
  NAND2_X1 U898 ( .A1(n920), .A2(n816), .ZN(n802) );
  XNOR2_X1 U899 ( .A(n802), .B(KEYINPUT88), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n819) );
  XOR2_X1 U901 ( .A(KEYINPUT39), .B(KEYINPUT102), .Z(n811) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n881), .ZN(n957) );
  INV_X1 U903 ( .A(n805), .ZN(n808) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n806) );
  AND2_X1 U905 ( .A1(n928), .A2(n864), .ZN(n960) );
  NOR2_X1 U906 ( .A1(n806), .A2(n960), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n957), .A2(n809), .ZN(n810) );
  XOR2_X1 U909 ( .A(n811), .B(n810), .Z(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n887), .A2(n814), .ZN(n971) );
  NAND2_X1 U912 ( .A1(n815), .A2(n971), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(n821), .A2(G2106), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U919 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U922 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G57), .ZN(G237) );
  NOR2_X1 U927 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n828), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XOR2_X1 U930 ( .A(G2100), .B(KEYINPUT107), .Z(n830) );
  XNOR2_X1 U931 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U933 ( .A(KEYINPUT42), .B(G2090), .Z(n832) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2072), .ZN(n831) );
  XNOR2_X1 U935 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U936 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U937 ( .A(G2678), .B(G2096), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n838) );
  XOR2_X1 U939 ( .A(G2084), .B(G2078), .Z(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1956), .B(G1961), .Z(n840) );
  XNOR2_X1 U942 ( .A(G1981), .B(G1966), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U944 ( .A(n841), .B(G2474), .Z(n843) );
  XNOR2_X1 U945 ( .A(G1976), .B(G1971), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U947 ( .A(KEYINPUT41), .B(G1986), .Z(n845) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U949 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G124), .A2(n873), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n868), .A2(G100), .ZN(n849) );
  NAND2_X1 U954 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G136), .A2(n867), .ZN(n852) );
  NAND2_X1 U956 ( .A1(G112), .A2(n871), .ZN(n851) );
  NAND2_X1 U957 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U958 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n866) );
  NAND2_X1 U960 ( .A1(n873), .A2(G130), .ZN(n856) );
  NAND2_X1 U961 ( .A1(G118), .A2(n871), .ZN(n855) );
  NAND2_X1 U962 ( .A1(n856), .A2(n855), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G142), .A2(n867), .ZN(n858) );
  NAND2_X1 U964 ( .A1(G106), .A2(n868), .ZN(n857) );
  NAND2_X1 U965 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U966 ( .A(KEYINPUT109), .B(n859), .ZN(n860) );
  XNOR2_X1 U967 ( .A(KEYINPUT45), .B(n860), .ZN(n861) );
  NOR2_X1 U968 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U969 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n880) );
  NAND2_X1 U971 ( .A1(G139), .A2(n867), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G103), .A2(n868), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G115), .A2(n871), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n872), .B(KEYINPUT110), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G127), .A2(n873), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(KEYINPUT111), .B(n876), .ZN(n877) );
  XNOR2_X1 U979 ( .A(KEYINPUT47), .B(n877), .ZN(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n951) );
  XOR2_X1 U981 ( .A(n880), .B(n951), .Z(n883) );
  XOR2_X1 U982 ( .A(G160), .B(n881), .Z(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(n884), .B(n959), .Z(n886) );
  XNOR2_X1 U985 ( .A(G164), .B(G162), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n888) );
  XOR2_X1 U987 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U988 ( .A1(G37), .A2(n889), .ZN(G395) );
  XOR2_X1 U989 ( .A(KEYINPUT112), .B(G286), .Z(n891) );
  XNOR2_X1 U990 ( .A(G171), .B(n910), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U993 ( .A1(G37), .A2(n894), .ZN(G397) );
  NOR2_X1 U994 ( .A1(G227), .A2(G229), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n895), .B(KEYINPUT49), .ZN(n896) );
  NOR2_X1 U996 ( .A1(G401), .A2(n896), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G319), .A2(n897), .ZN(n898) );
  XNOR2_X1 U998 ( .A(KEYINPUT113), .B(n898), .ZN(n900) );
  NOR2_X1 U999 ( .A1(G395), .A2(G397), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U1001 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1002 ( .A(KEYINPUT56), .B(G16), .ZN(n924) );
  XOR2_X1 U1003 ( .A(G1966), .B(G168), .Z(n901) );
  NOR2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1005 ( .A(KEYINPUT57), .B(n903), .Z(n904) );
  XNOR2_X1 U1006 ( .A(KEYINPUT120), .B(n904), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(G301), .B(G1961), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n905), .B(G1341), .ZN(n906) );
  NOR2_X1 U1009 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n912) );
  XOR2_X1 U1011 ( .A(G1348), .B(n910), .Z(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n922) );
  NAND2_X1 U1013 ( .A1(G1971), .A2(G303), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(G1956), .B(G299), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n1008) );
  XNOR2_X1 U1021 ( .A(KEYINPUT115), .B(G2090), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n925), .B(G35), .ZN(n943) );
  XNOR2_X1 U1023 ( .A(G2067), .B(G26), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(G2072), .B(G33), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n936) );
  XNOR2_X1 U1026 ( .A(n928), .B(G25), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n929), .A2(G28), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(KEYINPUT116), .ZN(n934) );
  XOR2_X1 U1029 ( .A(n931), .B(G32), .Z(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT117), .B(n932), .ZN(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1033 ( .A(G27), .B(n937), .Z(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1035 ( .A(n940), .B(KEYINPUT118), .Z(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT53), .B(n941), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G34), .B(G2084), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(KEYINPUT54), .B(n944), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1041 ( .A(KEYINPUT119), .B(n947), .Z(n948) );
  NOR2_X1 U1042 ( .A1(G29), .A2(n948), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT55), .B(n949), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(G11), .ZN(n1006) );
  XOR2_X1 U1045 ( .A(G2072), .B(n951), .Z(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT114), .B(n952), .ZN(n954) );
  XOR2_X1 U1047 ( .A(G164), .B(G2078), .Z(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT50), .B(n955), .ZN(n968) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n958), .Z(n962) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G160), .B(G2084), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n972) );
  NAND2_X1 U1060 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(n973), .B(KEYINPUT52), .ZN(n974) );
  NAND2_X1 U1062 ( .A1(n974), .A2(G29), .ZN(n1004) );
  XNOR2_X1 U1063 ( .A(G1961), .B(G5), .ZN(n990) );
  XOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .Z(n975) );
  XNOR2_X1 U1065 ( .A(G4), .B(n975), .ZN(n984) );
  XOR2_X1 U1066 ( .A(G1341), .B(G19), .Z(n978) );
  XOR2_X1 U1067 ( .A(G20), .B(KEYINPUT122), .Z(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(G1956), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1070 ( .A(KEYINPUT123), .B(G1981), .Z(n979) );
  XNOR2_X1 U1071 ( .A(G6), .B(n979), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1073 ( .A(KEYINPUT124), .B(n982), .Z(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1075 ( .A(KEYINPUT60), .B(n985), .Z(n987) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G21), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(KEYINPUT125), .B(n988), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1080 ( .A(KEYINPUT126), .B(n991), .Z(n999) );
  XNOR2_X1 U1081 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n997) );
  XOR2_X1 U1082 ( .A(G1986), .B(G24), .Z(n995) );
  XNOR2_X1 U1083 ( .A(G1976), .B(G23), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G1971), .B(G22), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(n997), .B(n996), .Z(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(n1000), .B(KEYINPUT61), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G16), .B(KEYINPUT121), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(KEYINPUT62), .B(n1009), .Z(G311) );
  INV_X1 U1096 ( .A(G311), .ZN(G150) );
endmodule

