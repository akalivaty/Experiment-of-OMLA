//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n221), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  OAI211_X1 g0051(.A(G1), .B(G13), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G222), .A3(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT65), .Z(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n254), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n261), .A2(G223), .B1(G77), .B2(new_n260), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n252), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n251), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n252), .A2(G274), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n252), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G226), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OR2_X1    g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G169), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n216), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n217), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n217), .B1(new_n201), .B2(new_n202), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n267), .A2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G50), .ZN(new_n287));
  XOR2_X1   g0087(.A(new_n287), .B(KEYINPUT66), .Z(new_n288));
  INV_X1    g0088(.A(new_n276), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n285), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n284), .B1(G50), .B2(new_n285), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n263), .A2(new_n271), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n274), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n272), .A2(G200), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(G190), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n291), .B(KEYINPUT9), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n297), .A2(new_n302), .A3(new_n298), .A4(new_n299), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n296), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT70), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT68), .ZN(new_n306));
  XOR2_X1   g0106(.A(KEYINPUT8), .B(G58), .Z(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n280), .B1(G20), .B2(G77), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT15), .B(G87), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(new_n278), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n289), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n286), .A2(G77), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n290), .A2(new_n313), .B1(G77), .B2(new_n285), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n306), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n277), .A2(new_n281), .B1(new_n217), .B2(new_n203), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n276), .B1(new_n316), .B2(new_n310), .ZN(new_n317));
  INV_X1    g0117(.A(new_n285), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n276), .ZN(new_n319));
  INV_X1    g0119(.A(new_n313), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n319), .A2(new_n320), .B1(new_n203), .B2(new_n318), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(KEYINPUT68), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G244), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n266), .B1(new_n269), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n261), .A2(G238), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT67), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n254), .A2(G232), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n260), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n260), .A2(G107), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n253), .A2(KEYINPUT67), .A3(G232), .A4(new_n254), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n326), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(G169), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n305), .B1(new_n323), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n293), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n315), .A2(new_n322), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(KEYINPUT70), .C1(G169), .C2(new_n334), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT69), .ZN(new_n341));
  INV_X1    g0141(.A(G200), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n323), .B(new_n341), .C1(new_n342), .C2(new_n334), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n334), .A2(new_n342), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT69), .B1(new_n344), .B2(new_n338), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n334), .A2(G190), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n304), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G58), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n221), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n350), .B2(new_n201), .ZN(new_n351));
  INV_X1    g0151(.A(G159), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n281), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n253), .B2(G20), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n353), .B1(new_n357), .B2(G68), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n289), .B1(new_n358), .B2(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT74), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n258), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n257), .A2(KEYINPUT74), .A3(G33), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n259), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n354), .A2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n221), .B1(new_n366), .B2(new_n355), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n360), .B1(new_n367), .B2(new_n353), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(G223), .A2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n270), .A2(G1698), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n253), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n252), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n266), .B1(new_n269), .B2(new_n233), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n375), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n373), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n333), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(G200), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n307), .A2(new_n286), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n383), .A2(new_n290), .B1(new_n285), .B2(new_n307), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n369), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n369), .A2(new_n385), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n374), .A2(new_n375), .A3(new_n293), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(G169), .B2(new_n381), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT18), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(KEYINPUT18), .A3(new_n392), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(KEYINPUT75), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n384), .B1(new_n359), .B2(new_n368), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n396), .A2(new_n397), .A3(new_n391), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT75), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n388), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(KEYINPUT76), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n233), .A2(G1698), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n253), .B(new_n404), .C1(G226), .C2(G1698), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n252), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n266), .B1(new_n269), .B2(new_n222), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT13), .B1(new_n407), .B2(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n403), .B1(new_n413), .B2(G169), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n413), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G179), .ZN(new_n417));
  INV_X1    g0217(.A(new_n412), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n407), .A2(KEYINPUT13), .A3(new_n408), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n403), .B(G169), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n415), .A2(KEYINPUT73), .A3(new_n417), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT73), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n420), .B1(new_n293), .B2(new_n413), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n414), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n319), .A2(G68), .A3(new_n286), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n318), .A2(new_n221), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT12), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(KEYINPUT71), .A3(new_n428), .ZN(new_n429));
  XOR2_X1   g0229(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n430));
  OAI211_X1 g0230(.A(new_n426), .B(new_n429), .C1(new_n427), .C2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(KEYINPUT72), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(KEYINPUT72), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n281), .A2(new_n202), .B1(new_n217), .B2(G68), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n278), .A2(new_n203), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n276), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT11), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n425), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n416), .B2(G190), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n413), .A2(G200), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n394), .A2(KEYINPUT75), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n397), .B1(new_n396), .B2(new_n391), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n400), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n386), .B(KEYINPUT17), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n446), .A2(KEYINPUT76), .A3(new_n447), .ZN(new_n448));
  NOR4_X1   g0248(.A1(new_n348), .A2(new_n402), .A3(new_n443), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(G97), .B(G107), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI22_X1  g0254(.A1(new_n454), .A2(new_n217), .B1(new_n203), .B2(new_n281), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n207), .B1(new_n366), .B2(new_n355), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n276), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n267), .A2(G33), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n289), .A2(new_n285), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n318), .A2(new_n206), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n264), .A2(G1), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT5), .B(G41), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n333), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G257), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n467), .A2(new_n252), .A3(G274), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n253), .A2(G244), .A3(new_n254), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G250), .A2(G1698), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT4), .A2(G244), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(G1698), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n253), .A2(new_n477), .B1(G33), .B2(G283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n252), .B1(new_n479), .B2(KEYINPUT77), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT77), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n474), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  AOI211_X1 g0282(.A(G190), .B(new_n471), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(KEYINPUT77), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n333), .A3(new_n482), .ZN(new_n485));
  INV_X1    g0285(.A(new_n471), .ZN(new_n486));
  AOI21_X1  g0286(.A(G200), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n465), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n293), .A3(new_n486), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n471), .B1(new_n480), .B2(new_n482), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n464), .C1(G169), .C2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n309), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n285), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n253), .A2(new_n217), .A3(G68), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT19), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n217), .B1(new_n406), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G87), .B2(new_n208), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n278), .B2(new_n206), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  OR2_X1    g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n289), .B1(new_n499), .B2(new_n500), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n493), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n460), .A2(new_n492), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n252), .B(G250), .C1(G1), .C2(new_n264), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n252), .A2(G274), .A3(new_n466), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT78), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n254), .A2(G238), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n260), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n253), .A2(KEYINPUT78), .A3(G238), .A4(new_n254), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n253), .A2(G244), .A3(G1698), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n508), .B1(new_n515), .B2(new_n333), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n273), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n293), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n505), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n459), .A2(new_n223), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n493), .B(new_n521), .C1(new_n501), .C2(new_n502), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(G200), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(G190), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n488), .A2(new_n491), .A3(new_n520), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT25), .B1(new_n318), .B2(new_n207), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n318), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n460), .A2(G107), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n258), .A2(new_n259), .A3(new_n217), .A4(G87), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT22), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n217), .A3(G87), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n260), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n223), .A2(KEYINPUT22), .A3(G20), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT81), .B1(new_n253), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n534), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT82), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n535), .B1(new_n260), .B2(new_n537), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n253), .A2(KEYINPUT81), .A3(new_n539), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT82), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n534), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n513), .A2(G20), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT23), .B1(new_n207), .B2(G20), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n532), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n553), .ZN(new_n555));
  AOI211_X1 g0355(.A(KEYINPUT24), .B(new_n555), .C1(new_n542), .C2(new_n547), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n276), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT83), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI221_X4 g0359(.A(KEYINPUT82), .B1(new_n533), .B2(KEYINPUT22), .C1(new_n543), .C2(new_n544), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n546), .B1(new_n545), .B2(new_n534), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n553), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT24), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n548), .A2(new_n532), .A3(new_n553), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(KEYINPUT83), .A3(new_n276), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n531), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT84), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n254), .A2(G250), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n260), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n253), .A2(KEYINPUT84), .A3(G250), .A4(new_n254), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n253), .A2(G257), .A3(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n333), .B1(G264), .B2(new_n468), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n470), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n342), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G190), .B2(new_n576), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n526), .B1(new_n567), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n319), .A2(G116), .A3(new_n458), .ZN(new_n581));
  INV_X1    g0381(.A(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n318), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n275), .A2(new_n216), .B1(G20), .B2(new_n582), .ZN(new_n584));
  AOI21_X1  g0384(.A(G20), .B1(G33), .B2(G283), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G33), .B2(new_n206), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n584), .A2(new_n586), .A3(KEYINPUT20), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT20), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n581), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G169), .ZN(new_n590));
  NAND2_X1  g0390(.A1(KEYINPUT5), .A2(G41), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT5), .A2(G41), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n466), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(G270), .A3(new_n252), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n470), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n258), .A2(new_n259), .A3(G257), .A4(new_n254), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n258), .A2(new_n259), .A3(G264), .A4(G1698), .ZN(new_n598));
  INV_X1    g0398(.A(G303), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n253), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n596), .B1(new_n333), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n580), .B1(new_n590), .B2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n595), .A2(new_n470), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n333), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(G190), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n587), .A2(new_n588), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n583), .B1(new_n459), .B2(new_n582), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n605), .B(new_n608), .C1(new_n601), .C2(new_n342), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n601), .A2(G179), .A3(new_n589), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n604), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n611), .A2(KEYINPUT21), .A3(new_n589), .A4(G169), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n602), .A2(new_n609), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT80), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT83), .B1(new_n565), .B2(new_n276), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n558), .B(new_n289), .C1(new_n563), .C2(new_n564), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n530), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n576), .A2(G179), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n273), .B2(new_n576), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n615), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n449), .A2(new_n579), .A3(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n301), .A2(new_n303), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n339), .A2(new_n337), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n442), .A2(new_n336), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n388), .B1(new_n439), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n393), .B2(new_n398), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n394), .A2(KEYINPUT85), .A3(new_n445), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n623), .B1(new_n626), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n295), .ZN(new_n633));
  INV_X1    g0433(.A(new_n449), .ZN(new_n634));
  INV_X1    g0434(.A(new_n491), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(KEYINPUT26), .A3(new_n520), .A4(new_n525), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n520), .A2(new_n525), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(new_n491), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n518), .A2(new_n519), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n636), .A2(new_n639), .B1(new_n505), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n602), .A2(new_n610), .A3(new_n612), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n618), .B2(new_n620), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n530), .B(new_n578), .C1(new_n616), .C2(new_n617), .ZN(new_n645));
  INV_X1    g0445(.A(new_n526), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n642), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n633), .B1(new_n634), .B2(new_n649), .ZN(G369));
  NAND3_X1  g0450(.A1(new_n267), .A2(new_n217), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n618), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n657), .A2(new_n645), .B1(new_n618), .B2(new_n620), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n618), .A2(new_n620), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n656), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n613), .B(KEYINPUT80), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n589), .A2(new_n656), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT86), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n643), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n661), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n656), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n645), .B1(new_n567), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n659), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n666), .A2(new_n656), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n660), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n211), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n214), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n648), .A2(new_n685), .A3(new_n672), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n648), .B2(new_n672), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n621), .A2(new_n579), .A3(new_n672), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n485), .A2(new_n486), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n575), .A2(new_n516), .A3(new_n601), .A4(G179), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n516), .A2(new_n601), .A3(G179), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n691), .A3(new_n576), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n575), .A2(new_n516), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n611), .A2(new_n293), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n490), .A3(KEYINPUT30), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT87), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT87), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n693), .A2(new_n695), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n656), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n672), .A2(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n703), .A2(new_n704), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n688), .B1(new_n689), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n686), .A2(new_n687), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n684), .B1(new_n708), .B2(G1), .ZN(G364));
  AND2_X1   g0509(.A1(new_n217), .A2(G13), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n267), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n679), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(G355), .A2(new_n253), .A3(new_n211), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n248), .A2(new_n264), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n678), .A2(new_n253), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(G45), .B2(new_n214), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n715), .B1(G116), .B2(new_n211), .C1(new_n716), .C2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n216), .B1(G20), .B2(new_n273), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n714), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n723), .ZN(new_n726));
  NAND2_X1  g0526(.A1(G20), .A2(G179), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT88), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n376), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G311), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n729), .A2(new_n342), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(KEYINPUT33), .B(G317), .Z(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(G20), .A3(new_n376), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n253), .B1(new_n738), .B2(G329), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n217), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(new_n376), .A3(G200), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT89), .Z(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G283), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n739), .B1(new_n599), .B2(new_n741), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n728), .A2(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n735), .B(new_n746), .C1(G322), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n342), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n736), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n750), .A2(G326), .B1(G294), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT90), .Z(new_n754));
  NOR2_X1   g0554(.A1(new_n733), .A2(new_n221), .ZN(new_n755));
  INV_X1    g0555(.A(new_n730), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n203), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n755), .B(new_n757), .C1(G107), .C2(new_n743), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G50), .A2(new_n750), .B1(new_n748), .B2(G58), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n737), .A2(new_n352), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n741), .A2(new_n223), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n260), .B(new_n762), .C1(G97), .C2(new_n752), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n749), .A2(new_n754), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n722), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n725), .B1(new_n726), .B2(new_n765), .C1(new_n668), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n669), .A2(new_n714), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n668), .A2(G330), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(G396));
  NAND2_X1  g0570(.A1(new_n648), .A2(new_n672), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n323), .A2(new_n672), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n347), .A2(new_n340), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT92), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n624), .A2(new_n775), .A3(new_n336), .A4(new_n772), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n336), .A2(new_n337), .A3(new_n772), .A4(new_n339), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(KEYINPUT92), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n774), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT93), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n774), .A2(new_n776), .A3(new_n778), .A4(KEYINPUT93), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n771), .B(new_n783), .Z(new_n784));
  INV_X1    g0584(.A(new_n707), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n713), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n744), .A2(new_n223), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G311), .B2(new_n738), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT91), .Z(new_n790));
  INV_X1    g0590(.A(new_n752), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n260), .B1(new_n741), .B2(new_n207), .C1(new_n791), .C2(new_n206), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(G303), .B2(new_n750), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n582), .A2(new_n756), .B1(new_n733), .B2(new_n745), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G294), .B2(new_n748), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n790), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G137), .A2(new_n750), .B1(new_n732), .B2(G150), .ZN(new_n797));
  INV_X1    g0597(.A(G143), .ZN(new_n798));
  INV_X1    g0598(.A(new_n748), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(new_n798), .B2(new_n799), .C1(new_n352), .C2(new_n756), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT34), .ZN(new_n801));
  INV_X1    g0601(.A(G132), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n253), .B1(new_n737), .B2(new_n802), .C1(new_n741), .C2(new_n202), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n744), .A2(new_n221), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(G58), .C2(new_n752), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n726), .B1(new_n796), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n723), .A2(new_n720), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n714), .B(new_n807), .C1(new_n203), .C2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n721), .B2(new_n783), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n787), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G384));
  INV_X1    g0612(.A(new_n454), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(KEYINPUT35), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(KEYINPUT35), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n814), .A2(G116), .A3(new_n218), .A4(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT36), .Z(new_n817));
  OAI211_X1 g0617(.A(new_n215), .B(G77), .C1(new_n349), .C2(new_n221), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n267), .B(G13), .C1(new_n818), .C2(new_n244), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT38), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT94), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n358), .A2(KEYINPUT16), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n221), .B1(new_n355), .B2(new_n356), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n360), .B1(new_n824), .B2(new_n353), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n823), .A2(new_n276), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n385), .ZN(new_n827));
  INV_X1    g0627(.A(new_n654), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(KEYINPUT94), .B(new_n654), .C1(new_n826), .C2(new_n385), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n446), .B2(new_n447), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n386), .B1(new_n396), .B2(new_n391), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n396), .A2(new_n654), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n833), .A2(KEYINPUT37), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n827), .A2(new_n828), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(KEYINPUT94), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n827), .A2(new_n822), .A3(new_n828), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n827), .A2(new_n392), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n837), .A2(new_n386), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n835), .B1(KEYINPUT37), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n821), .B1(new_n832), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n834), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n389), .A2(new_n392), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n386), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n839), .A2(new_n386), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n847), .A2(new_n829), .A3(new_n830), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n846), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n849), .B(KEYINPUT38), .C1(new_n401), .C2(new_n831), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n842), .A2(new_n850), .A3(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n843), .B1(new_n630), .B2(new_n447), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n833), .B2(new_n834), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(new_n846), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n821), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT39), .B1(new_n855), .B2(new_n850), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n439), .A2(new_n656), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n438), .A2(new_n656), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n439), .A2(new_n442), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n442), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n438), .B(new_n656), .C1(new_n425), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n783), .A2(new_n648), .A3(new_n672), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n340), .A2(new_n656), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n842), .A2(new_n850), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n631), .A2(new_n654), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n859), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n449), .B1(new_n686), .B2(new_n687), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n633), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n874), .B(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n855), .A2(new_n850), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n700), .A2(new_n705), .A3(new_n702), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n704), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n689), .B(new_n879), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n862), .A2(new_n864), .B1(new_n781), .B2(new_n782), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n878), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT40), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT40), .B1(new_n842), .B2(new_n850), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n883), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n449), .A2(new_n883), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n891), .A2(new_n892), .A3(new_n688), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n877), .A2(new_n893), .B1(new_n267), .B2(new_n710), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n877), .A2(new_n893), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n820), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n896), .B(KEYINPUT96), .Z(G367));
  INV_X1    g0697(.A(new_n750), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n202), .A2(new_n756), .B1(new_n898), .B2(new_n798), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n791), .A2(new_n221), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n260), .B1(new_n738), .B2(G137), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n349), .B2(new_n741), .ZN(new_n902));
  INV_X1    g0702(.A(new_n742), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n900), .B(new_n902), .C1(G77), .C2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n279), .B2(new_n799), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n899), .B(new_n905), .C1(G159), .C2(new_n732), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT103), .ZN(new_n907));
  AOI22_X1  g0707(.A1(G303), .A2(new_n748), .B1(new_n750), .B2(G311), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT102), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(KEYINPUT102), .ZN(new_n910));
  INV_X1    g0710(.A(G317), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n260), .B1(new_n911), .B2(new_n737), .C1(new_n791), .C2(new_n207), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(G97), .B2(new_n903), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n741), .A2(new_n582), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT46), .Z(new_n915));
  AOI22_X1  g0715(.A1(G283), .A2(new_n730), .B1(new_n732), .B2(G294), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n910), .A2(new_n913), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n907), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT47), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n723), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n522), .A2(new_n672), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n638), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n641), .A2(new_n921), .A3(new_n505), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n722), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n239), .A2(new_n717), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n723), .B(new_n722), .C1(new_n678), .C2(new_n492), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n714), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n920), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n620), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n567), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n672), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n675), .B1(new_n674), .B2(new_n931), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n673), .A2(new_n930), .A3(new_n666), .A4(new_n656), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n670), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n675), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n658), .B2(new_n660), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n559), .A2(new_n566), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n672), .B1(new_n937), .B2(new_n530), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n576), .A2(G190), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n342), .B2(new_n576), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n531), .B(new_n940), .C1(new_n559), .C2(new_n566), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n942), .A2(new_n643), .A3(new_n659), .A4(new_n672), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n936), .A2(new_n669), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n708), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n671), .A2(KEYINPUT100), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n464), .A2(new_n656), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n488), .A2(new_n491), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT97), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n488), .A2(KEYINPUT97), .A3(new_n491), .A4(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n635), .A2(new_n656), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n931), .B(new_n954), .C1(new_n658), .C2(new_n935), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n943), .A2(KEYINPUT45), .A3(new_n931), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT99), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n676), .B2(new_n954), .ZN(new_n962));
  INV_X1    g0762(.A(new_n954), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n933), .C2(new_n660), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n959), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n946), .B1(new_n947), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n671), .A2(KEYINPUT100), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n968), .A2(new_n959), .A3(new_n962), .A4(new_n965), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT101), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n957), .A2(new_n958), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n962), .A2(new_n965), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n947), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n945), .A2(new_n708), .ZN(new_n974));
  AND4_X1   g0774(.A1(KEYINPUT101), .A2(new_n973), .A3(new_n969), .A4(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n708), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n679), .B(new_n977), .Z(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n712), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n933), .A2(new_n954), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT42), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n951), .A2(new_n952), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n491), .B1(new_n983), .B2(new_n659), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n981), .A2(KEYINPUT42), .B1(new_n672), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n922), .A2(new_n923), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n982), .A2(new_n985), .B1(KEYINPUT43), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n671), .A2(new_n963), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n990), .B1(new_n989), .B2(new_n991), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n928), .B1(new_n980), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT104), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n928), .ZN(new_n999));
  INV_X1    g0799(.A(new_n708), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n973), .A2(new_n969), .A3(new_n974), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT101), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT101), .A4(new_n969), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n711), .B1(new_n1005), .B2(new_n978), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n999), .B1(new_n1006), .B2(new_n994), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT104), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n998), .A2(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n945), .A2(new_n712), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n253), .B1(new_n737), .B2(new_n279), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n791), .A2(new_n309), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n741), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1012), .C1(G77), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n748), .A2(G50), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n743), .A2(G97), .B1(new_n732), .B2(new_n307), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G68), .A2(new_n730), .B1(new_n750), .B2(G159), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n253), .B1(new_n738), .B2(G326), .ZN(new_n1019));
  INV_X1    g0819(.A(G294), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n791), .A2(new_n745), .B1(new_n741), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G311), .A2(new_n732), .B1(new_n750), .B2(G322), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n599), .B2(new_n756), .C1(new_n911), .C2(new_n799), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1019), .B1(new_n582), .B2(new_n742), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1018), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n723), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n236), .A2(G45), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT105), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n307), .A2(new_n202), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n681), .B(new_n264), .C1(new_n221), .C2(new_n203), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n717), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n253), .A2(new_n211), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(G107), .B2(new_n211), .C1(new_n681), .C2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n714), .B1(new_n1039), .B2(new_n724), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1031), .B(new_n1040), .C1(new_n661), .C2(new_n766), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n946), .A2(new_n679), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n945), .A2(new_n708), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1010), .B(new_n1041), .C1(new_n1042), .C2(new_n1043), .ZN(G393));
  INV_X1    g0844(.A(new_n671), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n971), .B2(new_n972), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n959), .A2(new_n671), .A3(new_n962), .A4(new_n965), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n680), .B1(new_n1048), .B2(new_n946), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n970), .B2(new_n975), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n717), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n724), .B1(new_n206), .B2(new_n211), .C1(new_n243), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n713), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n791), .A2(new_n203), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n260), .B(new_n1054), .C1(G143), .C2(new_n738), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n221), .B2(new_n741), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n202), .A2(new_n733), .B1(new_n756), .B2(new_n277), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n788), .B(new_n1056), .C1(KEYINPUT106), .C2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G150), .A2(new_n750), .B1(new_n748), .B2(G159), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT51), .Z(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(KEYINPUT106), .C2(new_n1057), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT107), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G311), .A2(new_n748), .B1(new_n750), .B2(G317), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  AOI22_X1  g0865(.A1(new_n732), .A2(G303), .B1(G116), .B2(new_n752), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1020), .B2(new_n756), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n253), .B1(new_n738), .B2(G322), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n745), .B2(new_n741), .C1(new_n744), .C2(new_n207), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT108), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1065), .B(new_n1071), .C1(new_n1070), .C2(new_n1069), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1063), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1053), .B1(new_n1074), .B2(new_n723), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n963), .A2(new_n722), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1048), .B2(new_n711), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1050), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT109), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1050), .A2(KEYINPUT109), .A3(new_n1079), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(new_n808), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n732), .A2(G137), .ZN(new_n1086));
  INV_X1    g0886(.A(G128), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n898), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(G125), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n253), .B1(new_n737), .B2(new_n1089), .C1(new_n742), .C2(new_n202), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G159), .B2(new_n752), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n802), .B2(new_n799), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(KEYINPUT54), .B(G143), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT111), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1088), .B(new_n1092), .C1(new_n730), .C2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n741), .A2(new_n279), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT112), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT53), .Z(new_n1098));
  OAI21_X1  g0898(.A(new_n260), .B1(new_n737), .B2(new_n1020), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n804), .A2(new_n762), .A3(new_n1054), .A4(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n206), .A2(new_n756), .B1(new_n733), .B2(new_n207), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n582), .A2(new_n799), .B1(new_n898), .B2(new_n745), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1095), .A2(new_n1098), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n713), .B1(new_n307), .B2(new_n1085), .C1(new_n1104), .C2(new_n726), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT39), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n878), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n842), .A2(new_n850), .A3(KEYINPUT39), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1105), .B1(new_n1109), .B2(new_n720), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n707), .A2(new_n783), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n865), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n867), .A2(new_n869), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n865), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n858), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1109), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n870), .A2(new_n858), .A3(new_n878), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n878), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n857), .B1(new_n870), .B2(new_n858), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n883), .A2(new_n884), .A3(G330), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1111), .B1(new_n1125), .B2(new_n711), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1121), .A2(new_n1122), .B1(new_n865), .B2(new_n1112), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n449), .A2(G330), .A3(new_n883), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n875), .A2(new_n1131), .A3(new_n633), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n883), .A2(G330), .A3(new_n783), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n866), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT110), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1114), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(KEYINPUT110), .A3(new_n866), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1113), .A4(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n865), .B1(new_n707), .B2(new_n783), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1114), .B1(new_n1123), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1132), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n679), .B1(new_n1130), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1113), .A3(new_n1137), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT110), .B1(new_n1133), .B2(new_n866), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1132), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1125), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1127), .B1(new_n1143), .B2(new_n1149), .ZN(G378));
  NAND3_X1  g0950(.A1(new_n859), .A2(new_n872), .A3(new_n873), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n291), .A2(new_n828), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n304), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n304), .A2(new_n1152), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n889), .B2(G330), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n688), .B(new_n1158), .C1(new_n886), .C2(new_n888), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1151), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n883), .A2(new_n884), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n887), .B1(new_n885), .B2(KEYINPUT40), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1158), .B1(new_n1164), .B2(new_n688), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n889), .A2(G330), .A3(new_n1159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n874), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1158), .A2(new_n720), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n713), .B1(new_n1085), .B2(G50), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G97), .A2(new_n732), .B1(new_n730), .B2(new_n492), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT114), .Z(new_n1172));
  AOI21_X1  g0972(.A(new_n900), .B1(new_n750), .B2(G116), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT115), .Z(new_n1174));
  NOR2_X1   g0974(.A1(new_n799), .A2(new_n207), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n260), .A2(new_n251), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G283), .B2(new_n738), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n349), .B2(new_n742), .C1(new_n203), .C2(new_n741), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT116), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1176), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT113), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n1094), .A2(new_n1013), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n279), .B2(new_n791), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G128), .B2(new_n748), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G132), .A2(new_n732), .B1(new_n730), .B2(G137), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1188), .A2(KEYINPUT117), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(KEYINPUT117), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1187), .B1(new_n1089), .B2(new_n898), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n738), .C2(G124), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n352), .B2(new_n742), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1191), .B2(KEYINPUT59), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1184), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1181), .A2(new_n1182), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1170), .B1(new_n1197), .B2(new_n723), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1168), .A2(new_n712), .B1(new_n1169), .B2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1160), .A2(new_n1161), .A3(new_n1151), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n874), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1132), .B(KEYINPUT118), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1130), .B2(new_n1142), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n679), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1203), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1148), .B2(new_n1125), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1168), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1199), .B1(new_n1205), .B2(new_n1208), .ZN(G375));
  NAND3_X1  g1009(.A1(new_n1139), .A2(new_n1141), .A3(new_n1132), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1148), .A2(new_n979), .A3(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT119), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1146), .A2(new_n712), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n713), .B1(new_n1085), .B2(G68), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n253), .B(new_n1012), .C1(G303), .C2(new_n738), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n206), .B2(new_n741), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G283), .B2(new_n748), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n203), .B2(new_n744), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G116), .A2(new_n732), .B1(new_n750), .B2(G294), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n207), .B2(new_n756), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT120), .Z(new_n1221));
  AOI21_X1  g1021(.A(new_n260), .B1(new_n903), .B2(G58), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n748), .A2(G137), .B1(new_n1222), .B2(KEYINPUT122), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n732), .A2(new_n1094), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(KEYINPUT122), .C2(new_n1222), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n898), .B2(new_n802), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n750), .A2(KEYINPUT121), .A3(G132), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n730), .A2(G150), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n741), .A2(new_n352), .B1(new_n1087), .B2(new_n737), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G50), .B2(new_n752), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1218), .A2(new_n1221), .B1(new_n1225), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1214), .B1(new_n1233), .B2(new_n723), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n865), .B2(new_n721), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1213), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1212), .A2(new_n1237), .ZN(G381));
  NOR4_X1   g1038(.A1(G378), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1081), .B(new_n1078), .C1(new_n1240), .C2(new_n1049), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT109), .B1(new_n1050), .B2(new_n1079), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  OR4_X1    g1044(.A1(G387), .A2(new_n1244), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1045(.A(new_n1143), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1149), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1126), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n655), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G375), .C2(new_n1249), .ZN(G409));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1146), .A2(new_n1251), .A3(new_n1147), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(new_n680), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1210), .B1(new_n1142), .B2(new_n1251), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1236), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(G384), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(G384), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n655), .A2(G213), .ZN(new_n1259));
  INV_X1    g1059(.A(G2897), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1258), .A3(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1255), .A2(G384), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n1263), .A2(new_n1256), .B1(new_n1260), .B2(new_n1259), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1199), .C1(new_n1205), .C2(new_n1208), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1207), .A2(new_n979), .A3(new_n1168), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1199), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1248), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1259), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT61), .B1(new_n1265), .B2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1263), .A2(new_n1256), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1273), .A3(new_n1259), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT123), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1270), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1266), .A2(new_n1269), .A3(KEYINPUT123), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(new_n1273), .A3(new_n1278), .A4(new_n1259), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1272), .B(new_n1275), .C1(new_n1279), .C2(KEYINPUT62), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(G393), .B(G396), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n996), .A2(new_n1243), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(G390), .A2(new_n1007), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT125), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n996), .A2(new_n1243), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1006), .A2(new_n994), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1288), .B(new_n928), .C1(new_n1242), .C2(new_n1241), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1282), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n998), .A2(new_n1008), .A3(new_n1243), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(new_n1281), .A3(new_n1289), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT126), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1291), .B1(new_n1290), .B2(new_n1282), .ZN(new_n1297));
  AOI211_X1 g1097(.A(KEYINPUT125), .B(new_n1281), .C1(new_n1287), .C2(new_n1289), .ZN(new_n1298));
  OAI211_X1 g1098(.A(KEYINPUT126), .B(new_n1295), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1280), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1274), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1279), .A2(KEYINPUT124), .A3(new_n1303), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1279), .A2(new_n1303), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT124), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1277), .A2(new_n1278), .A3(new_n1259), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1265), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1305), .A2(new_n1306), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1301), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1273), .A2(KEYINPUT127), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G375), .A2(new_n1248), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1266), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1315), .B(new_n1317), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1314), .B(new_n1318), .ZN(G402));
endmodule


