//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906;
  XOR2_X1   g000(.A(KEYINPUT66), .B(G190gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT28), .Z(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  OR3_X1    g005(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(new_n206), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n202), .A2(KEYINPUT67), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n206), .B(KEYINPUT24), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G190gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G183gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  OAI22_X1  g022(.A1(new_n222), .A2(new_n223), .B1(new_n209), .B2(new_n210), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n220), .A2(KEYINPUT68), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT68), .B1(new_n220), .B2(new_n226), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n216), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n224), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n227), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n213), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G226gat), .A2(G233gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(KEYINPUT74), .A3(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n235), .B(KEYINPUT73), .Z(new_n238));
  NOR2_X1   g037(.A1(new_n213), .A2(new_n233), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(KEYINPUT29), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT74), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n239), .B2(new_n235), .ZN(new_n242));
  XNOR2_X1  g041(.A(G197gat), .B(G204gat), .ZN(new_n243));
  INV_X1    g042(.A(G211gat), .ZN(new_n244));
  INV_X1    g043(.A(G218gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n243), .B1(KEYINPUT22), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n237), .A2(new_n240), .A3(new_n242), .A4(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n252), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n236), .B1(new_n234), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n239), .A2(new_n238), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n249), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT38), .B1(new_n259), .B2(KEYINPUT37), .ZN(new_n260));
  XNOR2_X1  g059(.A(G8gat), .B(G36gat), .ZN(new_n261));
  INV_X1    g060(.A(G64gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G92gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n237), .A2(new_n240), .A3(new_n242), .A4(new_n249), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT37), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI211_X1 g070(.A(KEYINPUT85), .B(KEYINPUT37), .C1(new_n267), .C2(new_n268), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n260), .B(new_n265), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n265), .B1(new_n271), .B2(new_n272), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n269), .A2(new_n270), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT38), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G134gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n280), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n286));
  INV_X1    g085(.A(G127gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G134gat), .ZN(new_n288));
  OAI221_X1 g087(.A(new_n286), .B1(KEYINPUT69), .B2(new_n288), .C1(KEYINPUT1), .C2(new_n279), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291));
  INV_X1    g090(.A(G155gat), .ZN(new_n292));
  INV_X1    g091(.A(G162gat), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT2), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G155gat), .B(G162gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  OR3_X1    g096(.A1(new_n290), .A2(new_n297), .A3(KEYINPUT4), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n290), .ZN(new_n301));
  INV_X1    g100(.A(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT4), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(new_n299), .A3(new_n298), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(new_n290), .ZN(new_n308));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n300), .A2(new_n305), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n290), .B(new_n297), .ZN(new_n312));
  INV_X1    g111(.A(new_n309), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n304), .A2(new_n298), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n316), .A2(new_n311), .A3(new_n308), .A4(new_n309), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT0), .B(G57gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(G85gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT6), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n315), .A2(new_n322), .A3(new_n317), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n327), .A2(new_n325), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n273), .A2(new_n276), .A3(new_n278), .A4(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G78gat), .B(G106gat), .Z(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT31), .ZN(new_n332));
  INV_X1    g131(.A(G50gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n249), .A2(KEYINPUT29), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT3), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT79), .B1(new_n249), .B2(KEYINPUT29), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n302), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n250), .B1(new_n306), .B2(new_n255), .ZN(new_n341));
  INV_X1    g140(.A(G228gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n340), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n341), .ZN(new_n345));
  AOI211_X1 g144(.A(new_n342), .B(new_n343), .C1(new_n336), .C2(new_n297), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n307), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G22gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n335), .B1(new_n349), .B2(KEYINPUT78), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(G22gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT80), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n348), .A2(G22gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n352), .A2(new_n353), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n335), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n316), .A2(new_n308), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n313), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT82), .B1(new_n312), .B2(new_n313), .ZN(new_n364));
  OR3_X1    g163(.A1(new_n312), .A2(KEYINPUT82), .A3(new_n313), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n363), .A2(KEYINPUT39), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT81), .B(KEYINPUT39), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n366), .B(new_n322), .C1(new_n363), .C2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT40), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n368), .A2(KEYINPUT83), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT83), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n368), .A2(new_n369), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n265), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT30), .B1(new_n269), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(new_n277), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n277), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n373), .A2(new_n377), .A3(new_n324), .A4(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n330), .A2(new_n361), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT86), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT71), .B(G71gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(G99gat), .ZN(new_n383));
  XOR2_X1   g182(.A(G15gat), .B(G43gat), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386));
  XOR2_X1   g185(.A(new_n386), .B(KEYINPUT64), .Z(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n234), .A2(new_n290), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n239), .A2(new_n301), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n385), .B1(new_n391), .B2(KEYINPUT33), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n388), .A3(new_n390), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT34), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n392), .A2(new_n394), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n398), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n392), .A2(new_n394), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n395), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT36), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n400), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT72), .B1(new_n402), .B2(new_n395), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n398), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT72), .B(new_n401), .C1(new_n402), .C2(new_n395), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n405), .B1(new_n409), .B2(KEYINPUT36), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n327), .A2(KEYINPUT76), .A3(new_n325), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n324), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT76), .B1(new_n327), .B2(new_n325), .ZN(new_n413));
  OAI22_X1  g212(.A1(new_n412), .A2(new_n413), .B1(new_n325), .B2(new_n324), .ZN(new_n414));
  INV_X1    g213(.A(new_n378), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n376), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT77), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n377), .A2(new_n378), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT77), .A3(new_n414), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n410), .B1(new_n421), .B2(new_n360), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n330), .A2(new_n423), .A3(new_n361), .A4(new_n379), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n381), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n360), .B1(new_n407), .B2(new_n408), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT35), .B1(new_n427), .B2(new_n421), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n400), .A2(new_n403), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(new_n360), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT35), .ZN(new_n432));
  INV_X1    g231(.A(new_n329), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n419), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G57gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G64gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n262), .A2(G57gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G78gat), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n443), .B2(new_n440), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G85gat), .A2(G92gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT98), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(G85gat), .A3(G92gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT7), .ZN(new_n452));
  XNOR2_X1  g251(.A(G99gat), .B(G106gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454));
  INV_X1    g253(.A(G85gat), .ZN(new_n455));
  AOI22_X1  g254(.A1(KEYINPUT8), .A2(new_n454), .B1(new_n455), .B2(new_n264), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT7), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n448), .A2(KEYINPUT98), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n452), .A2(new_n453), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n452), .A2(new_n456), .A3(new_n458), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT99), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(G71gat), .A2(G78gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(G71gat), .A2(G78gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n442), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n470), .A2(new_n444), .A3(KEYINPUT94), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT94), .B1(new_n470), .B2(new_n444), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n462), .A2(new_n459), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT99), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n465), .B1(new_n475), .B2(new_n463), .ZN(new_n476));
  NAND2_X1  g275(.A1(G230gat), .A2(G233gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G120gat), .B(G148gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G204gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT103), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(new_n210), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT102), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT10), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n473), .A2(new_n485), .A3(new_n474), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n444), .A3(KEYINPUT94), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n445), .B2(new_n446), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n464), .A3(new_n463), .ZN(new_n492));
  INV_X1    g291(.A(new_n474), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT99), .A3(new_n447), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT100), .B1(new_n495), .B2(new_n485), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT100), .ZN(new_n497));
  AOI211_X1 g296(.A(new_n497), .B(KEYINPUT10), .C1(new_n492), .C2(new_n494), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n487), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT101), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT101), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n487), .C1(new_n496), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n484), .B1(new_n503), .B2(new_n477), .ZN(new_n504));
  AOI211_X1 g303(.A(KEYINPUT102), .B(new_n478), .C1(new_n500), .C2(new_n502), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n479), .B(new_n483), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT104), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n497), .B1(new_n476), .B2(KEYINPUT10), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n495), .A2(KEYINPUT100), .A3(new_n485), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n501), .B1(new_n511), .B2(new_n487), .ZN(new_n512));
  AOI211_X1 g311(.A(KEYINPUT101), .B(new_n486), .C1(new_n509), .C2(new_n510), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n477), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT102), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n503), .A2(new_n484), .A3(new_n477), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(KEYINPUT104), .A3(new_n479), .A4(new_n483), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n477), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n479), .ZN(new_n521));
  INV_X1    g320(.A(new_n483), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT16), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(G1gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G1gat), .B2(new_n525), .ZN(new_n528));
  INV_X1    g327(.A(G8gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT21), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n473), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT96), .Z(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n473), .A2(new_n531), .ZN(new_n536));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT95), .ZN(new_n540));
  XOR2_X1   g339(.A(G183gat), .B(G211gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n538), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n535), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  INV_X1    g347(.A(G36gat), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(KEYINPUT87), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n546), .B(new_n550), .C1(new_n553), .C2(KEYINPUT87), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n333), .A2(G43gat), .ZN(new_n555));
  INV_X1    g354(.A(G43gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G50gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(KEYINPUT15), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT15), .B1(new_n555), .B2(KEYINPUT88), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n558), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n555), .B(new_n557), .C1(KEYINPUT88), .C2(KEYINPUT15), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(new_n553), .A3(new_n546), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(KEYINPUT17), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT89), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n560), .A2(new_n569), .A3(new_n564), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n572));
  AOI21_X1  g371(.A(new_n566), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n560), .A2(new_n569), .A3(new_n564), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n569), .B1(new_n560), .B2(new_n564), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n566), .B(new_n572), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n565), .B(new_n474), .C1(new_n573), .C2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n571), .A2(new_n493), .B1(KEYINPUT41), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G190gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n581), .B(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT97), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G218gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n584), .B(new_n587), .Z(new_n588));
  NOR3_X1   g387(.A1(new_n524), .A2(new_n545), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n436), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n530), .A2(new_n565), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n573), .B2(new_n577), .ZN(new_n592));
  INV_X1    g391(.A(new_n571), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n593), .A2(new_n530), .ZN(new_n594));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n571), .B(new_n530), .Z(new_n599));
  XOR2_X1   g398(.A(new_n595), .B(KEYINPUT13), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n592), .A2(KEYINPUT18), .A3(new_n594), .A4(new_n595), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT11), .B(G169gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G197gat), .ZN(new_n605));
  XOR2_X1   g404(.A(G113gat), .B(G141gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n598), .A2(new_n608), .A3(new_n601), .A4(new_n602), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(KEYINPUT92), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n603), .A2(new_n613), .A3(new_n609), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT93), .B1(new_n612), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n414), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g421(.A1(new_n618), .A2(new_n419), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n526), .A2(new_n529), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n626), .A2(KEYINPUT42), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(KEYINPUT42), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n627), .B(new_n628), .C1(new_n529), .C2(new_n623), .ZN(G1325gat));
  AOI21_X1  g428(.A(G15gat), .B1(new_n619), .B2(new_n429), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT105), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n410), .A2(G15gat), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n619), .B2(new_n632), .ZN(G1326gat));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n361), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT43), .B(G22gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(G1327gat));
  NAND2_X1  g435(.A1(new_n436), .A2(new_n588), .ZN(new_n637));
  INV_X1    g436(.A(new_n617), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n524), .A2(new_n544), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n548), .A3(new_n620), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT45), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n612), .A2(new_n614), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n588), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n425), .B2(new_n435), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT44), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n645), .A2(new_n647), .A3(new_n650), .A4(new_n640), .ZN(new_n651));
  OAI21_X1  g450(.A(G29gat), .B1(new_n651), .B2(new_n414), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n643), .A2(new_n652), .ZN(G1328gat));
  INV_X1    g452(.A(new_n419), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n641), .A2(new_n549), .A3(new_n654), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n655), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(KEYINPUT46), .ZN(new_n657));
  OAI21_X1  g456(.A(G36gat), .B1(new_n651), .B2(new_n419), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT106), .B1(new_n655), .B2(KEYINPUT46), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n659), .ZN(G1329gat));
  INV_X1    g459(.A(new_n410), .ZN(new_n661));
  OAI21_X1  g460(.A(G43gat), .B1(new_n651), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT47), .B1(new_n662), .B2(KEYINPUT107), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n641), .A2(new_n556), .A3(new_n429), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n662), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n663), .B(new_n665), .ZN(G1330gat));
  AND4_X1   g465(.A1(new_n333), .A2(new_n639), .A3(new_n360), .A4(new_n640), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n651), .A2(new_n361), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(G50gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g469(.A(new_n524), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n425), .B2(new_n435), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n647), .A2(new_n588), .A3(new_n545), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n414), .B(KEYINPUT108), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g477(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n419), .B(KEYINPUT109), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n675), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT110), .ZN(new_n683));
  NOR2_X1   g482(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1333gat));
  NAND3_X1  g484(.A1(new_n675), .A2(G71gat), .A3(new_n410), .ZN(new_n686));
  INV_X1    g485(.A(G71gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n674), .B2(new_n430), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT111), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT111), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n360), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g495(.A1(new_n647), .A2(new_n544), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n645), .A2(new_n524), .A3(new_n650), .A4(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G85gat), .B1(new_n698), .B2(new_n414), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT51), .ZN(new_n700));
  INV_X1    g499(.A(new_n697), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n637), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n649), .A2(KEYINPUT51), .A3(new_n697), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n524), .A2(new_n455), .A3(new_n620), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT112), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n699), .B1(new_n705), .B2(new_n707), .ZN(G1336gat));
  NAND4_X1  g507(.A1(new_n704), .A2(new_n264), .A3(new_n524), .A4(new_n681), .ZN(new_n709));
  OAI21_X1  g508(.A(G92gat), .B1(new_n698), .B2(new_n680), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT52), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G92gat), .B1(new_n698), .B2(new_n419), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT113), .B(G92gat), .C1(new_n698), .C2(new_n419), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n715), .A2(new_n709), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n712), .B1(new_n717), .B2(new_n711), .ZN(G1337gat));
  INV_X1    g517(.A(G99gat), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n698), .A2(new_n719), .A3(new_n661), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n524), .A3(new_n429), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n719), .B2(new_n721), .ZN(G1338gat));
  XNOR2_X1  g521(.A(KEYINPUT114), .B(G106gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n698), .B2(new_n361), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT115), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(G106gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n704), .A2(new_n727), .A3(new_n524), .A4(new_n360), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT115), .B(new_n723), .C1(new_n698), .C2(new_n361), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT53), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT117), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n698), .A2(new_n732), .A3(new_n361), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n698), .B2(new_n361), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n723), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n728), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n731), .A2(new_n737), .ZN(G1339gat));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT54), .B1(new_n499), .B2(new_n477), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n515), .B2(new_n516), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n522), .B1(new_n520), .B2(KEYINPUT54), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n742), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n504), .A2(new_n505), .ZN(new_n745));
  OAI211_X1 g544(.A(KEYINPUT55), .B(new_n744), .C1(new_n745), .C2(new_n740), .ZN(new_n746));
  AND4_X1   g545(.A1(new_n647), .A2(new_n519), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n595), .B1(new_n592), .B2(new_n594), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n599), .A2(new_n600), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n607), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n611), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n519), .B2(new_n523), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n648), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n751), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n519), .A2(new_n743), .A3(new_n746), .A4(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n648), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n544), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n671), .A2(new_n673), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT118), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n524), .A2(new_n754), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n519), .A2(new_n647), .A3(new_n743), .A4(new_n746), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n588), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n545), .B1(new_n764), .B2(new_n756), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(new_n759), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n681), .A2(new_n414), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n431), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G113gat), .B1(new_n770), .B2(new_n638), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n768), .A2(new_n426), .A3(new_n676), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n680), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n646), .A2(G113gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT120), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n773), .A2(new_n778), .ZN(G1340gat));
  INV_X1    g578(.A(G120gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n775), .A2(new_n780), .A3(new_n524), .ZN(new_n781));
  OAI21_X1  g580(.A(G120gat), .B1(new_n770), .B2(new_n671), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1341gat));
  NOR3_X1   g582(.A1(new_n770), .A2(new_n287), .A3(new_n545), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n775), .A2(new_n544), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n287), .ZN(G1342gat));
  INV_X1    g585(.A(G134gat), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n654), .A2(new_n648), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n774), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT56), .ZN(new_n790));
  OAI21_X1  g589(.A(G134gat), .B1(new_n770), .B2(new_n648), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(KEYINPUT56), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(G1343gat));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n410), .A2(new_n361), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n761), .A2(new_n795), .A3(new_n676), .A4(new_n767), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n681), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n638), .A2(G141gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT122), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n769), .A2(new_n661), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n617), .A2(new_n519), .A3(new_n743), .A4(new_n746), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n762), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n648), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n544), .B1(new_n804), .B2(new_n757), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n360), .B1(new_n805), .B2(new_n760), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n801), .B1(new_n806), .B2(KEYINPUT57), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n761), .A2(new_n808), .A3(new_n360), .A4(new_n767), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G141gat), .B1(new_n810), .B2(new_n638), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n812), .A3(new_n798), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n800), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n797), .A2(KEYINPUT121), .A3(new_n798), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT121), .B1(new_n797), .B2(new_n798), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n807), .A2(new_n647), .A3(new_n809), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n794), .B1(new_n818), .B2(G141gat), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n794), .A2(new_n814), .B1(new_n817), .B2(new_n819), .ZN(G1344gat));
  INV_X1    g619(.A(G148gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n797), .A2(new_n821), .A3(new_n524), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n761), .A2(new_n360), .A3(new_n767), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT57), .ZN(new_n825));
  INV_X1    g624(.A(new_n801), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n589), .A2(new_n638), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n804), .A2(new_n757), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n545), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n808), .A3(new_n360), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n825), .A2(new_n524), .A3(new_n826), .A4(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n821), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT57), .B1(new_n829), .B2(new_n831), .ZN(new_n837));
  AOI22_X1  g636(.A1(KEYINPUT57), .A2(new_n824), .B1(new_n837), .B2(new_n360), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(KEYINPUT125), .A3(new_n524), .A4(new_n826), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n823), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n807), .A2(new_n524), .A3(new_n809), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n823), .A3(G148gat), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n841), .A2(KEYINPUT123), .A3(new_n823), .A4(G148gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n822), .B1(new_n840), .B2(new_n846), .ZN(G1345gat));
  NOR3_X1   g646(.A1(new_n810), .A2(new_n292), .A3(new_n545), .ZN(new_n848));
  AOI21_X1  g647(.A(G155gat), .B1(new_n797), .B2(new_n544), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n810), .B2(new_n648), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n788), .A2(new_n293), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n796), .B2(new_n852), .ZN(G1347gat));
  NOR2_X1   g652(.A1(new_n676), .A2(new_n419), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n768), .A2(new_n431), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G169gat), .B1(new_n855), .B2(new_n638), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n761), .A2(new_n414), .A3(new_n681), .A4(new_n767), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(new_n427), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n209), .A3(new_n647), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1348gat));
  NOR3_X1   g659(.A1(new_n855), .A2(new_n210), .A3(new_n671), .ZN(new_n861));
  AOI21_X1  g660(.A(G176gat), .B1(new_n858), .B2(new_n524), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(G1349gat));
  OAI21_X1  g662(.A(G183gat), .B1(new_n855), .B2(new_n545), .ZN(new_n864));
  INV_X1    g663(.A(new_n858), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n544), .A2(new_n203), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT60), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n864), .B(new_n869), .C1(new_n865), .C2(new_n866), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n855), .B2(new_n648), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n865), .A2(new_n218), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT126), .B1(new_n876), .B2(new_n588), .ZN(new_n877));
  AND4_X1   g676(.A1(KEYINPUT126), .A2(new_n858), .A3(new_n588), .A4(new_n202), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n874), .B(new_n875), .C1(new_n877), .C2(new_n878), .ZN(G1351gat));
  NOR3_X1   g678(.A1(new_n410), .A2(new_n419), .A3(new_n676), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n838), .A2(new_n617), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G197gat), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n857), .A2(new_n361), .A3(new_n410), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n646), .A2(G197gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1352gat));
  NAND4_X1  g685(.A1(new_n825), .A2(new_n524), .A3(new_n833), .A4(new_n880), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G204gat), .ZN(new_n888));
  INV_X1    g687(.A(new_n857), .ZN(new_n889));
  INV_X1    g688(.A(G204gat), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n524), .A4(new_n795), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT62), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n883), .A2(new_n893), .A3(new_n890), .A4(new_n524), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n888), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT127), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n888), .A2(new_n892), .A3(new_n894), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1353gat));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n244), .A3(new_n544), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n838), .A2(new_n544), .A3(new_n880), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n901), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT63), .B1(new_n901), .B2(G211gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(G1354gat));
  NAND3_X1  g703(.A1(new_n883), .A2(new_n245), .A3(new_n588), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n838), .A2(new_n588), .A3(new_n880), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n245), .ZN(G1355gat));
endmodule


