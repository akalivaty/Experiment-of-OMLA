//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n216), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G250), .B(G257), .Z(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n231), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G68), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n214), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n206), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI22_X1  g0053(.A1(new_n252), .A2(new_n253), .B1(new_n206), .B2(G68), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n247), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT11), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT71), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n205), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G68), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(KEYINPUT12), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n257), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n256), .B(new_n264), .C1(KEYINPUT12), .C2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n247), .B1(new_n259), .B2(new_n260), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G1), .B2(new_n206), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n268), .B2(KEYINPUT12), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n279), .A2(new_n233), .A3(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n276), .A2(new_n278), .A3(G226), .A4(new_n280), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G97), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n274), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n205), .B(G274), .C1(G41), .C2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n273), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n273), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g0091(.A(G238), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AND4_X1   g0092(.A1(new_n271), .A2(new_n285), .A3(new_n286), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n286), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n273), .A2(new_n288), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n289), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n294), .B1(new_n297), .B2(G238), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n271), .B1(new_n298), .B2(new_n285), .ZN(new_n299));
  OAI21_X1  g0099(.A(G169), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n293), .A2(new_n299), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n300), .A2(KEYINPUT14), .B1(new_n301), .B2(G179), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n285), .A2(new_n286), .A3(new_n292), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT13), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n298), .A2(new_n271), .A3(new_n285), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(G179), .A3(new_n306), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n307), .B2(new_n308), .ZN(new_n313));
  AOI211_X1 g0113(.A(KEYINPUT14), .B(new_n303), .C1(new_n305), .C2(new_n306), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n270), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n301), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n270), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n301), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT3), .B(G33), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(G222), .A3(new_n280), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(G223), .A3(G1698), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n325), .B(new_n326), .C1(new_n253), .C2(new_n324), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n273), .B1(new_n327), .B2(KEYINPUT68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(KEYINPUT68), .B2(new_n327), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n294), .B1(new_n297), .B2(G226), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n303), .ZN(new_n332));
  INV_X1    g0132(.A(new_n247), .ZN(new_n333));
  INV_X1    g0133(.A(G58), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n275), .A2(G20), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT8), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT70), .B1(new_n341), .B2(G58), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n339), .B(new_n340), .C1(new_n337), .C2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n250), .A2(new_n334), .A3(new_n263), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(G20), .B1(G150), .B2(new_n248), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n333), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n265), .A2(new_n250), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n333), .B1(G1), .B2(new_n206), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n250), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n332), .B(new_n352), .C1(G179), .C2(new_n331), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n347), .A2(KEYINPUT9), .A3(new_n351), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(new_n357), .C1(new_n318), .C2(new_n331), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n331), .A2(G200), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT10), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n356), .A2(new_n357), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n329), .A2(new_n330), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G190), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT10), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .A4(new_n359), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n354), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n268), .A2(new_n253), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G20), .A2(G77), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT8), .B(G58), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n369), .B1(new_n370), .B2(new_n252), .C1(new_n249), .C2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n372), .A2(new_n247), .B1(new_n253), .B2(new_n262), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT72), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n324), .A2(G238), .A3(G1698), .ZN(new_n377));
  INV_X1    g0177(.A(G107), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n324), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n279), .A2(new_n233), .A3(G1698), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n274), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n297), .A2(G244), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n286), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G190), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT72), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n374), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(G200), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n376), .A2(new_n385), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G179), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n383), .A2(new_n303), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(new_n374), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n323), .A2(new_n367), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G20), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n248), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n277), .A2(G33), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n206), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT75), .B1(new_n277), .B2(G33), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(new_n275), .A3(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n407), .A3(new_n278), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n401), .A2(G20), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n401), .A2(new_n404), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n400), .B1(new_n410), .B2(new_n263), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n333), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT74), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n401), .B1(new_n324), .B2(G20), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n399), .B1(new_n417), .B2(G68), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n414), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n263), .B1(new_n415), .B2(new_n416), .ZN(new_n420));
  NOR4_X1   g0220(.A1(new_n420), .A2(KEYINPUT74), .A3(new_n399), .A4(new_n412), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n413), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n339), .B1(new_n337), .B2(new_n342), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n257), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n349), .B(new_n339), .C1(new_n337), .C2(new_n342), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(G223), .A2(G1698), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n280), .A2(G226), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n324), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n273), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n286), .B1(new_n295), .B2(new_n233), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n432), .A2(new_n390), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n274), .ZN(new_n436));
  INV_X1    g0236(.A(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(G169), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT76), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n439), .B1(new_n422), .B2(new_n426), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT76), .A3(KEYINPUT18), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  INV_X1    g0246(.A(new_n426), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT7), .B1(new_n279), .B2(new_n206), .ZN(new_n448));
  AOI211_X1 g0248(.A(new_n401), .B(G20), .C1(new_n276), .C2(new_n278), .ZN(new_n449));
  OAI21_X1  g0249(.A(G68), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT74), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n418), .A2(new_n414), .A3(KEYINPUT16), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n447), .B1(new_n454), .B2(new_n413), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n446), .B1(new_n455), .B2(new_n439), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n443), .A2(new_n445), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(G200), .B1(new_n436), .B2(new_n437), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n432), .A2(G190), .A3(new_n433), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n422), .A2(new_n426), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT17), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT77), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n395), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n457), .A2(KEYINPUT77), .A3(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n468), .B(new_n206), .C1(G33), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G20), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n247), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n470), .A2(KEYINPUT20), .A3(new_n247), .A4(new_n472), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n471), .B1(new_n205), .B2(G33), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n475), .A2(new_n476), .B1(new_n267), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT83), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n261), .B2(G116), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n259), .A2(KEYINPUT83), .A3(new_n471), .A4(new_n260), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n478), .A2(new_n482), .A3(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT78), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(G41), .ZN(new_n490));
  INV_X1    g0290(.A(G41), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(G45), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G1), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G270), .A3(new_n273), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(new_n273), .A3(new_n490), .A4(new_n492), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n276), .A2(new_n278), .A3(G257), .A4(new_n280), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT81), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT81), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n324), .A2(new_n503), .A3(G257), .A4(new_n280), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n279), .A2(G303), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n324), .A2(G264), .A3(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n502), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n507), .A2(new_n508), .A3(new_n274), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n507), .B2(new_n274), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n487), .A2(KEYINPUT21), .A3(G169), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n487), .A2(G169), .A3(new_n511), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(G200), .ZN(new_n516));
  OAI211_X1 g0316(.A(G190), .B(new_n500), .C1(new_n509), .C2(new_n510), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n485), .A3(new_n486), .A4(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G179), .B(new_n500), .C1(new_n509), .C2(new_n510), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n487), .ZN(new_n521));
  AND4_X1   g0321(.A1(new_n512), .A2(new_n515), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n276), .A2(new_n278), .A3(G250), .A4(new_n280), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n276), .A2(new_n278), .A3(G257), .A4(G1698), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n274), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n495), .A2(G264), .A3(new_n273), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n498), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G169), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(KEYINPUT88), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT88), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n495), .A2(new_n535), .A3(G264), .A4(new_n273), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(new_n536), .B1(new_n274), .B2(new_n527), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(G179), .A3(new_n498), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(KEYINPUT87), .A3(G169), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n533), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n276), .A2(new_n278), .A3(new_n206), .A4(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT22), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT22), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n324), .A2(new_n543), .A3(new_n206), .A4(G87), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g0345(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G20), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT23), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n206), .B2(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n378), .A2(KEYINPUT23), .A3(G20), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n545), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n546), .B1(new_n545), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n247), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n205), .A2(G33), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n333), .A2(new_n257), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n378), .B1(KEYINPUT86), .B2(KEYINPUT25), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n257), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n265), .A2(KEYINPUT86), .A3(KEYINPUT25), .A4(new_n378), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n557), .A2(G107), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n540), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(G200), .B1(new_n537), .B2(new_n498), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n530), .A2(G190), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n555), .B(new_n562), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT89), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT89), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n564), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n370), .B(KEYINPUT80), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n557), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n324), .A2(new_n206), .A3(G68), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n206), .B1(new_n283), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G87), .B2(new_n203), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n252), .B2(new_n469), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n247), .B1(new_n262), .B2(new_n370), .ZN(new_n582));
  INV_X1    g0382(.A(new_n497), .ZN(new_n583));
  OAI21_X1  g0383(.A(G250), .B1(new_n493), .B2(G1), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n274), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n324), .A2(G238), .A3(new_n280), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n324), .A2(G244), .A3(G1698), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n547), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n588), .B2(new_n274), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n575), .A2(new_n582), .B1(new_n589), .B2(new_n390), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n274), .ZN(new_n591));
  INV_X1    g0391(.A(new_n585), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n303), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(G200), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n557), .A2(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n589), .A2(G190), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(new_n582), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n469), .A2(new_n378), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n202), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n378), .A2(KEYINPUT6), .A3(G97), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n605), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n378), .B2(new_n410), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n247), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n257), .A2(G97), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n557), .B2(G97), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n276), .A2(new_n278), .A3(G244), .A4(new_n280), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT4), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n324), .A2(KEYINPUT4), .A3(G244), .A4(new_n280), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n324), .A2(G250), .A3(G1698), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n468), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n274), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n495), .A2(G257), .A3(new_n273), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n498), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n303), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n617), .B2(new_n274), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n390), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n611), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(G200), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT79), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(G190), .B2(new_n624), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n624), .A2(new_n628), .A3(G190), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n608), .A3(new_n610), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n600), .B(new_n626), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n572), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n467), .A2(new_n523), .A3(new_n634), .ZN(G372));
  NOR2_X1   g0435(.A1(new_n322), .A2(new_n393), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n463), .B1(new_n316), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n638));
  AOI211_X1 g0438(.A(new_n446), .B(new_n439), .C1(new_n422), .C2(new_n426), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n361), .A2(new_n366), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n354), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n626), .B1(new_n629), .B2(new_n631), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n596), .A2(new_n598), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n582), .A2(new_n597), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT90), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n582), .A2(KEYINPUT90), .A3(new_n597), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n567), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n515), .A2(new_n564), .A3(new_n512), .A4(new_n521), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n654), .A2(new_n655), .B1(new_n594), .B2(new_n590), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n595), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n626), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n595), .A2(new_n599), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n626), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n644), .B1(new_n467), .B2(new_n664), .ZN(G369));
  AOI22_X1  g0465(.A1(new_n513), .A2(new_n514), .B1(new_n487), .B2(new_n520), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n512), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n487), .A2(new_n673), .ZN(new_n674));
  MUX2_X1   g0474(.A(new_n667), .B(new_n522), .S(new_n674), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n563), .A2(new_n673), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n572), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n673), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n678), .B1(new_n564), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n564), .A2(new_n673), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n667), .A2(new_n679), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n686), .B2(new_n572), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n209), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n212), .B2(new_n691), .ZN(new_n694));
  XOR2_X1   g0494(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n695));
  XNOR2_X1  g0495(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n673), .B1(new_n656), .B2(new_n663), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n657), .B2(new_n626), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n660), .A2(new_n661), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n673), .B1(new_n656), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n698), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n572), .A2(new_n522), .A3(new_n633), .A4(new_n679), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n624), .A2(new_n537), .A3(new_n589), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n519), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n507), .A2(new_n274), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT82), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n507), .A2(new_n508), .A3(new_n274), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n499), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n624), .A2(new_n537), .A3(new_n589), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(KEYINPUT30), .A4(G179), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT92), .B1(new_n591), .B2(new_n592), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT92), .ZN(new_n718));
  AOI211_X1 g0518(.A(new_n718), .B(new_n585), .C1(new_n588), .C2(new_n274), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n537), .A2(new_n498), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n624), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n511), .A2(new_n720), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n710), .A2(new_n716), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT31), .B1(new_n724), .B2(new_n673), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n707), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n673), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(KEYINPUT93), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n706), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n705), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n696), .B1(new_n736), .B2(G1), .ZN(G364));
  AND2_X1   g0537(.A1(new_n206), .A2(G13), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n205), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n690), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n675), .B2(G330), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n675), .ZN(new_n743));
  XOR2_X1   g0543(.A(KEYINPUT33), .B(G317), .Z(new_n744));
  NOR2_X1   g0544(.A1(new_n390), .A2(new_n320), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n206), .A2(G190), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n279), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n206), .A2(new_n318), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n745), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n390), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G326), .A2(new_n751), .B1(new_n754), .B2(G322), .ZN(new_n755));
  INV_X1    g0555(.A(G303), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n320), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n746), .A2(new_n752), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n755), .B1(new_n756), .B2(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n206), .B1(new_n762), .B2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n748), .B(new_n761), .C1(G294), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n746), .A2(new_n757), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n746), .A2(new_n762), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G283), .A2(new_n767), .B1(new_n769), .B2(G329), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT97), .Z(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n768), .A2(KEYINPUT32), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT32), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n769), .B2(G159), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n773), .B(new_n775), .C1(G97), .C2(new_n764), .ZN(new_n776));
  INV_X1    g0576(.A(new_n760), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G50), .A2(new_n751), .B1(new_n777), .B2(G77), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n263), .B2(new_n747), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n766), .A2(new_n378), .ZN(new_n780));
  INV_X1    g0580(.A(G87), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n334), .A2(new_n753), .B1(new_n758), .B2(new_n781), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n779), .A2(new_n279), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n765), .A2(new_n771), .B1(new_n776), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n214), .B1(G20), .B2(new_n303), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n741), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n209), .A2(G116), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n689), .A2(new_n324), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G45), .B2(new_n212), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(new_n241), .B2(G45), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n209), .A2(new_n324), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n793), .B(new_n796), .C1(G355), .C2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n792), .B(new_n785), .C1(new_n799), .C2(KEYINPUT95), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n799), .A2(KEYINPUT95), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n787), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n675), .B2(new_n791), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n743), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  OAI21_X1  g0605(.A(new_n389), .B1(new_n375), .B2(new_n679), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n393), .ZN(new_n807));
  INV_X1    g0607(.A(new_n393), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n679), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n697), .B(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n741), .B1(new_n812), .B2(new_n734), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n734), .B2(new_n812), .ZN(new_n814));
  INV_X1    g0614(.A(new_n741), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n785), .A2(new_n788), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n253), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n747), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G143), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n753), .A2(new_n820), .B1(new_n760), .B2(new_n772), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n821), .C1(G137), .C2(new_n751), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n822), .A2(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(KEYINPUT34), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n324), .B1(new_n768), .B2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n758), .A2(new_n250), .B1(new_n766), .B2(new_n263), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G58), .C2(new_n764), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n823), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n766), .A2(new_n781), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n747), .A2(new_n831), .B1(new_n760), .B2(new_n471), .ZN(new_n832));
  INV_X1    g0632(.A(new_n758), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n830), .B(new_n832), .C1(G107), .C2(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n750), .A2(new_n756), .B1(new_n768), .B2(new_n759), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n324), .B(new_n835), .C1(G294), .C2(new_n754), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n469), .C2(new_n763), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n817), .B1(new_n786), .B2(new_n838), .C1(new_n811), .C2(new_n789), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n814), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  OR2_X1    g0641(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n605), .A2(KEYINPUT35), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n842), .A2(G116), .A3(new_n215), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT36), .Z(new_n845));
  OAI211_X1 g0645(.A(new_n213), .B(G77), .C1(new_n334), .C2(new_n263), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n250), .A2(G68), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n205), .B(G13), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n466), .B(new_n465), .C1(new_n699), .C2(new_n704), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n644), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT103), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n456), .B1(new_n639), .B2(KEYINPUT76), .ZN(new_n853));
  INV_X1    g0653(.A(new_n445), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n463), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n247), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n453), .A2(new_n452), .B1(new_n856), .B2(KEYINPUT99), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT99), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n858), .B(new_n247), .C1(new_n418), .C2(KEYINPUT16), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n447), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n671), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n462), .B1(new_n860), .B2(new_n439), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n864), .B2(KEYINPUT100), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT100), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n866), .B(new_n462), .C1(new_n860), .C2(new_n439), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n427), .A2(new_n440), .ZN(new_n869));
  INV_X1    g0669(.A(new_n671), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n408), .A2(new_n409), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n415), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n399), .B1(new_n872), .B2(G68), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n247), .B1(new_n873), .B2(KEYINPUT16), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n453), .B2(new_n452), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n870), .B1(new_n875), .B2(new_n447), .ZN(new_n876));
  AND4_X1   g0676(.A1(new_n863), .A2(new_n869), .A3(new_n876), .A4(new_n462), .ZN(new_n877));
  OAI211_X1 g0677(.A(KEYINPUT38), .B(new_n862), .C1(new_n868), .C2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n450), .B2(new_n400), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT99), .B1(new_n880), .B2(new_n333), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n454), .A2(new_n859), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n439), .B1(new_n882), .B2(new_n426), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n447), .B(new_n460), .C1(new_n454), .C2(new_n413), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT100), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n882), .A2(new_n426), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n870), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n867), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n877), .B1(new_n888), .B2(KEYINPUT37), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n457), .B2(new_n463), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n878), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n809), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n697), .B2(new_n811), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n270), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT73), .B1(new_n302), .B2(new_n309), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n313), .A2(new_n311), .A3(new_n314), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n322), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n270), .A2(new_n679), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI211_X1 g0703(.A(KEYINPUT98), .B(new_n902), .C1(new_n310), .C2(new_n315), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT98), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n310), .A2(new_n315), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n901), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n903), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n892), .A2(new_n895), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n641), .B2(new_n870), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n316), .A2(new_n679), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n892), .A2(KEYINPUT39), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n884), .A2(new_n444), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n863), .B1(new_n913), .B2(new_n876), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT101), .B1(new_n914), .B2(new_n877), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n462), .B1(new_n455), .B2(new_n439), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n455), .A2(new_n671), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT101), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n869), .A2(new_n876), .A3(new_n863), .A4(new_n462), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT17), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n462), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n884), .A2(KEYINPUT17), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(new_n638), .C2(new_n639), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n917), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n915), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n879), .ZN(new_n928));
  XOR2_X1   g0728(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n878), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n911), .B1(new_n912), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n910), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n852), .B(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(G330), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n878), .A2(new_n891), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n725), .A2(new_n726), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n810), .B1(new_n706), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT104), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT40), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n908), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n908), .A2(new_n938), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n939), .A2(new_n943), .B1(new_n928), .B2(new_n878), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n942), .B1(new_n944), .B2(new_n935), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n467), .B1(new_n937), .B2(new_n706), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n934), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n945), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n933), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n951), .B1(new_n205), .B2(new_n738), .C1(new_n933), .C2(new_n948), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n849), .B1(new_n952), .B2(new_n953), .ZN(G367));
  AOI21_X1  g0754(.A(new_n679), .B1(new_n608), .B2(new_n610), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n645), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n626), .B2(new_n679), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(new_n686), .A3(new_n572), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT42), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n626), .B1(new_n956), .B2(new_n564), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n679), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n651), .A2(new_n679), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(new_n595), .A3(new_n652), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT106), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n966), .A2(new_n967), .B1(new_n595), .B2(new_n965), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n966), .ZN(new_n969));
  NOR2_X1   g0769(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n970));
  AND2_X1   g0770(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT43), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n963), .B(new_n972), .C1(new_n973), .C2(new_n969), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(new_n963), .C2(new_n972), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n682), .A2(new_n957), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n977), .B(new_n978), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n690), .B(KEYINPUT41), .Z(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n687), .A2(KEYINPUT109), .A3(new_n957), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT109), .B1(new_n687), .B2(new_n957), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n687), .A2(new_n957), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT45), .Z(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n682), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n986), .A2(new_n683), .A3(new_n987), .A4(new_n989), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n681), .A2(new_n685), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n686), .A2(new_n572), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n676), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n676), .B1(new_n995), .B2(new_n996), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n735), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n994), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n992), .A2(new_n993), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n982), .B1(new_n1003), .B2(new_n735), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n980), .B1(new_n1004), .B2(new_n739), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n792), .A2(new_n785), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n209), .B2(new_n370), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n230), .A2(new_n689), .A3(new_n324), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n741), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n750), .A2(new_n820), .B1(new_n758), .B2(new_n334), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n279), .B(new_n1010), .C1(G150), .C2(new_n754), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G77), .A2(new_n767), .B1(new_n769), .B2(G137), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n747), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G159), .A2(new_n1013), .B1(new_n777), .B2(G50), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n764), .A2(G68), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(KEYINPUT111), .B(G317), .Z(new_n1017));
  OAI22_X1  g0817(.A1(new_n759), .A2(new_n750), .B1(new_n1017), .B2(new_n768), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G283), .B2(new_n777), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n324), .B1(new_n1013), .B2(G294), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G303), .A2(new_n754), .B1(new_n767), .B2(G97), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n833), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT46), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n758), .B2(new_n471), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n378), .C2(new_n763), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1016), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT47), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1009), .B1(new_n1028), .B2(new_n785), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT112), .Z(new_n1030));
  NAND2_X1  g0830(.A1(new_n969), .A2(new_n792), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1005), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT113), .ZN(G387));
  INV_X1    g0834(.A(new_n1001), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1000), .A2(new_n735), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n690), .A3(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n833), .A2(G294), .B1(new_n764), .B2(G283), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G322), .A2(new_n751), .B1(new_n1013), .B2(G311), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n756), .B2(new_n760), .C1(new_n753), .C2(new_n1017), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT49), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n324), .B1(new_n769), .B2(G326), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n471), .B2(new_n766), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n574), .A2(new_n764), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n750), .A2(new_n772), .B1(new_n768), .B2(new_n818), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n758), .A2(new_n253), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n279), .B1(new_n767), .B2(G97), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G50), .A2(new_n754), .B1(new_n777), .B2(G68), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n423), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n1013), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n785), .B1(new_n1047), .B2(new_n1056), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n236), .A2(new_n493), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n692), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1058), .A2(new_n794), .B1(new_n1059), .B2(new_n798), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT50), .B1(new_n371), .B2(G50), .ZN(new_n1061));
  AOI21_X1  g0861(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n692), .A3(new_n1062), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n371), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1060), .A2(new_n1065), .B1(G107), .B2(new_n209), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n815), .B1(new_n1066), .B2(new_n1006), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n681), .B2(new_n792), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1000), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n740), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1037), .A2(new_n1071), .ZN(G393));
  NAND2_X1  g0872(.A1(new_n991), .A2(new_n994), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n691), .B1(new_n1073), .B2(new_n1035), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n992), .A2(new_n1002), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n993), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1073), .A2(new_n739), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n957), .A2(new_n791), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1006), .B1(new_n469), .B2(new_n209), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n794), .A2(new_n244), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n741), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n750), .A2(new_n818), .B1(new_n753), .B2(new_n772), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n747), .A2(new_n250), .B1(new_n760), .B2(new_n371), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT114), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n758), .A2(new_n263), .B1(new_n768), .B2(new_n820), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n763), .A2(new_n253), .ZN(new_n1087));
  NOR4_X1   g0887(.A1(new_n1086), .A2(new_n830), .A3(new_n1087), .A4(new_n279), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1083), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n751), .B1(new_n754), .B2(G311), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n324), .B(new_n780), .C1(G116), .C2(new_n764), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G303), .A2(new_n1013), .B1(new_n777), .B2(G294), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G283), .A2(new_n833), .B1(new_n769), .B2(G322), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1089), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1081), .B1(new_n1096), .B2(new_n785), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1077), .B1(new_n1078), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1076), .A2(new_n1098), .ZN(G390));
  NAND2_X1  g0899(.A1(new_n706), .A2(new_n937), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n465), .A2(G330), .A3(new_n466), .A4(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n850), .A2(new_n644), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n893), .B1(new_n703), .B2(new_n807), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n934), .B(new_n810), .C1(new_n706), .C2(new_n937), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n908), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n733), .A2(G330), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT115), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1106), .A2(new_n1107), .A3(new_n811), .A4(new_n908), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n908), .A2(new_n733), .A3(G330), .A4(new_n811), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT115), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1105), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n907), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n904), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1112), .A2(new_n1113), .B1(new_n323), .B2(new_n902), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n734), .B2(new_n810), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1104), .A2(new_n908), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n894), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1102), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT116), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n911), .B1(new_n894), .B2(new_n1114), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n912), .A2(new_n1120), .A3(new_n930), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n928), .A2(new_n878), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1123), .B(new_n911), .C1(new_n1114), .C2(new_n1103), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1116), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1118), .B(new_n1119), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n850), .A2(new_n644), .A3(new_n1101), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1105), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1109), .A2(KEYINPUT115), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1109), .A2(KEYINPUT115), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1117), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1128), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1116), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1127), .A2(new_n1139), .A3(new_n690), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT116), .B1(new_n1142), .B2(new_n1134), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n912), .A2(new_n788), .A3(new_n930), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n816), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n751), .A2(G128), .B1(new_n769), .B2(G125), .ZN(new_n1147));
  INV_X1    g0947(.A(G137), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n747), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n324), .B1(new_n753), .B2(new_n825), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n250), .A2(new_n766), .B1(new_n760), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n758), .A2(new_n818), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1153), .B(new_n1155), .C1(new_n772), .C2(new_n763), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n279), .B1(new_n758), .B2(new_n781), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT117), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n750), .A2(new_n831), .B1(new_n747), .B2(new_n378), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n753), .A2(new_n471), .B1(new_n766), .B2(new_n263), .ZN(new_n1160));
  INV_X1    g0960(.A(G294), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n760), .A2(new_n469), .B1(new_n768), .B2(new_n1161), .ZN(new_n1162));
  OR4_X1    g0962(.A1(new_n1087), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1156), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1165), .A2(KEYINPUT118), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n785), .B1(new_n1165), .B2(KEYINPUT118), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n741), .B1(new_n1055), .B2(new_n1146), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1141), .A2(new_n739), .B1(new_n1145), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1144), .A2(new_n1170), .ZN(G378));
  OR2_X1    g0971(.A1(new_n910), .A2(new_n931), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n352), .A2(new_n870), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n367), .B(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n918), .A2(new_n920), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1177), .A2(KEYINPUT101), .B1(new_n917), .B2(new_n925), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT38), .B1(new_n1178), .B2(new_n921), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n889), .A2(new_n879), .A3(new_n890), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT104), .B1(new_n908), .B2(new_n938), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT40), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n934), .B(new_n1176), .C1(new_n1183), .C2(new_n942), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1176), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n945), .B2(G330), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1172), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n943), .A2(new_n939), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n1123), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1189), .A2(KEYINPUT40), .B1(new_n936), .B2(new_n941), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1176), .B1(new_n1190), .B2(new_n934), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n945), .A2(G330), .A3(new_n1185), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n932), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1139), .A2(new_n1102), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n690), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n741), .B1(new_n1146), .B2(G50), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1185), .A2(new_n789), .ZN(new_n1201));
  INV_X1    g1001(.A(G128), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1202), .A2(new_n753), .B1(new_n758), .B2(new_n1151), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT121), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n764), .A2(G150), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1013), .A2(G132), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G125), .A2(new_n751), .B1(new_n777), .B2(G137), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1209));
  XNOR2_X1  g1009(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n275), .B(new_n491), .C1(new_n766), .C2(new_n772), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G124), .B2(new_n769), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(KEYINPUT3), .A2(G33), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G50), .B1(new_n1214), .B2(new_n491), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT119), .Z(new_n1216));
  NAND2_X1  g1016(.A1(new_n574), .A2(new_n777), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n753), .A2(new_n378), .B1(new_n768), .B2(new_n831), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1218), .A2(new_n1050), .A3(G41), .A4(new_n324), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n750), .A2(new_n471), .B1(new_n766), .B2(new_n334), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G97), .B2(new_n1013), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1217), .A2(new_n1219), .A3(new_n1015), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT120), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1213), .B(new_n1225), .C1(new_n1223), .C2(new_n1222), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1200), .B(new_n1201), .C1(new_n785), .C2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1194), .B2(new_n740), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1199), .A2(new_n1228), .ZN(G375));
  OAI22_X1  g1029(.A1(new_n758), .A2(new_n772), .B1(new_n760), .B2(new_n818), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n747), .A2(new_n1151), .B1(new_n768), .B2(new_n1202), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n324), .B1(new_n766), .B2(new_n334), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n750), .A2(new_n825), .B1(new_n753), .B2(new_n1148), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(G50), .C2(new_n764), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n750), .A2(new_n1161), .B1(new_n747), .B2(new_n471), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n758), .A2(new_n469), .B1(new_n760), .B2(new_n378), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n753), .A2(new_n831), .B1(new_n768), .B2(new_n756), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n279), .B1(new_n766), .B2(new_n253), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1232), .A2(new_n1235), .B1(new_n1240), .B2(new_n1048), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n741), .B1(G68), .B2(new_n1146), .C1(new_n1241), .C2(new_n786), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1114), .B2(new_n788), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1243), .B1(new_n1244), .B2(new_n740), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1118), .A2(new_n982), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1244), .A2(new_n1102), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(G381));
  AOI21_X1  g1048(.A(new_n1169), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1199), .A2(new_n1249), .A3(new_n1228), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1037), .A2(new_n804), .A3(new_n1071), .ZN(new_n1251));
  OR3_X1    g1051(.A1(G390), .A2(G384), .A3(new_n1251), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G387), .A2(new_n1250), .A3(G381), .A4(new_n1252), .ZN(G407));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  INV_X1    g1054(.A(new_n1005), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1032), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n804), .B1(new_n1037), .B2(new_n1071), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1251), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT113), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1076), .A2(new_n1098), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1076), .A2(new_n1098), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1255), .B(new_n1256), .C1(new_n1263), .C2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G390), .A2(new_n1259), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1266), .B(new_n1262), .C1(new_n1005), .C2(new_n1032), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1247), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n690), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1269), .A2(new_n1247), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1245), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n840), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n672), .A2(G213), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G384), .B(new_n1245), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1277));
  AND4_X1   g1077(.A1(G2897), .A2(new_n1274), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1274), .A2(new_n1277), .B1(G2897), .B2(new_n1276), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G378), .B(new_n1228), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1194), .A2(new_n1195), .A3(new_n982), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1228), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1284), .A2(new_n1285), .A3(new_n1249), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1284), .B2(new_n1249), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1282), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1275), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1281), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT62), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1276), .B1(new_n1288), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1292), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1282), .B(KEYINPUT124), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1268), .B1(new_n1294), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1288), .A2(new_n1297), .A3(KEYINPUT63), .A4(new_n1275), .ZN(new_n1303));
  AND4_X1   g1103(.A1(new_n1291), .A2(new_n1303), .A3(new_n1265), .A4(new_n1267), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1288), .A2(new_n1295), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1275), .A3(new_n1298), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1305), .B1(new_n1307), .B2(new_n1281), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1292), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1302), .B(new_n1304), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1280), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1299), .B1(new_n1312), .B2(new_n1305), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1302), .B1(new_n1313), .B2(new_n1304), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1301), .B1(new_n1311), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT126), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1317), .B(new_n1301), .C1(new_n1311), .C2(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(G405));
  INV_X1    g1119(.A(new_n1268), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1249), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1321), .A2(new_n1297), .A3(new_n1282), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1297), .B1(new_n1321), .B2(new_n1282), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1320), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1320), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .ZN(G402));
endmodule


