//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n251), .A3(G274), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n256), .A2(G226), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  OR2_X1    g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n261), .A2(G223), .B1(new_n264), .B2(G77), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n260), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G222), .A3(new_n258), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n269));
  AOI211_X1 g0069(.A(new_n253), .B(new_n257), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G179), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n216), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n207), .A2(G20), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G50), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT8), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  INV_X1    g0089(.A(G58), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(KEYINPUT68), .A2(KEYINPUT8), .A3(G58), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n208), .A2(G33), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n284), .B1(new_n285), .B2(new_n287), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n295), .A2(new_n276), .B1(new_n296), .B2(new_n280), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n283), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n272), .B(new_n298), .C1(G169), .C2(new_n270), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  AOI22_X1  g0100(.A1(G190), .A2(new_n270), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n270), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n283), .A2(new_n297), .A3(KEYINPUT9), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT69), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n305), .B1(new_n304), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n299), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n274), .B(KEYINPUT67), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n219), .A2(G20), .ZN(new_n312));
  INV_X1    g0112(.A(G33), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(G20), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(G77), .B1(new_n286), .B2(G50), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT12), .B1(new_n280), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  INV_X1    g0120(.A(new_n278), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n312), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n280), .A2(new_n274), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n207), .B2(G20), .ZN(new_n324));
  AOI211_X1 g0124(.A(new_n319), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n316), .A2(KEYINPUT11), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n317), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n266), .A2(G226), .A3(new_n258), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT70), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT70), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n266), .A2(new_n330), .A3(G226), .A4(new_n258), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n251), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n251), .A2(G238), .A3(new_n254), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n252), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n252), .A2(new_n338), .A3(KEYINPUT71), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT73), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n342), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT73), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n335), .B1(new_n331), .B2(new_n329), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n345), .B(new_n346), .C1(new_n347), .C2(new_n251), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n344), .A2(KEYINPUT13), .A3(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n345), .B(new_n350), .C1(new_n347), .C2(new_n251), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G179), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  INV_X1    g0153(.A(new_n350), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n337), .B2(new_n343), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n355), .B2(new_n351), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n349), .A2(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n327), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n351), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n327), .B1(new_n362), .B2(G200), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n344), .A2(KEYINPUT13), .A3(new_n348), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n351), .A2(G190), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n293), .B1(new_n207), .B2(G20), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n281), .A2(new_n370), .B1(new_n280), .B2(new_n293), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n287), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n202), .B1(new_n219), .B2(new_n290), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n372), .B(new_n374), .C1(new_n375), .C2(G20), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n318), .A2(KEYINPUT64), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT64), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G68), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n290), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n380), .B2(new_n201), .ZN(new_n381));
  INV_X1    g0181(.A(new_n374), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT74), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n259), .A2(new_n208), .A3(new_n260), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n260), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(KEYINPUT75), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT75), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n390), .A3(new_n386), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n220), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT16), .B1(new_n384), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n378), .A2(G68), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n318), .A2(KEYINPUT64), .ZN(new_n395));
  OAI21_X1  g0195(.A(G58), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n208), .B1(new_n396), .B2(new_n202), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n372), .B1(new_n397), .B2(new_n374), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n387), .A2(new_n388), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(G68), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n381), .A2(KEYINPUT74), .A3(new_n382), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n274), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n371), .B1(new_n393), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n258), .A2(G226), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n266), .B(new_n406), .C1(G223), .C2(G1698), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n251), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G232), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n252), .B1(new_n410), .B2(new_n255), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G179), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n353), .B2(new_n412), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n405), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  INV_X1    g0218(.A(G190), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n412), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n302), .B1(new_n409), .B2(new_n411), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n371), .B(new_n422), .C1(new_n393), .C2(new_n404), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT17), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n371), .ZN(new_n426));
  INV_X1    g0226(.A(new_n274), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n384), .B2(new_n401), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n398), .A2(new_n392), .A3(new_n402), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n399), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT17), .A3(new_n422), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n416), .A2(new_n418), .A3(new_n425), .A4(new_n432), .ZN(new_n433));
  XOR2_X1   g0233(.A(KEYINPUT15), .B(G87), .Z(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n294), .ZN(new_n436));
  XNOR2_X1  g0236(.A(KEYINPUT8), .B(G58), .ZN(new_n437));
  INV_X1    g0237(.A(G77), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n437), .A2(new_n287), .B1(new_n208), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n274), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n282), .A2(G77), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n323), .A2(new_n442), .B1(new_n438), .B2(new_n280), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n261), .A2(G238), .B1(new_n264), .B2(G107), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n266), .A2(G232), .A3(new_n258), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n251), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n256), .A2(G244), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n447), .A2(new_n253), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n444), .B1(new_n449), .B2(G190), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n302), .B2(new_n449), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n271), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n444), .C1(G169), .C2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR4_X1   g0254(.A1(new_n310), .A2(new_n369), .A3(new_n433), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G20), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n321), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n207), .A2(G33), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n456), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n323), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n274), .A2(new_n457), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT80), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n274), .A2(KEYINPUT80), .A3(new_n457), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(G20), .B1(G33), .B2(G283), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(G33), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT20), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n274), .A2(KEYINPUT80), .A3(new_n457), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT80), .B1(new_n274), .B2(new_n457), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT20), .B(new_n470), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n462), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n248), .A2(G1), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT5), .B(G41), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n269), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n478), .A2(new_n477), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n269), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n479), .A2(G270), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G264), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n484));
  OAI211_X1 g0284(.A(G257), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n259), .A2(G303), .A3(new_n260), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT79), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n487), .A2(new_n488), .A3(new_n269), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n487), .B2(new_n269), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n483), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n476), .B1(G200), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n419), .B2(new_n491), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n476), .A2(KEYINPUT21), .A3(G169), .A4(new_n491), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n479), .A2(G270), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n480), .A2(new_n482), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n487), .A2(new_n269), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT79), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n487), .A2(new_n488), .A3(new_n269), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n476), .A2(new_n501), .A3(G179), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n476), .A2(G169), .A3(new_n491), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n493), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G257), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n508));
  OAI211_X1 g0308(.A(G250), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n269), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n479), .A2(G264), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n496), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n302), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G190), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n208), .B(G87), .C1(new_n262), .C2(new_n263), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(KEYINPUT22), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n266), .A2(new_n208), .A3(G87), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT24), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n208), .B2(G107), .ZN(new_n526));
  INV_X1    g0326(.A(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(KEYINPUT23), .A3(G20), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n526), .A2(new_n528), .B1(new_n314), .B2(G116), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n524), .B1(new_n523), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n274), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n279), .A2(G107), .ZN(new_n533));
  XOR2_X1   g0333(.A(KEYINPUT82), .B(KEYINPUT25), .Z(new_n534));
  XNOR2_X1  g0334(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n311), .A2(new_n279), .A3(new_n459), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(G107), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n516), .A2(new_n532), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n514), .A2(G169), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n511), .A2(new_n269), .B1(new_n479), .B2(G264), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G179), .A3(new_n496), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n532), .A2(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT83), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n532), .A2(new_n538), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n542), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT83), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n516), .A2(new_n532), .A3(new_n538), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(G33), .B2(G283), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT76), .B1(new_n261), .B2(G250), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT76), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n269), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n479), .A2(G257), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n496), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(G179), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n269), .B2(new_n560), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n353), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT78), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n389), .A2(G107), .A3(new_n391), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n527), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n469), .A2(new_n527), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n204), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n572), .B2(KEYINPUT6), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(G20), .B1(G77), .B2(new_n286), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n274), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n279), .A2(G97), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n536), .B2(new_n469), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n568), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n427), .B1(new_n569), .B2(new_n574), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n582), .A2(new_n579), .A3(KEYINPUT78), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n567), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n566), .A2(G190), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n582), .A2(new_n579), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n566), .B2(KEYINPUT77), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n561), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n434), .A2(new_n279), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n208), .B1(new_n334), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G87), .B2(new_n205), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n208), .B(G68), .C1(new_n262), .C2(new_n263), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n294), .B2(new_n469), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n590), .B1(new_n596), .B2(new_n274), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n311), .A2(G87), .A3(new_n279), .A4(new_n459), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n251), .A2(G274), .A3(new_n477), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n207), .A2(G45), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n251), .A2(G250), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G244), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n603));
  OAI211_X1 g0403(.A(G238), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n313), .C2(new_n456), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n605), .B2(new_n269), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n597), .B(new_n598), .C1(new_n606), .C2(new_n302), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n419), .B(new_n602), .C1(new_n269), .C2(new_n605), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n597), .B1(new_n435), .B2(new_n536), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n606), .A2(G169), .ZN(new_n611));
  AOI211_X1 g0411(.A(G179), .B(new_n602), .C1(new_n269), .C2(new_n605), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n584), .A2(new_n589), .A3(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n455), .A2(new_n507), .A3(new_n551), .A4(new_n615), .ZN(G372));
  OR2_X1    g0416(.A1(new_n308), .A2(new_n309), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n432), .A2(new_n425), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n367), .A2(new_n453), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n361), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n416), .A2(new_n418), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n622), .A2(new_n299), .ZN(new_n623));
  INV_X1    g0423(.A(new_n455), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n608), .B1(new_n607), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n605), .A2(new_n269), .ZN(new_n627));
  OAI21_X1  g0427(.A(G200), .B1(new_n627), .B2(new_n602), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(KEYINPUT84), .A3(new_n597), .A4(new_n598), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n626), .A2(new_n629), .B1(new_n610), .B2(new_n613), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n584), .A2(new_n589), .A3(new_n630), .A4(new_n549), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT85), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n494), .A2(new_n502), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n499), .A2(new_n500), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n353), .B1(new_n634), .B2(new_n483), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT21), .B1(new_n635), .B2(new_n476), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n506), .A2(KEYINPUT85), .A3(new_n502), .A4(new_n494), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n631), .B1(new_n639), .B2(new_n547), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n613), .A2(new_n610), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n608), .B2(new_n607), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT26), .B1(new_n584), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n586), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n567), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(new_n630), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n647), .A3(new_n641), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n623), .B1(new_n624), .B2(new_n649), .ZN(G369));
  OR3_X1    g0450(.A1(new_n321), .A2(KEYINPUT27), .A3(G20), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n321), .B2(G20), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n476), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n507), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n639), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G330), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n545), .A2(new_n655), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n551), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n543), .A2(new_n655), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n547), .A2(new_n655), .ZN(new_n667));
  INV_X1    g0467(.A(new_n655), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n633), .B2(new_n636), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT87), .Z(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n211), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n214), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n633), .A2(new_n636), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n547), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT88), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT88), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n683), .A3(new_n547), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n631), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n584), .A2(new_n642), .A3(KEYINPUT26), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n645), .A2(new_n630), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n686), .B(new_n641), .C1(new_n687), .C2(new_n646), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n668), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT29), .ZN(new_n690));
  INV_X1    g0490(.A(new_n649), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n668), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n551), .A2(new_n615), .A3(new_n507), .A4(new_n668), .ZN(new_n694));
  OAI211_X1 g0494(.A(G179), .B(new_n483), .C1(new_n489), .C2(new_n490), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n541), .A2(new_n606), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n566), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n606), .A2(G179), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n514), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n566), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n698), .A2(new_n699), .B1(new_n702), .B2(new_n491), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n696), .A2(KEYINPUT30), .A3(new_n566), .A4(new_n697), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n668), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT31), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n698), .A2(new_n699), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n702), .A2(new_n491), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n655), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n694), .A2(new_n706), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n690), .A2(new_n693), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n679), .B1(new_n716), .B2(G1), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT89), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n277), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n207), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n674), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n658), .A2(G330), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n659), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n245), .A2(G45), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT90), .Z(new_n726));
  NAND2_X1  g0526(.A1(new_n211), .A2(new_n264), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT91), .Z(new_n728));
  OAI211_X1 g0528(.A(new_n726), .B(new_n728), .C1(G45), .C2(new_n214), .ZN(new_n729));
  INV_X1    g0529(.A(G355), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n211), .A2(new_n266), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n729), .B1(G116), .B2(new_n211), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n216), .B1(G20), .B2(new_n353), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n208), .A2(new_n271), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n419), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G326), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n208), .A2(G179), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n741), .A2(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n739), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT33), .B(G317), .Z(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(new_n419), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(G283), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n302), .A2(G190), .ZN(new_n754));
  OAI21_X1  g0554(.A(G20), .B1(new_n754), .B2(G179), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT95), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G294), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n743), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G329), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n738), .A2(new_n762), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n754), .A2(new_n208), .A3(new_n271), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n266), .B(new_n771), .C1(G322), .C2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n753), .A2(new_n761), .A3(new_n768), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n266), .B1(new_n769), .B2(new_n438), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G58), .B2(new_n772), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n750), .A2(new_n527), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(G50), .B2(new_n740), .ZN(new_n778));
  INV_X1    g0578(.A(G87), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n744), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(G68), .B2(new_n747), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n776), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n760), .A2(G97), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n767), .A2(G159), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n784), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n766), .B2(new_n373), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n783), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n774), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n732), .A2(new_n737), .B1(new_n736), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n735), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n658), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n724), .B1(new_n722), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT96), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  NAND2_X1  g0595(.A1(new_n444), .A2(new_n655), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n451), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n453), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n453), .A2(new_n655), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n649), .B2(new_n655), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n454), .A2(new_n655), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n640), .B2(new_n648), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n714), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT98), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT98), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n722), .B1(new_n805), .B2(new_n806), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n736), .A2(new_n733), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n722), .B1(G77), .B2(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n741), .A2(new_n745), .B1(new_n750), .B2(new_n779), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT97), .B(G283), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n748), .A2(new_n816), .B1(new_n744), .B2(new_n527), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n767), .A2(G311), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n264), .B1(new_n769), .B2(new_n456), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G294), .B2(new_n772), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n818), .A2(new_n783), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n769), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n823), .A2(G159), .B1(new_n772), .B2(G143), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n285), .B2(new_n748), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G137), .B2(new_n740), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n266), .B1(new_n750), .B2(new_n318), .ZN(new_n828));
  INV_X1    g0628(.A(new_n744), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(G50), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n766), .B2(new_n831), .C1(new_n290), .C2(new_n759), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n822), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n814), .B1(new_n833), .B2(new_n736), .ZN(new_n834));
  INV_X1    g0634(.A(new_n801), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n734), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n812), .A2(new_n836), .ZN(G384));
  OR2_X1    g0637(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n573), .A2(KEYINPUT35), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n838), .A2(G116), .A3(new_n217), .A4(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT36), .Z(new_n841));
  NAND3_X1  g0641(.A1(new_n215), .A2(G77), .A3(new_n396), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n296), .A2(G68), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n207), .B(G13), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n690), .A2(new_n693), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n455), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n847), .A2(new_n623), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT103), .ZN(new_n849));
  INV_X1    g0649(.A(new_n653), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n416), .B2(new_n418), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n804), .A2(new_n800), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n327), .A2(new_n655), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n361), .A2(new_n368), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n362), .A2(G169), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT14), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n364), .A2(G179), .A3(new_n351), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n359), .A3(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n327), .B(new_n655), .C1(new_n858), .C2(new_n367), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n400), .A2(G68), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT16), .B1(new_n384), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n403), .A2(new_n276), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n371), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n850), .A2(new_n866), .B1(new_n431), .B2(new_n422), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n414), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n414), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n423), .B1(new_n431), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n428), .A2(new_n430), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n653), .B1(new_n872), .B2(new_n371), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n871), .A2(KEYINPUT37), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT100), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n311), .B1(new_n384), .B2(new_n401), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n398), .A2(new_n402), .A3(new_n863), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n399), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n426), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n423), .B1(new_n879), .B2(new_n653), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n870), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT100), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n405), .A2(new_n850), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n415), .A2(new_n884), .A3(new_n862), .A4(new_n423), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n879), .A2(new_n653), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n433), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n875), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n886), .A4(new_n888), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n861), .A2(KEYINPUT99), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n860), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n804), .B2(new_n800), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT99), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n851), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n858), .A2(new_n327), .A3(new_n668), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n433), .A2(new_n873), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n871), .B2(new_n873), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n885), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n882), .A2(new_n885), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n909), .A2(KEYINPUT100), .B1(new_n433), .B2(new_n887), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT102), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT38), .A4(new_n886), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n907), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n900), .B(new_n901), .C1(new_n913), .C2(KEYINPUT39), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n898), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n849), .B(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n801), .B1(new_n854), .B2(new_n859), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT104), .B1(new_n705), .B2(KEYINPUT31), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT104), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n710), .A2(new_n919), .A3(new_n711), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n694), .A2(new_n918), .A3(new_n920), .A4(new_n706), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n917), .A2(new_n921), .A3(KEYINPUT40), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n908), .A2(new_n912), .ZN(new_n923));
  INV_X1    g0723(.A(new_n907), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n917), .A2(new_n921), .ZN(new_n927));
  INV_X1    g0727(.A(new_n892), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n910), .B2(new_n886), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n926), .A2(new_n455), .A3(new_n921), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G330), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n926), .A2(new_n932), .B1(new_n455), .B2(new_n921), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n916), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n207), .B2(new_n719), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n916), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n845), .B1(new_n938), .B2(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n665), .A2(new_n670), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n584), .B(new_n589), .C1(new_n586), .C2(new_n668), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n645), .A2(new_n655), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n941), .A2(KEYINPUT42), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n584), .B1(new_n945), .B2(new_n547), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n668), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT42), .B1(new_n941), .B2(new_n945), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n597), .A2(new_n598), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n655), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n641), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n630), .B2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT43), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT106), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n666), .A2(new_n945), .ZN(new_n962));
  INV_X1    g0762(.A(new_n960), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n950), .A2(new_n963), .A3(new_n956), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n666), .B2(new_n945), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n674), .B(KEYINPUT41), .Z(new_n968));
  NAND2_X1  g0768(.A1(new_n671), .A2(new_n944), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  OR3_X1    g0772(.A1(new_n671), .A2(new_n972), .A3(new_n944), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n671), .B2(new_n944), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n666), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n665), .B(new_n670), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n659), .A2(KEYINPUT107), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n715), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n971), .A2(new_n975), .A3(new_n666), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n978), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n968), .B1(new_n984), .B2(new_n716), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n965), .B(new_n967), .C1(new_n985), .C2(new_n721), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n728), .A2(new_n238), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n737), .C1(new_n211), .C2(new_n435), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n748), .A2(new_n373), .B1(new_n744), .B2(new_n290), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n767), .A2(G137), .ZN(new_n990));
  INV_X1    g0790(.A(G143), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n741), .A2(new_n991), .B1(new_n750), .B2(new_n438), .ZN(new_n992));
  INV_X1    g0792(.A(new_n772), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n266), .B1(new_n296), .B2(new_n769), .C1(new_n993), .C2(new_n285), .ZN(new_n994));
  OR4_X1    g0794(.A1(new_n989), .A2(new_n990), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n759), .A2(new_n318), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n264), .B1(new_n769), .B2(new_n816), .C1(new_n993), .C2(new_n745), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n829), .A2(G116), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n998), .B2(new_n999), .C1(new_n1001), .C2(new_n766), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n750), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n747), .A2(G294), .B1(new_n1003), .B2(G97), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n770), .B2(new_n741), .C1(new_n759), .C2(new_n527), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n995), .A2(new_n996), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  INV_X1    g0807(.A(new_n736), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n722), .B(new_n988), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n954), .A2(new_n735), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n986), .A2(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n981), .A2(new_n715), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT112), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n982), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(KEYINPUT112), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n674), .B(KEYINPUT111), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n981), .A2(new_n720), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n662), .A2(new_n664), .A3(new_n735), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n731), .A2(new_n676), .B1(G107), .B2(new_n211), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n728), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n235), .B2(G45), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n437), .A2(G50), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n248), .B1(new_n318), .B2(new_n438), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n676), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT108), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1026), .B(new_n1029), .C1(KEYINPUT108), .C2(new_n1028), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1022), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n737), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n722), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n741), .A2(new_n373), .B1(new_n750), .B2(new_n469), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n748), .A2(new_n293), .B1(new_n438), .B2(new_n744), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n760), .A2(new_n434), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n767), .A2(G150), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n266), .B1(new_n993), .B2(new_n296), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G68), .B2(new_n823), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n993), .A2(new_n1001), .B1(new_n769), .B2(new_n745), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT109), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n747), .A2(G311), .B1(new_n740), .B2(G322), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n816), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n760), .A2(new_n1050), .B1(G294), .B2(new_n829), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT49), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT110), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n266), .B1(new_n1003), .B2(G116), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n742), .C2(new_n766), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1053), .A2(KEYINPUT110), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1041), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1033), .B1(new_n1058), .B2(new_n736), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1020), .B1(new_n1021), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1019), .A2(new_n1060), .ZN(G393));
  INV_X1    g0861(.A(new_n983), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n666), .B1(new_n971), .B2(new_n975), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1016), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(new_n984), .A3(new_n1018), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n728), .A2(new_n242), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n737), .C1(new_n469), .C2(new_n211), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n760), .A2(G77), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n296), .B2(new_n748), .C1(new_n437), .C2(new_n769), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n740), .A2(G150), .B1(G159), .B2(new_n772), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT51), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n264), .B1(new_n1003), .B2(G87), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n219), .B2(new_n744), .C1(new_n766), .C2(new_n991), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT113), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n740), .A2(G317), .B1(G311), .B2(new_n772), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT52), .Z(new_n1077));
  NAND2_X1  g0877(.A1(new_n767), .A2(G322), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n266), .B(new_n777), .C1(G294), .C2(new_n823), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n747), .A2(G303), .B1(new_n829), .B2(new_n1050), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G116), .B2(new_n760), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1072), .A2(new_n1075), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n722), .B(new_n1067), .C1(new_n1083), .C2(new_n1008), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n945), .B2(new_n735), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n721), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1065), .A2(new_n1087), .ZN(G390));
  INV_X1    g0888(.A(new_n293), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n722), .B1(new_n1089), .B2(new_n813), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n527), .A2(new_n748), .B1(new_n741), .B2(new_n751), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n780), .B(new_n1091), .C1(G68), .C2(new_n1003), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n767), .A2(G294), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n264), .B1(new_n993), .B2(new_n456), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G97), .B2(new_n823), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1092), .A2(new_n1068), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n744), .A2(new_n285), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT54), .B(G143), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n266), .B1(new_n769), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G132), .B2(new_n772), .ZN(new_n1101));
  INV_X1    g0901(.A(G125), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1098), .B(new_n1101), .C1(new_n1102), .C2(new_n766), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n740), .A2(G128), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n747), .A2(G137), .B1(new_n1003), .B2(G50), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n759), .C2(new_n373), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1096), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1090), .B1(new_n1107), .B2(new_n736), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n923), .A2(new_n924), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT39), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1108), .B1(new_n1112), .B2(new_n734), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n668), .B(new_n798), .C1(new_n685), .C2(new_n688), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n860), .B1(new_n1115), .B2(new_n799), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1110), .A2(new_n1116), .A3(new_n899), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n806), .A2(new_n835), .A3(new_n860), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n895), .A2(new_n900), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1117), .B(new_n1118), .C1(new_n1112), .C2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n901), .B1(new_n913), .B2(KEYINPUT39), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1119), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n913), .A2(new_n900), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1121), .A2(new_n1122), .B1(new_n1123), .B2(new_n1116), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n917), .A2(new_n921), .A3(G330), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1113), .B1(new_n1126), .B2(new_n720), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n455), .A2(G330), .A3(new_n921), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n847), .A2(new_n623), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n860), .B1(new_n806), .B2(new_n835), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1125), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n852), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n921), .A2(G330), .A3(new_n835), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n894), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1118), .A2(new_n800), .A3(new_n1134), .A4(new_n1114), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1129), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1120), .B(new_n1136), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1137), .A2(new_n1018), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1136), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1126), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1127), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(G378));
  AND2_X1   g0942(.A1(new_n898), .A2(new_n914), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n298), .A2(new_n850), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n617), .A2(new_n299), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n310), .A2(new_n298), .A3(new_n850), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(G330), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n930), .B2(new_n931), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n926), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n917), .A2(new_n921), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n891), .B2(new_n892), .ZN(new_n1158));
  OAI21_X1  g0958(.A(G330), .B1(new_n1158), .B2(KEYINPUT40), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1159), .A2(new_n925), .A3(new_n1152), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1143), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n926), .A2(new_n1155), .A3(new_n1153), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1152), .B1(new_n1159), .B2(new_n925), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n915), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(KEYINPUT116), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT116), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1162), .A2(new_n915), .A3(new_n1163), .A4(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n721), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n722), .B1(G50), .B2(new_n813), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n264), .A2(new_n247), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n434), .B2(new_n823), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n527), .B2(new_n993), .C1(new_n766), .C2(new_n751), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n748), .A2(new_n469), .B1(new_n744), .B2(new_n438), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n741), .A2(new_n456), .B1(new_n750), .B2(new_n290), .ZN(new_n1174));
  OR4_X1    g0974(.A1(new_n996), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1170), .B(new_n296), .C1(G33), .C2(G41), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1180), .B2(KEYINPUT114), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n823), .A2(G137), .B1(new_n772), .B2(G128), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n744), .B2(new_n1099), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G132), .B2(new_n747), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n760), .A2(G150), .B1(G125), .B2(new_n740), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1185), .A2(KEYINPUT115), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(KEYINPUT115), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1184), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n767), .A2(G124), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n1003), .C2(G159), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1181), .B1(KEYINPUT114), .B2(new_n1180), .C1(new_n1189), .C2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1169), .B1(new_n1194), .B2(new_n736), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1152), .B2(new_n734), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1168), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT117), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT117), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1168), .A2(new_n1199), .A3(new_n1196), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1129), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1137), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT118), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1162), .A2(new_n915), .A3(new_n1163), .A4(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1161), .A2(KEYINPUT118), .A3(new_n1164), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(KEYINPUT57), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1203), .A2(new_n1167), .A3(new_n1165), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1018), .B(new_n1207), .C1(new_n1208), .C2(KEYINPUT57), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1201), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(G375));
  INV_X1    g1011(.A(new_n968), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1129), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1139), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT119), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n720), .B(KEYINPUT120), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n894), .A2(new_n733), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n722), .B1(G68), .B2(new_n813), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1037), .B1(new_n751), .B2(new_n993), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT121), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n264), .B1(new_n769), .B2(new_n527), .C1(new_n438), .C2(new_n750), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n747), .A2(G116), .B1(new_n740), .B2(G294), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n469), .B2(new_n744), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1222), .B(new_n1224), .C1(G303), .C2(new_n767), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT122), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n264), .B1(new_n1003), .B2(G58), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n760), .A2(G50), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n823), .A2(G150), .B1(new_n772), .B2(G137), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n748), .B2(new_n1099), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n741), .A2(new_n831), .B1(new_n744), .B2(new_n373), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n767), .A2(G128), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1228), .A2(new_n1227), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1229), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1226), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1219), .B1(new_n1237), .B2(new_n736), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1216), .A2(new_n1217), .B1(new_n1218), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1215), .A2(new_n1239), .ZN(G381));
  NAND2_X1  g1040(.A1(new_n1210), .A2(new_n1141), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  INV_X1    g1042(.A(G390), .ZN(new_n1243));
  INV_X1    g1043(.A(G384), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  OR4_X1    g1045(.A1(G387), .A2(new_n1241), .A3(G381), .A4(new_n1245), .ZN(G407));
  OAI211_X1 g1046(.A(G407), .B(G213), .C1(G343), .C2(new_n1241), .ZN(G409));
  AOI21_X1  g1047(.A(new_n794), .B1(new_n1019), .B2(new_n1060), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n986), .A2(new_n1012), .A3(G390), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G390), .B1(new_n986), .B2(new_n1012), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n967), .A2(new_n965), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n984), .A2(new_n716), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1212), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1255), .B2(new_n720), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1243), .B1(new_n1256), .B2(new_n1011), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n986), .A2(new_n1012), .A3(G390), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n654), .A2(G213), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1203), .A2(new_n1212), .A3(new_n1167), .A4(new_n1165), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1206), .A2(new_n1205), .A3(new_n1217), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1196), .A3(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1268), .A2(KEYINPUT123), .A3(new_n1141), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT123), .B1(new_n1268), .B2(new_n1141), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1201), .A2(G378), .A3(new_n1209), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1265), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1213), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1213), .A2(new_n1274), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1139), .A3(new_n1018), .A4(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1277), .A2(G384), .A3(new_n1239), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1277), .B2(new_n1239), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(G2897), .A3(new_n1265), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1265), .A2(G2897), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1262), .B(new_n1263), .C1(new_n1273), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1270), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1268), .A2(KEYINPUT123), .A3(new_n1141), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1272), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n1264), .A3(new_n1280), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT62), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1273), .A2(new_n1292), .A3(new_n1280), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1286), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1264), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1284), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1262), .B1(new_n1296), .B2(new_n1263), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1261), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1252), .A2(new_n1263), .A3(new_n1260), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT126), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1289), .A2(KEYINPUT63), .A3(new_n1264), .A4(new_n1280), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(KEYINPUT125), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1273), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1305), .A3(new_n1284), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT124), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1290), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1307), .B1(new_n1290), .B2(new_n1308), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1302), .B(new_n1306), .C1(new_n1309), .C2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1298), .A2(new_n1311), .ZN(G405));
  XNOR2_X1  g1112(.A(new_n1210), .B(G378), .ZN(new_n1313));
  OR2_X1    g1113(.A1(new_n1313), .A2(new_n1280), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1280), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1261), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1314), .A2(new_n1260), .A3(new_n1252), .A4(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


