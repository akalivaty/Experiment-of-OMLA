//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1259, new_n1260, new_n1261;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  XOR2_X1   g028(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n460), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(new_n463), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n471), .B1(new_n462), .B2(G2104), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n469), .A2(G137), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT68), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(G160));
  NAND3_X1  g051(.A1(new_n469), .A2(G2105), .A3(new_n472), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n477), .A2(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n469), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n486), .B1(new_n470), .B2(G114), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI211_X1 g067(.A(KEYINPUT70), .B(new_n485), .C1(new_n487), .C2(new_n489), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n484), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n472), .A2(new_n468), .A3(new_n496), .A4(new_n463), .ZN(new_n497));
  INV_X1    g072(.A(new_n464), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n494), .A2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n505), .A2(new_n507), .A3(G62), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n517), .A2(new_n518), .A3(new_n505), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n517), .B2(new_n505), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n514), .B2(new_n516), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n511), .A2(new_n522), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  XNOR2_X1  g102(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n530), .A2(new_n531), .B1(new_n505), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n523), .B1(new_n517), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n514), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G51), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n517), .A2(new_n505), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT72), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n517), .A2(new_n518), .A3(new_n505), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n540), .A2(G89), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n541), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n517), .A2(new_n534), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(G543), .A3(new_n536), .ZN(new_n548));
  INV_X1    g123(.A(G52), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n513), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n546), .A2(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n503), .A2(new_n504), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n558), .B2(new_n548), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(G81), .B2(new_n521), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT76), .Z(G188));
  AND2_X1   g141(.A1(KEYINPUT77), .A2(G53), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n535), .A2(new_n536), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n535), .A2(new_n570), .A3(new_n536), .A4(new_n567), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n513), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n521), .B2(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  OR2_X1    g152(.A1(new_n538), .A2(new_n542), .ZN(G286));
  NAND3_X1  g153(.A1(new_n540), .A2(G87), .A3(new_n541), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n580));
  INV_X1    g155(.A(G49), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n548), .ZN(G288));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  NOR3_X1   g158(.A1(new_n519), .A2(new_n520), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n524), .A2(G48), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n513), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AND2_X1   g164(.A1(new_n521), .A2(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n548), .A2(new_n591), .B1(new_n513), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n590), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n554), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  INV_X1    g174(.A(G54), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n548), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n544), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(G868), .B2(new_n606), .ZN(G284));
  OAI21_X1  g182(.A(new_n595), .B1(G868), .B2(new_n606), .ZN(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n609), .B2(G168), .ZN(G280));
  XNOR2_X1  g187(.A(KEYINPUT78), .B(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(G860), .B2(new_n613), .ZN(G148));
  INV_X1    g189(.A(G81), .ZN(new_n615));
  OAI221_X1 g190(.A(new_n557), .B1(new_n548), .B2(new_n558), .C1(new_n544), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n609), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n606), .A2(new_n613), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n619), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n623));
  INV_X1    g198(.A(G111), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n622), .A2(new_n623), .B1(new_n624), .B2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n623), .B2(new_n622), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n477), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G135), .B2(new_n482), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n460), .A2(G2105), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n498), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT13), .B(G2100), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n630), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2454), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(KEYINPUT84), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(KEYINPUT84), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT82), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2451), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n655), .B1(new_n650), .B2(new_n651), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n642), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n641), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT85), .Z(new_n664));
  OAI21_X1  g239(.A(G14), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n641), .B1(new_n660), .B2(new_n656), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT86), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n670), .B(new_n664), .C1(new_n666), .C2(new_n667), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n665), .B1(new_n669), .B2(new_n671), .ZN(G401));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2100), .ZN(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n676), .B2(KEYINPUT18), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2096), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n688), .A2(new_n693), .A3(new_n691), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(KEYINPUT20), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n688), .B2(new_n693), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n692), .B(new_n694), .C1(new_n696), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G1981), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(G1981), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n686), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n701), .A2(new_n686), .A3(new_n702), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n685), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(new_n685), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n706), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n706), .B2(new_n709), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(G229));
  NAND2_X1  g290(.A1(G162), .A2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G29), .B2(G35), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT29), .B(G2090), .Z(new_n718));
  XOR2_X1   g293(.A(new_n717), .B(new_n718), .Z(new_n719));
  INV_X1    g294(.A(G1341), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n560), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n721), .B2(G19), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n719), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(G29), .A2(G33), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT25), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n728));
  INV_X1    g303(.A(G139), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n727), .B1(new_n728), .B2(new_n729), .C1(new_n730), .C2(new_n470), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G2072), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G11), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G11), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(G28), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n732), .B1(new_n740), .B2(G28), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n738), .B(new_n739), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n629), .B2(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G34), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT24), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT24), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G160), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n732), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2084), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n482), .A2(G141), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT26), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n755), .A2(new_n756), .B1(G105), .B2(new_n632), .ZN(new_n757));
  INV_X1    g332(.A(G129), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n477), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(new_n732), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n732), .B2(G32), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n751), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n724), .A2(new_n735), .A3(new_n745), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n721), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n721), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1966), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n762), .A2(new_n763), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  NAND2_X1  g345(.A1(G164), .A2(G29), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G27), .B2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n768), .B(new_n773), .C1(new_n770), .C2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n765), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(G171), .A2(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G5), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n779), .B(new_n780), .C1(new_n720), .C2(new_n723), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT97), .B(KEYINPUT23), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n721), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G299), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1956), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n787), .A2(G4), .A3(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(G4), .B2(G16), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n604), .A2(new_n605), .ZN(new_n790));
  INV_X1    g365(.A(new_n601), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n788), .B(new_n789), .C1(new_n792), .C2(new_n721), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n732), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT96), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  AND4_X1   g372(.A1(G2105), .A2(new_n472), .A3(new_n468), .A4(new_n463), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G128), .ZN(new_n799));
  INV_X1    g374(.A(G140), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G116), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n803), .A2(KEYINPUT94), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n799), .B1(new_n728), .B2(new_n800), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n806), .A2(KEYINPUT95), .A3(G29), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(KEYINPUT95), .B1(new_n806), .B2(G29), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n797), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G2067), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n781), .A2(new_n786), .A3(new_n794), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n775), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n721), .A2(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G166), .B2(new_n721), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1971), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT92), .ZN(new_n819));
  NOR2_X1   g394(.A1(G6), .A2(G16), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n588), .B2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT32), .ZN(new_n822));
  INV_X1    g397(.A(G1981), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n721), .A2(G23), .ZN(new_n825));
  INV_X1    g400(.A(G288), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n721), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT33), .B(G1976), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n818), .A2(KEYINPUT92), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n819), .A2(new_n824), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n824), .A2(new_n829), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n835), .A2(new_n832), .A3(new_n819), .A4(new_n830), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n732), .A2(G25), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT89), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(KEYINPUT89), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n798), .A2(G119), .ZN(new_n840));
  OR2_X1    g415(.A1(G95), .A2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n841), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G131), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n728), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT90), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n838), .B(new_n839), .C1(new_n847), .C2(new_n732), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G1991), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n721), .A2(G24), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n590), .A2(new_n593), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(new_n721), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(G1986), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(G1986), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n851), .A2(new_n852), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n834), .A2(new_n836), .A3(new_n859), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(KEYINPUT36), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(KEYINPUT36), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n815), .B1(new_n861), .B2(new_n862), .ZN(G311));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n860), .A2(KEYINPUT36), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n814), .B1(new_n864), .B2(new_n865), .ZN(G150));
  NAND2_X1  g441(.A1(new_n606), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT98), .B(G93), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n544), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n513), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n535), .A2(G55), .A3(new_n536), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT99), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n521), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n873), .A4(new_n872), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n879), .A3(new_n616), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n873), .A3(new_n872), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n560), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n868), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(KEYINPUT39), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT100), .Z(new_n886));
  AOI21_X1  g461(.A(G860), .B1(new_n884), .B2(KEYINPUT39), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n875), .A2(new_n879), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(G860), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT37), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(G145));
  XNOR2_X1  g467(.A(G162), .B(new_n629), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n749), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n728), .A2(new_n800), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G164), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n752), .A2(new_n759), .ZN(new_n900));
  INV_X1    g475(.A(new_n485), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n488), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT69), .B1(new_n488), .B2(G2105), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT70), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n490), .A2(new_n491), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n498), .A2(new_n499), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n910), .A3(new_n484), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n806), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n899), .A2(new_n900), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n900), .B1(new_n899), .B2(new_n912), .ZN(new_n914));
  OAI211_X1 g489(.A(KEYINPUT101), .B(new_n731), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n899), .A2(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n760), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n731), .A2(KEYINPUT101), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n731), .A2(KEYINPUT101), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n899), .A2(new_n900), .A3(new_n912), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n922));
  INV_X1    g497(.A(G118), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n922), .A2(KEYINPUT102), .B1(new_n923), .B2(G2105), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(KEYINPUT102), .B2(new_n922), .ZN(new_n925));
  INV_X1    g500(.A(G130), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n477), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G142), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n728), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n843), .B2(new_n845), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n482), .A2(G131), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(KEYINPUT103), .A3(new_n840), .A4(new_n842), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n930), .B1(new_n934), .B2(new_n932), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n635), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n934), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n927), .B1(G142), .B2(new_n482), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n635), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(new_n935), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n915), .A2(new_n921), .A3(new_n938), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n915), .A2(new_n921), .B1(new_n938), .B2(new_n943), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n895), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n915), .A2(new_n921), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n938), .A2(new_n943), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n894), .A3(new_n944), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n947), .A2(KEYINPUT104), .A3(new_n952), .A4(new_n948), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n880), .A2(new_n882), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n880), .B2(new_n882), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n618), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n962), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(new_n619), .A3(new_n960), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n792), .A2(G299), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT41), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n606), .A2(new_n572), .A3(new_n575), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n967), .B2(new_n969), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G290), .A2(new_n588), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n854), .A2(G305), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(G166), .A2(G288), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n826), .A2(G303), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n975), .A2(new_n978), .A3(new_n979), .A4(new_n976), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n984), .A2(KEYINPUT42), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n981), .A2(new_n984), .A3(KEYINPUT42), .A4(new_n982), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n967), .A2(new_n969), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n963), .A2(new_n965), .A3(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n974), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n991), .B2(new_n974), .ZN(new_n993));
  OAI21_X1  g568(.A(G868), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n889), .A2(new_n609), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(G295));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n996), .ZN(G331));
  INV_X1    g575(.A(new_n983), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n972), .A2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT110), .B(new_n968), .C1(new_n967), .C2(new_n969), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n970), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G286), .A2(G171), .ZN(new_n1008));
  OAI21_X1  g583(.A(G168), .B1(new_n546), .B2(new_n551), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n880), .A2(new_n882), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n880), .A2(new_n882), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1005), .A2(new_n1007), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1012), .A2(new_n967), .A3(new_n969), .A4(new_n1010), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1001), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1010), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n971), .A2(new_n972), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(new_n1014), .A3(KEYINPUT108), .A4(new_n983), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1014), .A3(new_n983), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n1021));
  AOI21_X1  g596(.A(G37), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1016), .A2(KEYINPUT43), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(new_n1014), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n1001), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1024), .A2(new_n1026), .A3(new_n948), .A4(new_n1019), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT44), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1016), .A2(new_n1028), .A3(new_n1019), .A4(new_n1022), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1027), .A2(KEYINPUT43), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(G397));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n494), .B2(new_n500), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(KEYINPUT111), .B(G40), .Z(new_n1042));
  NAND4_X1  g617(.A1(new_n467), .A2(new_n473), .A3(new_n475), .A4(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n846), .B(KEYINPUT112), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n850), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n850), .B2(new_n1046), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n806), .B(new_n811), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n900), .A2(G1996), .ZN(new_n1050));
  INV_X1    g625(.A(G1996), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n760), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1044), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G290), .A2(G1986), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n854), .A2(new_n686), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1045), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT113), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1062));
  NOR2_X1   g637(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1043), .B1(new_n911), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1961), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1040), .A2(G1384), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1043), .B1(new_n911), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G2078), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1041), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n905), .A2(new_n906), .B1(G126), .B2(new_n798), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1384), .B1(new_n1071), .B2(new_n910), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT114), .B1(new_n1072), .B2(KEYINPUT45), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1039), .A2(new_n1074), .A3(new_n1040), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1073), .A2(new_n770), .A3(new_n1067), .A4(new_n1075), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1065), .B(new_n1070), .C1(new_n1076), .C2(new_n1068), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1061), .B1(new_n1077), .B2(G301), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1066), .B1(new_n494), .B2(new_n500), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(G40), .A3(G160), .A4(new_n1069), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT45), .B1(new_n911), .B2(new_n1038), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1065), .B(new_n1082), .C1(new_n1076), .C2(new_n1068), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  OAI21_X1  g659(.A(G171), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1065), .B1(new_n1076), .B2(new_n1068), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1082), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1086), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1078), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(G301), .A3(new_n1087), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1070), .ZN(new_n1091));
  AOI21_X1  g666(.A(G301), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1061), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1043), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n1038), .A3(new_n911), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G8), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G288), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT52), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G8), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1072), .B2(new_n1094), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT116), .B(G1976), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(G288), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1101), .B(new_n1103), .C1(new_n1097), .C2(G288), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G73), .A2(G543), .ZN(new_n1107));
  INV_X1    g682(.A(G61), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n554), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1109), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n540), .A2(G86), .A3(new_n541), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n823), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1106), .A2(KEYINPUT117), .A3(new_n1112), .A4(KEYINPUT49), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT49), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1112), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n823), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1115), .A2(new_n1116), .A3(new_n1120), .A4(new_n1101), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT118), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT49), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1096), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1116), .A4(new_n1115), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1105), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  OR2_X1    g702(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1128));
  NAND3_X1  g703(.A1(G303), .A2(G8), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G166), .A2(new_n1100), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1079), .A2(new_n1094), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1971), .B1(new_n1134), .B2(new_n1073), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(G2090), .ZN(new_n1137));
  OAI211_X1 g712(.A(G8), .B(new_n1132), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1131), .B1(G303), .B2(G8), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1130), .B2(new_n1128), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1073), .A2(new_n1067), .A3(new_n1075), .ZN(new_n1141));
  INV_X1    g716(.A(G1971), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1143));
  INV_X1    g718(.A(G2090), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1140), .B1(new_n1145), .B2(new_n1100), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1127), .A2(new_n1138), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(G1966), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1133), .B2(new_n1081), .ZN(new_n1149));
  INV_X1    g724(.A(G2084), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1062), .A2(new_n1064), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(G168), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1100), .A2(KEYINPUT124), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT51), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1062), .A2(new_n1064), .A3(new_n1150), .ZN(new_n1156));
  AOI21_X1  g731(.A(G1966), .B1(new_n1041), .B2(new_n1067), .ZN(new_n1157));
  OAI211_X1 g732(.A(G8), .B(G286), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1152), .A2(new_n1159), .A3(new_n1153), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1155), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1089), .A2(new_n1093), .A3(new_n1147), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT57), .B1(new_n572), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(G299), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n572), .B(new_n575), .C1(new_n1163), .C2(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT56), .B(G2072), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1073), .A2(new_n1067), .A3(new_n1075), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(G1956), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1136), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1167), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT121), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1167), .A2(new_n1169), .A3(new_n1174), .A4(new_n1171), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n1095), .A2(KEYINPUT122), .A3(G2067), .ZN(new_n1177));
  INV_X1    g752(.A(G1348), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1136), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT122), .B1(new_n1095), .B2(G2067), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n606), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1167), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1176), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1176), .A2(new_n1185), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OR3_X1    g765(.A1(new_n1141), .A2(KEYINPUT123), .A3(G1996), .ZN(new_n1191));
  XOR2_X1   g766(.A(KEYINPUT58), .B(G1341), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n1095), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT123), .B1(new_n1141), .B2(G1996), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n560), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1181), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n606), .A2(KEYINPUT60), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1189), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1202), .A2(new_n1203), .B1(new_n1204), .B2(new_n1172), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1195), .A2(KEYINPUT59), .A3(new_n560), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1190), .A2(new_n1198), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1162), .B1(new_n1187), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1209));
  NOR2_X1   g784(.A1(G288), .A2(G1976), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1096), .B1(new_n1211), .B2(new_n1112), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1105), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1209), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(KEYINPUT119), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT119), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1127), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1138), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1212), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g795(.A(G8), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1221), .A2(new_n1222), .A3(G286), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1146), .A2(new_n1138), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1127), .A2(new_n1216), .ZN(new_n1225));
  AOI211_X1 g800(.A(KEYINPUT119), .B(new_n1105), .C1(new_n1122), .C2(new_n1126), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1221), .A2(G286), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1127), .A2(new_n1138), .A3(new_n1146), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1229), .A2(new_n1222), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  AND4_X1   g806(.A1(new_n1092), .A2(new_n1127), .A3(new_n1138), .A4(new_n1146), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1160), .A2(new_n1158), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1159), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1234));
  OAI21_X1  g809(.A(KEYINPUT62), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1235), .A2(KEYINPUT126), .ZN(new_n1236));
  OR3_X1    g811(.A1(new_n1233), .A2(KEYINPUT62), .A3(new_n1234), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1161), .A2(new_n1238), .A3(KEYINPUT62), .ZN(new_n1239));
  NAND4_X1  g814(.A1(new_n1232), .A2(new_n1236), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1220), .A2(new_n1231), .A3(new_n1240), .ZN(new_n1241));
  OAI21_X1  g816(.A(new_n1060), .B1(new_n1208), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1243));
  XNOR2_X1  g818(.A(new_n1243), .B(KEYINPUT46), .ZN(new_n1244));
  AND2_X1   g819(.A1(new_n1049), .A2(new_n760), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1244), .B1(new_n1045), .B2(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g821(.A(new_n1246), .B(KEYINPUT127), .ZN(new_n1247));
  OR2_X1    g822(.A1(new_n1247), .A2(KEYINPUT47), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1247), .A2(KEYINPUT47), .ZN(new_n1249));
  INV_X1    g824(.A(new_n1055), .ZN(new_n1250));
  NOR2_X1   g825(.A1(new_n1045), .A2(new_n1057), .ZN(new_n1251));
  XOR2_X1   g826(.A(new_n1251), .B(KEYINPUT48), .Z(new_n1252));
  NAND3_X1  g827(.A1(new_n1054), .A2(new_n849), .A3(new_n847), .ZN(new_n1253));
  OAI21_X1  g828(.A(new_n1253), .B1(G2067), .B2(new_n806), .ZN(new_n1254));
  AOI22_X1  g829(.A1(new_n1250), .A2(new_n1252), .B1(new_n1044), .B2(new_n1254), .ZN(new_n1255));
  AND3_X1   g830(.A1(new_n1248), .A2(new_n1249), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1242), .A2(new_n1256), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g832(.A1(G227), .A2(new_n457), .ZN(new_n1259));
  OAI21_X1  g833(.A(new_n1259), .B1(new_n713), .B2(new_n714), .ZN(new_n1260));
  NOR2_X1   g834(.A1(G401), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g835(.A1(new_n1034), .A2(new_n1261), .A3(new_n957), .ZN(G225));
  INV_X1    g836(.A(G225), .ZN(G308));
endmodule


