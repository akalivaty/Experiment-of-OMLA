//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(KEYINPUT3), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n465), .A2(new_n466), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(new_n464), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  OAI22_X1  g051(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n468), .A2(new_n478), .A3(KEYINPUT64), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT64), .B1(new_n468), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g055(.A(G125), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G113), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n477), .B1(new_n485), .B2(G2105), .ZN(G160));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n465), .A2(G2105), .A3(new_n470), .A4(new_n471), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT68), .ZN(new_n491));
  INV_X1    g066(.A(new_n472), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n492), .A2(KEYINPUT67), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(KEYINPUT67), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G136), .ZN(new_n496));
  OAI221_X1 g071(.A(new_n488), .B1(new_n489), .B2(new_n491), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  NOR2_X1   g073(.A1(new_n466), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n490), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G126), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n465), .A2(new_n470), .A3(new_n471), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n504), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n479), .B2(new_n480), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  XOR2_X1   g087(.A(KEYINPUT5), .B(G543), .Z(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT69), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n523), .A2(new_n525), .B1(G651), .B2(new_n528), .ZN(G166));
  XNOR2_X1  g104(.A(KEYINPUT5), .B(G543), .ZN(new_n530));
  INV_X1    g105(.A(new_n516), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n520), .A2(G51), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(G168));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n513), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n540), .B1(new_n543), .B2(KEYINPUT70), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(KEYINPUT70), .B2(new_n543), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n517), .A2(G90), .B1(new_n520), .B2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(new_n520), .A2(G43), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n531), .A2(new_n530), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n540), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT72), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n520), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n517), .A2(G91), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n564), .B(new_n565), .C1(new_n540), .C2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n517), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n520), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n530), .A2(G61), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(new_n575), .B1(G73), .B2(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n530), .A2(KEYINPUT73), .A3(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n540), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n520), .A2(G48), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n551), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n520), .A2(G47), .ZN(new_n584));
  XOR2_X1   g159(.A(KEYINPUT74), .B(G85), .Z(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n551), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n540), .B2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n517), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n513), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G168), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  OAI21_X1  g182(.A(new_n602), .B1(new_n552), .B2(new_n554), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n598), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g186(.A(new_n495), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G135), .ZN(new_n613));
  OR2_X1    g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n614), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n491), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(G123), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT76), .B(G2096), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n468), .A2(new_n478), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT64), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n468), .A2(new_n478), .A3(KEYINPUT64), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n476), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n620), .A2(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT78), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  INV_X1    g224(.A(KEYINPUT18), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n630), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2096), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n666), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  AOI211_X1 g245(.A(new_n668), .B(new_n670), .C1(new_n663), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  NAND2_X1  g252(.A1(G166), .A2(G16), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G16), .B2(G22), .ZN(new_n679));
  INV_X1    g254(.A(G1971), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G6), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n582), .B2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT80), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(G23), .B(G288), .S(G16), .Z(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n679), .A2(new_n680), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n681), .A2(new_n687), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT34), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n682), .A2(G24), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G290), .B2(G16), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT79), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  OR2_X1    g272(.A1(G25), .A2(G29), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n700));
  INV_X1    g275(.A(G119), .ZN(new_n701));
  INV_X1    g276(.A(G131), .ZN(new_n702));
  OAI221_X1 g277(.A(new_n700), .B1(new_n701), .B2(new_n491), .C1(new_n495), .C2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n698), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT35), .B(G1991), .Z(new_n706));
  AOI21_X1  g281(.A(KEYINPUT81), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n705), .B2(new_n706), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n693), .A2(new_n697), .A3(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n709), .A2(KEYINPUT36), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n682), .A2(G20), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT23), .Z(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G299), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT92), .ZN(new_n714));
  INV_X1    g289(.A(G1956), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n704), .A2(G35), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G162), .B2(new_n704), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT29), .Z(new_n719));
  INV_X1    g294(.A(G2090), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT93), .Z(new_n722));
  NOR2_X1   g297(.A1(new_n709), .A2(KEYINPUT36), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n710), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G160), .A2(G29), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G34), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n725), .B1(G29), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2084), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT89), .Z(new_n731));
  INV_X1    g306(.A(G1961), .ZN(new_n732));
  NOR2_X1   g307(.A1(G171), .A2(new_n682), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G5), .B2(new_n682), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n731), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n704), .A2(G32), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT26), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n626), .A2(G105), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G129), .ZN(new_n742));
  INV_X1    g317(.A(G141), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n741), .B1(new_n742), .B2(new_n491), .C1(new_n495), .C2(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(KEYINPUT87), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(KEYINPUT87), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n745), .A2(KEYINPUT88), .A3(new_n746), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n736), .B1(new_n751), .B2(new_n704), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n735), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT90), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT90), .ZN(new_n757));
  NOR2_X1   g332(.A1(G4), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n599), .B2(G16), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1348), .Z(new_n760));
  INV_X1    g335(.A(KEYINPUT31), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(G11), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(G11), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(G28), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n704), .B1(new_n764), .B2(G28), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n762), .B(new_n763), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G168), .A2(new_n682), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n682), .B2(G21), .ZN(new_n769));
  INV_X1    g344(.A(G1966), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n760), .B(new_n771), .C1(new_n770), .C2(new_n769), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G19), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n555), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT82), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n618), .A2(G29), .B1(G1341), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n704), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n704), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n776), .B1(new_n732), .B2(new_n734), .C1(G2078), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(G2078), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n780), .B1(new_n729), .B2(new_n728), .C1(new_n775), .C2(G1341), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n772), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n719), .A2(new_n720), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(KEYINPUT91), .ZN(new_n784));
  INV_X1    g359(.A(G2072), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  INV_X1    g362(.A(G139), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n495), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT85), .Z(new_n790));
  AND2_X1   g365(.A1(new_n625), .A2(G127), .ZN(new_n791));
  AND2_X1   g366(.A1(G115), .A2(G2104), .ZN(new_n792));
  OAI21_X1  g367(.A(G2105), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n704), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n704), .B2(G33), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n782), .B(new_n784), .C1(new_n785), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n753), .A2(new_n754), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n617), .A2(G128), .ZN(new_n798));
  INV_X1    g373(.A(G140), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n466), .A2(G116), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n798), .B1(new_n495), .B2(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G29), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n704), .A2(G26), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT28), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT84), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT83), .B(G2067), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n807), .A2(new_n808), .B1(new_n795), .B2(new_n785), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n797), .B(new_n809), .C1(new_n807), .C2(new_n808), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n783), .A2(KEYINPUT91), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n796), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n724), .A2(new_n756), .A3(new_n757), .A4(new_n812), .ZN(G150));
  XOR2_X1   g388(.A(G150), .B(KEYINPUT94), .Z(G311));
  NAND2_X1  g389(.A1(G80), .A2(G543), .ZN(new_n815));
  INV_X1    g390(.A(G67), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n513), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n540), .B1(new_n817), .B2(KEYINPUT95), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(KEYINPUT95), .B2(new_n817), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n517), .A2(G93), .B1(new_n520), .B2(G55), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n555), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT96), .B1(new_n819), .B2(new_n820), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT38), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n599), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n831), .A2(new_n832), .A3(G860), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n821), .A2(G860), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n833), .A2(new_n835), .ZN(G145));
  NAND2_X1  g411(.A1(new_n790), .A2(new_n793), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n749), .B2(new_n750), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n802), .B(new_n511), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n747), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n842), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n840), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n612), .A2(G142), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT97), .Z(new_n848));
  OR2_X1    g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n617), .A2(G130), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n703), .B(KEYINPUT98), .ZN(new_n854));
  INV_X1    g429(.A(new_n628), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n855), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n852), .B1(new_n860), .B2(new_n856), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n846), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n843), .A2(new_n859), .A3(new_n861), .A4(new_n845), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n618), .B(G160), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G162), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(KEYINPUT100), .A3(new_n871), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT40), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT40), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(G395));
  NAND2_X1  g453(.A1(new_n821), .A2(new_n602), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n598), .B(G299), .Z(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n827), .B(new_n609), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n880), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n887), .B(KEYINPUT101), .C1(new_n888), .C2(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(KEYINPUT101), .B2(new_n887), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  XNOR2_X1  g466(.A(G290), .B(G303), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n582), .B(G288), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n892), .B(new_n893), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n891), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n879), .B1(new_n896), .B2(new_n602), .ZN(G295));
  OAI21_X1  g472(.A(new_n879), .B1(new_n896), .B2(new_n602), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n882), .B1(new_n900), .B2(new_n884), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n880), .A2(KEYINPUT103), .A3(new_n881), .ZN(new_n902));
  INV_X1    g477(.A(new_n827), .ZN(new_n903));
  XNOR2_X1  g478(.A(G301), .B(G168), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n825), .A2(new_n826), .A3(new_n904), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n901), .A2(new_n902), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n907), .B(KEYINPUT102), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n905), .A2(new_n888), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n909), .A2(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n895), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n906), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n917), .A2(new_n885), .B1(new_n908), .B2(new_n913), .ZN(new_n918));
  AOI21_X1  g493(.A(G37), .B1(new_n918), .B2(new_n894), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(KEYINPUT43), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n894), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n918), .A2(new_n894), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n899), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n916), .A2(new_n921), .A3(new_n919), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT105), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n920), .A2(new_n926), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT44), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n894), .B1(new_n911), .B2(new_n914), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n935), .A2(new_n924), .A3(KEYINPUT43), .ZN(new_n936));
  INV_X1    g511(.A(new_n925), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n921), .B1(new_n937), .B2(new_n919), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n899), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n932), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n931), .A2(new_n940), .ZN(G397));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n625), .A2(new_n508), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n943));
  INV_X1    g518(.A(G126), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n490), .A2(new_n944), .B1(new_n499), .B2(new_n500), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n942), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n466), .B1(new_n481), .B2(new_n484), .ZN(new_n948));
  INV_X1    g523(.A(G40), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n948), .A2(new_n477), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n951), .B(new_n942), .C1(new_n943), .C2(new_n945), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G8), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT49), .ZN(new_n956));
  INV_X1    g531(.A(G1981), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT109), .B1(new_n582), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  NOR4_X1   g534(.A1(new_n578), .A2(new_n581), .A3(new_n959), .A4(G1981), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n958), .A2(new_n960), .B1(new_n957), .B2(new_n582), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n956), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n961), .B2(new_n956), .ZN(new_n965));
  OAI221_X1 g540(.A(new_n955), .B1(new_n956), .B2(new_n961), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(G303), .A2(KEYINPUT107), .A3(KEYINPUT55), .A4(G8), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n968));
  INV_X1    g543(.A(G8), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(G166), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(G166), .A2(new_n969), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT107), .B1(new_n972), .B2(KEYINPUT55), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT108), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n970), .A4(new_n967), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT45), .B(new_n942), .C1(new_n943), .C2(new_n945), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n950), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n946), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n680), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n947), .A2(new_n987), .A3(new_n952), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n477), .A2(new_n949), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n485), .A2(G2105), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(KEYINPUT50), .B2(new_n946), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n986), .B1(G2090), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n974), .A2(new_n979), .A3(new_n994), .A4(G8), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n953), .B(G8), .C1(new_n996), .C2(G288), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT52), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n966), .A2(new_n995), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n988), .A2(new_n992), .A3(new_n729), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n947), .A2(new_n952), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n981), .B1(new_n1005), .B2(new_n983), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1004), .B1(new_n1006), .B2(G1966), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1007), .A2(G8), .A3(G168), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n951), .B1(new_n511), .B2(new_n942), .ZN(new_n1009));
  INV_X1    g584(.A(new_n952), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT50), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n950), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n987), .B1(new_n947), .B2(new_n952), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT113), .B1(new_n1014), .B2(new_n991), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n503), .B2(new_n510), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n987), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT114), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1013), .A2(new_n1015), .A3(new_n1020), .A4(new_n1017), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n720), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n969), .B1(new_n1022), .B2(new_n986), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n971), .A2(new_n973), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1003), .B(new_n1008), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT63), .ZN(new_n1029));
  AOI21_X1  g604(.A(G2090), .B1(new_n1018), .B2(KEYINPUT114), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1030), .A2(new_n1021), .B1(new_n680), .B2(new_n985), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1024), .B1(new_n1031), .B2(new_n969), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT115), .A3(new_n1003), .A4(new_n1008), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n995), .A2(KEYINPUT63), .A3(new_n1008), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1025), .B1(G8), .B2(new_n994), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n966), .A2(new_n1037), .A3(new_n1002), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n955), .B1(new_n956), .B2(new_n961), .ZN(new_n1039));
  INV_X1    g614(.A(new_n965), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(new_n963), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT111), .B1(new_n1041), .B2(new_n1001), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1036), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1045), .B(new_n1036), .C1(new_n1038), .C2(new_n1042), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1035), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1034), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT126), .ZN(new_n1049));
  INV_X1    g624(.A(G2078), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n984), .A2(new_n1050), .A3(new_n950), .A4(new_n980), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n993), .A2(new_n732), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n983), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1055), .A2(KEYINPUT121), .A3(new_n1050), .A4(new_n982), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT53), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT121), .B1(new_n1006), .B2(new_n1050), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1053), .B(new_n1054), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT45), .B1(new_n511), .B2(new_n942), .ZN(new_n1061));
  INV_X1    g636(.A(G125), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n623), .B2(new_n624), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT123), .B1(new_n1063), .B2(new_n483), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n481), .A2(new_n1065), .A3(new_n484), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(G2105), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n989), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT124), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n984), .A2(new_n1070), .A3(new_n989), .A4(new_n1067), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n980), .A2(KEYINPUT53), .A3(new_n1050), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1053), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1054), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n993), .A2(KEYINPUT122), .A3(new_n732), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G301), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1060), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(G171), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1054), .B(new_n1084), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(KEYINPUT54), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1079), .B2(G301), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n989), .B(new_n1067), .C1(new_n1016), .C2(KEYINPUT45), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1072), .B1(new_n1089), .B2(KEYINPUT124), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1090), .A2(new_n1071), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT122), .B1(new_n993), .B2(new_n732), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1076), .B(G1961), .C1(new_n988), .C2(new_n992), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1086), .A2(new_n1088), .A3(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1004), .B(G168), .C1(new_n1006), .C2(G1966), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G8), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1007), .A2(G286), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(G8), .A3(new_n1097), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1102), .B2(KEYINPUT51), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1083), .A2(new_n1096), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1032), .A2(new_n1003), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1049), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n966), .A2(new_n995), .A3(new_n1002), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1022), .A2(new_n986), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1108), .B1(new_n1110), .B2(new_n1024), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1094), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT125), .B1(new_n1094), .B2(G171), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1103), .B1(new_n1114), .B2(new_n1086), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1111), .A2(new_n1115), .A3(KEYINPUT126), .A4(new_n1083), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1348), .B1(new_n988), .B2(new_n992), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n953), .A2(G2067), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT118), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1125));
  OR3_X1    g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n598), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1018), .A2(new_n715), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n1129));
  OAI21_X1  g704(.A(G299), .B1(KEYINPUT117), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(KEYINPUT117), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n982), .A2(new_n984), .A3(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1128), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1127), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1132), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1128), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(G1341), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n953), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n985), .B2(G1996), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n555), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1125), .A2(new_n598), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1126), .A2(new_n1137), .A3(new_n1142), .A4(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1120), .A2(new_n599), .A3(new_n1123), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1141), .B1(new_n1136), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1107), .A2(new_n1116), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G288), .A2(G1976), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT112), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1041), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n958), .A2(new_n960), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n955), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n995), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1060), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n1169), .B2(new_n1111), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1048), .A2(new_n1159), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n984), .A2(new_n991), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n802), .B(G2067), .ZN(new_n1173));
  INV_X1    g748(.A(G1996), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n745), .B2(new_n746), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1173), .B(new_n1175), .C1(new_n751), .C2(new_n1174), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n703), .B(new_n706), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(G290), .B(G1986), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1172), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1171), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1172), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1182), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1184), .B1(new_n1178), .B2(new_n1172), .ZN(new_n1185));
  INV_X1    g760(.A(new_n706), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n703), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1176), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n802), .A2(G2067), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1182), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1172), .B1(new_n1173), .B2(new_n747), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT46), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT47), .Z(new_n1195));
  NOR3_X1   g770(.A1(new_n1185), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1181), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1181), .A2(KEYINPUT127), .A3(new_n1196), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g776(.A1(new_n874), .A2(new_n875), .ZN(new_n1203));
  OR3_X1    g777(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1204));
  AOI211_X1 g778(.A(G229), .B(new_n1204), .C1(new_n928), .C2(new_n929), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1203), .A2(new_n1205), .ZN(G225));
  INV_X1    g780(.A(G225), .ZN(G308));
endmodule


