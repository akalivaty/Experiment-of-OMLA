//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT27), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G190gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n205), .A2(new_n207), .A3(new_n209), .A4(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n206), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n202), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT69), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n218), .B(new_n202), .C1(new_n212), .C2(new_n215), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G190gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT27), .B(G183gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT28), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n224), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(G169gat), .ZN(new_n234));
  INV_X1    g033(.A(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT23), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT25), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT24), .B1(new_n206), .B2(new_n208), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n220), .A2(new_n206), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n235), .ZN(new_n248));
  NAND2_X1  g047(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n248), .A2(KEYINPUT23), .A3(new_n234), .A4(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n250), .A2(KEYINPUT65), .A3(new_n237), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT65), .B1(new_n250), .B2(new_n237), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n240), .A2(new_n242), .B1(new_n206), .B2(new_n208), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n246), .B1(new_n254), .B2(KEYINPUT25), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G127gat), .ZN(new_n257));
  INV_X1    g056(.A(G127gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G120gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(KEYINPUT1), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n262), .A2(new_n270), .A3(KEYINPUT70), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT70), .B1(new_n262), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n232), .A2(new_n255), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n273), .ZN(new_n275));
  INV_X1    g074(.A(new_n222), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n216), .B2(KEYINPUT69), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n230), .B1(new_n277), .B2(new_n219), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n234), .A2(KEYINPUT23), .ZN(new_n280));
  AND2_X1   g079(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n224), .B1(KEYINPUT23), .B2(new_n226), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n250), .A2(KEYINPUT65), .A3(new_n237), .ZN(new_n286));
  INV_X1    g085(.A(new_n253), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT25), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n245), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n275), .B1(new_n278), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G227gat), .ZN(new_n292));
  INV_X1    g091(.A(G233gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G15gat), .B(G43gat), .Z(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n274), .A2(new_n291), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT34), .B1(new_n302), .B2(new_n294), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n294), .B1(new_n274), .B2(new_n291), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT34), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n295), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n300), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n295), .B2(new_n296), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n304), .A2(new_n305), .ZN(new_n313));
  AOI211_X1 g112(.A(KEYINPUT34), .B(new_n294), .C1(new_n274), .C2(new_n291), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n307), .A2(new_n310), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n310), .B1(new_n307), .B2(new_n315), .ZN(new_n317));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT71), .B(G211gat), .Z(new_n322));
  AOI21_X1  g121(.A(KEYINPUT22), .B1(new_n322), .B2(G218gat), .ZN(new_n323));
  XOR2_X1   g122(.A(G197gat), .B(G204gat), .Z(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n326));
  INV_X1    g125(.A(new_n324), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT71), .B(G211gat), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n320), .B(new_n327), .C1(new_n330), .C2(KEYINPUT22), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(KEYINPUT72), .B(new_n321), .C1(new_n323), .C2(new_n324), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n342));
  INV_X1    g141(.A(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(G141gat), .ZN(new_n344));
  INV_X1    g143(.A(G141gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(G148gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n342), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n343), .B2(G141gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n343), .A2(G141gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n336), .B1(new_n339), .B2(KEYINPUT2), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n335), .B1(new_n356), .B2(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n332), .A2(new_n333), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n359), .B2(new_n335), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n341), .A2(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n319), .B(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n325), .B2(new_n331), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n356), .B1(new_n364), .B2(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n363), .B1(new_n366), .B2(new_n318), .ZN(new_n367));
  AOI211_X1 g166(.A(KEYINPUT80), .B(new_n319), .C1(new_n358), .C2(new_n365), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT31), .B(G50gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n376), .B2(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n377), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n362), .B(new_n379), .C1(new_n367), .C2(new_n368), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n316), .A2(new_n317), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(G226gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n293), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n232), .A2(new_n255), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n335), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n278), .B2(new_n290), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n391), .A3(new_n359), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT73), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n359), .B1(new_n389), .B2(new_n391), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n232), .A2(new_n255), .B1(new_n335), .B2(new_n388), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n278), .A2(new_n290), .A3(new_n387), .ZN(new_n398));
  OAI211_X1 g197(.A(KEYINPUT73), .B(new_n334), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT30), .B(new_n385), .C1(new_n396), .C2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n334), .B1(new_n397), .B2(new_n398), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n393), .A3(new_n392), .ZN(new_n403));
  INV_X1    g202(.A(new_n385), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n403), .B2(new_n399), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT74), .B1(new_n407), .B2(KEYINPUT30), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n385), .B1(new_n396), .B2(new_n400), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT74), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n406), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G1gat), .B(G29gat), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT0), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n418), .B(new_n361), .C1(new_n271), .C2(new_n272), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n262), .A2(new_n270), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT4), .B1(new_n356), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT78), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT78), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n424), .A3(new_n421), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n426));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT77), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n420), .B1(new_n361), .B2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n348), .A2(new_n429), .A3(new_n355), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n426), .B(new_n428), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n425), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n356), .A2(new_n420), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n361), .A2(new_n270), .A3(new_n262), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n428), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n426), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(KEYINPUT4), .B(new_n361), .C1(new_n271), .C2(new_n272), .ZN(new_n440));
  INV_X1    g239(.A(new_n436), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(KEYINPUT4), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n417), .B1(new_n434), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(KEYINPUT6), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n434), .A2(new_n444), .A3(new_n417), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n444), .ZN(new_n450));
  INV_X1    g249(.A(new_n417), .ZN(new_n451));
  AND4_X1   g250(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT6), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n445), .B2(KEYINPUT6), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n445), .A2(new_n449), .A3(KEYINPUT6), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT85), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n448), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT35), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n382), .A2(new_n413), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n452), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n448), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n382), .A2(new_n413), .A3(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n462), .A2(KEYINPUT87), .B1(new_n465), .B2(KEYINPUT35), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n454), .B1(new_n452), .B2(new_n453), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n457), .A2(KEYINPUT85), .A3(new_n458), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n467), .A2(new_n468), .B1(new_n447), .B2(new_n446), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(KEYINPUT35), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n382), .A4(new_n413), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n435), .A2(new_n436), .A3(new_n428), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT39), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n430), .A2(new_n431), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n423), .A2(new_n475), .A3(new_n425), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n476), .B2(new_n438), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT82), .B(KEYINPUT39), .Z(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n438), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n478), .A2(KEYINPUT40), .A3(new_n417), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n445), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT83), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n417), .A3(new_n480), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n480), .A2(new_n417), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n484), .B(new_n486), .C1(new_n489), .C2(new_n477), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n483), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n412), .A2(new_n408), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n403), .A2(new_n399), .A3(new_n404), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(KEYINPUT30), .B2(new_n407), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n381), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n404), .A2(KEYINPUT37), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n405), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n403), .A2(KEYINPUT37), .A3(new_n399), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT38), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(KEYINPUT86), .A3(KEYINPUT38), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT84), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n389), .A2(new_n391), .A3(new_n505), .A4(new_n359), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n506), .A2(KEYINPUT37), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n402), .A2(KEYINPUT84), .A3(new_n392), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT38), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n407), .B1(new_n498), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n503), .A2(new_n469), .A3(new_n504), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n316), .A2(new_n317), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT36), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n316), .B2(new_n317), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n407), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n464), .B(new_n494), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n514), .A2(new_n516), .B1(new_n519), .B2(new_n381), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n466), .A2(new_n472), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G197gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT11), .B(G169gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT88), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528));
  INV_X1    g327(.A(G29gat), .ZN(new_n529));
  INV_X1    g328(.A(G36gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT14), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(KEYINPUT14), .ZN(new_n534));
  NAND2_X1  g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n536), .A2(KEYINPUT90), .B1(KEYINPUT15), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(KEYINPUT15), .B2(new_n537), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT17), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(G1gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(G1gat), .B2(new_n545), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n540), .A2(new_n552), .A3(new_n541), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n543), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n542), .A2(new_n551), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n554), .A2(new_n556), .A3(KEYINPUT18), .A4(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(KEYINPUT13), .Z(new_n559));
  AND2_X1   g358(.A1(new_n542), .A2(new_n551), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n555), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n562), .A2(new_n563), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n527), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n558), .A2(new_n561), .A3(new_n526), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n565), .A2(KEYINPUT93), .A3(new_n566), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n521), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G64gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G57gat), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT94), .B(G57gat), .Z(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  OR2_X1    g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n583), .B(new_n584), .C1(new_n588), .C2(new_n585), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT95), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n551), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n591), .A2(new_n592), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT20), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n602), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n601), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n605), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n606), .B2(new_n610), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n598), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n611), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n606), .A2(new_n610), .A3(new_n612), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n597), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n542), .ZN(new_n621));
  NAND2_X1  g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT7), .ZN(new_n623));
  NAND2_X1  g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT8), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n623), .B(new_n625), .C1(G85gat), .C2(G92gat), .ZN(new_n626));
  XOR2_X1   g425(.A(G99gat), .B(G106gat), .Z(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(KEYINPUT98), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n621), .A2(new_n633), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n633), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n543), .A2(new_n553), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G190gat), .B(G218gat), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G134gat), .B(G162gat), .Z(new_n642));
  NOR2_X1   g441(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT99), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n641), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(G230gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n293), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n593), .A2(new_n633), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n626), .A2(KEYINPUT100), .A3(new_n627), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n628), .A2(new_n659), .A3(new_n630), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n591), .A2(new_n592), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n636), .A2(new_n593), .A3(new_n663), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n656), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n657), .A2(new_n656), .A3(new_n661), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n657), .A2(KEYINPUT101), .A3(new_n661), .A4(new_n656), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n654), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT10), .B1(new_n657), .B2(new_n661), .ZN(new_n674));
  OAI22_X1  g473(.A1(new_n674), .A2(new_n665), .B1(new_n655), .B2(new_n293), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n675), .A2(new_n653), .A3(new_n671), .A4(new_n670), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n620), .A2(new_n650), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n578), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n464), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g484(.A(new_n544), .B1(new_n682), .B2(new_n495), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n681), .A2(new_n413), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(KEYINPUT42), .B2(new_n688), .ZN(G1325gat));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n514), .A2(new_n691), .A3(new_n516), .ZN(new_n692));
  INV_X1    g491(.A(new_n317), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n307), .A2(new_n310), .A3(new_n315), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT36), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n316), .A2(new_n317), .A3(new_n515), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT102), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n681), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n513), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n681), .B2(new_n701), .ZN(G1326gat));
  NAND2_X1  g501(.A1(new_n682), .A2(new_n381), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT103), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n521), .B2(new_n650), .ZN(new_n707));
  INV_X1    g506(.A(new_n381), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n513), .A2(new_n708), .A3(new_n492), .A4(new_n494), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n460), .A2(new_n461), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT87), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n382), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT35), .B1(new_n712), .B2(new_n519), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n472), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n467), .A2(new_n468), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n510), .A3(new_n448), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT86), .B1(new_n500), .B2(KEYINPUT38), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT38), .ZN(new_n718));
  AOI211_X1 g517(.A(new_n502), .B(new_n718), .C1(new_n498), .C2(new_n499), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n481), .A2(new_n482), .ZN(new_n721));
  INV_X1    g520(.A(new_n490), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n487), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n708), .B1(new_n413), .B2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n692), .B(new_n697), .C1(new_n720), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n519), .A2(new_n381), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT104), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n519), .A2(new_n728), .A3(new_n381), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n714), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n650), .A2(KEYINPUT44), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n707), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n620), .A2(new_n577), .A3(new_n677), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n739), .B2(new_n464), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n521), .A2(new_n650), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n738), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n529), .A3(new_n683), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1328gat));
  OAI21_X1  g546(.A(G36gat), .B1(new_n739), .B2(new_n413), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n649), .A2(new_n530), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n620), .A2(new_n749), .A3(new_n677), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n578), .A2(new_n495), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n748), .A2(new_n753), .ZN(G1329gat));
  OAI21_X1  g553(.A(G43gat), .B1(new_n739), .B2(new_n698), .ZN(new_n755));
  INV_X1    g554(.A(G43gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n742), .A2(new_n756), .A3(new_n513), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(KEYINPUT108), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1330gat));
  NAND2_X1  g561(.A1(new_n381), .A2(G50gat), .ZN(new_n763));
  INV_X1    g562(.A(new_n742), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n708), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n739), .A2(new_n763), .B1(new_n765), .B2(G50gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g566(.A(new_n620), .ZN(new_n768));
  NOR4_X1   g567(.A1(new_n768), .A2(new_n576), .A3(new_n649), .A4(new_n678), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n731), .A2(KEYINPUT109), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT109), .B1(new_n731), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n683), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT110), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(new_n581), .ZN(G1332gat));
  INV_X1    g574(.A(new_n772), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n413), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT111), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1333gat));
  INV_X1    g580(.A(G71gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n776), .B2(new_n700), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n698), .A2(new_n782), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n772), .B2(new_n785), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n772), .A2(new_n784), .A3(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n381), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT113), .B(G78gat), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n620), .A2(new_n576), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n678), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n737), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n464), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n794), .A2(new_n650), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n798), .A2(new_n731), .A3(KEYINPUT51), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n798), .B2(new_n731), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n678), .A2(G85gat), .A3(new_n464), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT114), .Z(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n797), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT115), .ZN(G1336gat));
  NOR2_X1   g605(.A1(new_n413), .A2(G92gat), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n677), .B(new_n807), .C1(new_n799), .C2(new_n800), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n808), .A2(KEYINPUT118), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n495), .B(new_n795), .C1(new_n735), .C2(new_n736), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G92gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(KEYINPUT118), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n809), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n808), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n811), .B2(KEYINPUT116), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n810), .A2(new_n817), .A3(G92gat), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT117), .B(new_n812), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n811), .A2(KEYINPUT116), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n808), .A3(new_n818), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n822), .B2(KEYINPUT52), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n814), .B1(new_n819), .B2(new_n823), .ZN(G1337gat));
  INV_X1    g623(.A(new_n796), .ZN(new_n825));
  INV_X1    g624(.A(G99gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n698), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n801), .A2(new_n513), .A3(new_n677), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n825), .A2(new_n827), .B1(new_n826), .B2(new_n828), .ZN(G1338gat));
  INV_X1    g628(.A(G106gat), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n708), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n801), .A2(new_n381), .A3(new_n677), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n825), .A2(new_n831), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n653), .B1(new_n667), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n664), .A2(new_n666), .A3(new_n656), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n675), .A3(KEYINPUT54), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(KEYINPUT55), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n676), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT119), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n842), .A3(new_n676), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  INV_X1    g643(.A(new_n838), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n654), .B1(new_n675), .B2(KEYINPUT54), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n841), .A2(new_n576), .A3(new_n843), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n557), .B1(new_n554), .B2(new_n556), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n560), .A2(new_n555), .A3(new_n559), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n525), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT120), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n575), .A3(new_n677), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n649), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n841), .A2(new_n843), .A3(new_n847), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n649), .A2(new_n575), .A3(new_n852), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n768), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n679), .A2(new_n576), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n464), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n709), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n576), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n381), .B1(new_n858), .B2(new_n860), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n495), .A2(new_n464), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n866), .A2(new_n513), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n577), .A2(new_n265), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(G1340gat));
  AOI21_X1  g669(.A(G120gat), .B1(new_n864), .B2(new_n677), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n678), .A2(new_n263), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n868), .B2(new_n872), .ZN(G1341gat));
  NOR3_X1   g672(.A1(new_n863), .A2(G127gat), .A3(new_n768), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n620), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(G127gat), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT121), .Z(G1342gat));
  NOR3_X1   g676(.A1(new_n863), .A2(G134gat), .A3(new_n650), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n256), .B1(new_n868), .B2(new_n649), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(KEYINPUT56), .B2(new_n879), .ZN(G1343gat));
  AND3_X1   g682(.A1(new_n852), .A2(new_n575), .A3(new_n677), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n847), .A2(new_n676), .A3(new_n839), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n576), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT122), .B1(new_n886), .B2(new_n649), .ZN(new_n887));
  INV_X1    g686(.A(new_n857), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n847), .A2(new_n676), .A3(new_n839), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n853), .B1(new_n577), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n650), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n859), .B1(new_n893), .B2(new_n768), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n708), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n698), .A2(new_n867), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n708), .B1(new_n858), .B2(new_n860), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n899), .A3(new_n576), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G141gat), .ZN(new_n901));
  INV_X1    g700(.A(new_n698), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n708), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n861), .A2(new_n413), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n577), .A2(G141gat), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT58), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n895), .B2(new_n899), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n899), .A3(new_n908), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n576), .A3(new_n911), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n912), .A2(G141gat), .B1(new_n904), .B2(new_n905), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(G1344gat));
  NAND2_X1  g714(.A1(new_n343), .A2(KEYINPUT59), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n904), .B2(new_n677), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n895), .A2(new_n899), .A3(new_n908), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n909), .A3(new_n678), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n897), .A2(new_n898), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n890), .A2(new_n650), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n620), .B1(new_n888), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n898), .B(new_n381), .C1(new_n922), .C2(new_n859), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n677), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n698), .A2(KEYINPUT59), .A3(new_n867), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n919), .A2(KEYINPUT59), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n917), .B1(new_n927), .B2(G148gat), .ZN(G1345gat));
  AND2_X1   g727(.A1(new_n904), .A2(new_n620), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n911), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n620), .A2(G155gat), .ZN(new_n931));
  OAI221_X1 g730(.A(KEYINPUT124), .B1(G155gat), .B2(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n918), .A2(new_n909), .A3(new_n931), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n929), .A2(G155gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n936), .ZN(G1346gat));
  AOI21_X1  g736(.A(G162gat), .B1(new_n904), .B2(new_n649), .ZN(new_n938));
  INV_X1    g737(.A(new_n930), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n649), .A2(G162gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n413), .A2(new_n683), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(new_n700), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n866), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n945), .A2(new_n234), .A3(new_n577), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n683), .B1(new_n858), .B2(new_n860), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(new_n382), .A3(new_n495), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n576), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n234), .B2(new_n949), .ZN(G1348gat));
  AOI21_X1  g749(.A(G176gat), .B1(new_n948), .B2(new_n677), .ZN(new_n951));
  INV_X1    g750(.A(new_n945), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n678), .B1(new_n248), .B2(new_n249), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT125), .Z(G1349gat));
  OAI21_X1  g754(.A(G183gat), .B1(new_n945), .B2(new_n768), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n620), .A2(new_n221), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n948), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n948), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g761(.A1(new_n948), .A2(new_n220), .A3(new_n649), .ZN(new_n963));
  OAI21_X1  g762(.A(G190gat), .B1(new_n945), .B2(new_n650), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1351gat));
  NOR2_X1   g766(.A1(new_n902), .A2(new_n943), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT127), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n924), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n576), .A2(G197gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n947), .A2(new_n495), .A3(new_n903), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n973), .A2(new_n577), .ZN(new_n974));
  OAI22_X1  g773(.A1(new_n971), .A2(new_n972), .B1(G197gat), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(G1352gat));
  OAI21_X1  g775(.A(G204gat), .B1(new_n925), .B2(new_n969), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n973), .A2(G204gat), .A3(new_n678), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(G1353gat));
  NAND3_X1  g781(.A1(new_n924), .A2(new_n620), .A3(new_n968), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n620), .A2(new_n328), .ZN(new_n986));
  OAI22_X1  g785(.A1(new_n984), .A2(new_n985), .B1(new_n973), .B2(new_n986), .ZN(G1354gat));
  OAI21_X1  g786(.A(new_n329), .B1(new_n973), .B2(new_n650), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n649), .A2(G218gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n971), .B2(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(G1355gat));
endmodule


