//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT72), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT72), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G237), .ZN(new_n191));
  AOI21_X1  g005(.A(G953), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n192), .A2(G214), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n193), .B1(new_n194), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(KEYINPUT17), .A3(G131), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n210), .A3(KEYINPUT16), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(G146), .A3(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT91), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n218), .A3(new_n215), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n205), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT92), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n205), .A2(new_n217), .A3(new_n222), .A4(new_n219), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n204), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n200), .A2(KEYINPUT18), .A3(G131), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n207), .A2(new_n210), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n213), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n226), .B(KEYINPUT88), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n213), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(new_n201), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n225), .B(new_n229), .C1(new_n200), .C2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G113), .B(G122), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT90), .B(G104), .ZN(new_n234));
  XOR2_X1   g048(.A(new_n233), .B(new_n234), .Z(new_n235));
  NAND3_X1  g049(.A1(new_n224), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT19), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n238), .A2(KEYINPUT89), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n226), .A2(KEYINPUT89), .A3(new_n237), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n239), .B(new_n240), .C1(new_n237), .C2(new_n228), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n215), .B1(new_n241), .B2(G146), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n232), .B1(new_n242), .B2(new_n202), .ZN(new_n243));
  INV_X1    g057(.A(new_n235), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(G475), .A2(G902), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n187), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  AOI211_X1 g063(.A(KEYINPUT20), .B(new_n249), .C1(new_n236), .C2(new_n245), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n235), .B1(new_n224), .B2(new_n232), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(G902), .B1(new_n252), .B2(new_n236), .ZN(new_n253));
  INV_X1    g067(.A(G475), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n248), .A2(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(G234), .A2(G237), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(G952), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(G902), .A3(G953), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT21), .B(G898), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G478), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT15), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT64), .B(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G128), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G143), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G122), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G116), .ZN(new_n273));
  INV_X1    g087(.A(G116), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G122), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n275), .A3(G107), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n275), .ZN(new_n277));
  INV_X1    g091(.A(G107), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n267), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT93), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n266), .A2(KEYINPUT13), .A3(G128), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n266), .A2(G128), .B1(KEYINPUT13), .B2(new_n270), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n268), .B1(new_n286), .B2(KEYINPUT93), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n280), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n278), .B1(new_n273), .B2(KEYINPUT14), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n290), .A2(new_n277), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n277), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n267), .A2(new_n270), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G134), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n271), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  INV_X1    g112(.A(G217), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n298), .A2(new_n299), .A3(G953), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n289), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n300), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n288), .B2(new_n296), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT94), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n306), .B(G902), .C1(new_n301), .C2(new_n303), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n265), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI22_X1  g122(.A1(new_n304), .A2(KEYINPUT94), .B1(KEYINPUT15), .B2(new_n264), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n255), .A2(new_n263), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G210), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT87), .ZN(new_n314));
  OR2_X1    g128(.A1(KEYINPUT69), .A2(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT69), .A2(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(G116), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n274), .A2(G119), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(G113), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT86), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT2), .ZN(new_n323));
  INV_X1    g137(.A(G113), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT68), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(KEYINPUT2), .B2(G113), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n325), .A2(new_n327), .B1(KEYINPUT2), .B2(G113), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n317), .A3(new_n318), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n317), .A2(new_n318), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n328), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(KEYINPUT81), .A2(G104), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT81), .A2(G104), .ZN(new_n336));
  AOI21_X1  g150(.A(G107), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT82), .B1(new_n278), .B2(G104), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n339), .B(G101), .C1(new_n337), .C2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n335), .B(new_n336), .C1(KEYINPUT3), .C2(G107), .ZN(new_n342));
  AND2_X1   g156(.A1(KEYINPUT3), .A2(G107), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT3), .A2(G107), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(G104), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT86), .B1(new_n320), .B2(new_n321), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n322), .A2(new_n334), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G110), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT8), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n321), .B1(KEYINPUT5), .B2(new_n331), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n333), .B2(new_n330), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n350), .B(new_n352), .C1(new_n354), .C2(new_n348), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n213), .A2(G143), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n199), .B2(new_n213), .ZN(new_n357));
  AND2_X1   g171(.A1(KEYINPUT0), .A2(G128), .ZN(new_n358));
  NOR2_X1   g172(.A1(KEYINPUT0), .A2(G128), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT65), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n196), .A2(new_n198), .A3(G146), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n213), .A2(G143), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n358), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT65), .ZN(new_n366));
  AOI21_X1  g180(.A(G146), .B1(new_n196), .B2(new_n198), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n366), .B(new_n360), .C1(new_n367), .C2(new_n356), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G125), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n363), .A2(new_n371), .A3(G128), .A4(new_n364), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n269), .B1(new_n364), .B2(KEYINPUT1), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n357), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n209), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n257), .A2(G224), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n370), .A2(KEYINPUT7), .A3(new_n376), .A4(new_n379), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n355), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n346), .B1(new_n342), .B2(new_n345), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT4), .A3(new_n347), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n331), .A2(new_n328), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n330), .B2(new_n333), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n322), .A2(new_n334), .A3(new_n349), .ZN(new_n392));
  OAI221_X1 g206(.A(new_n351), .B1(new_n389), .B2(new_n391), .C1(new_n392), .C2(new_n348), .ZN(new_n393));
  AOI21_X1  g207(.A(G902), .B1(new_n383), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n351), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n392), .A2(new_n348), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n389), .A2(new_n391), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n393), .A3(KEYINPUT6), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(new_n395), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n377), .B(new_n380), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n314), .B1(new_n394), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n394), .A2(new_n403), .A3(new_n314), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G214), .B1(G237), .B2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n257), .A2(G227), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT11), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n268), .B2(G137), .ZN(new_n416));
  INV_X1    g230(.A(G137), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT11), .A3(G134), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n268), .A2(G137), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G131), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n416), .A2(new_n418), .A3(new_n201), .A4(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n372), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n363), .A2(new_n364), .ZN(new_n425));
  OAI21_X1  g239(.A(G128), .B1(new_n367), .B2(new_n371), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(new_n348), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n374), .B1(new_n341), .B2(new_n347), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(KEYINPUT12), .B(new_n423), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n375), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n348), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n435), .B1(new_n427), .B2(new_n348), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n368), .A2(new_n365), .ZN(new_n440));
  INV_X1    g254(.A(new_n356), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(new_n266), .B2(G146), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n366), .B1(new_n442), .B2(new_n360), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n386), .A3(new_n388), .ZN(new_n445));
  INV_X1    g259(.A(new_n423), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n438), .A2(new_n439), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n414), .B1(new_n434), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n426), .A2(new_n425), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n347), .B(new_n341), .C1(new_n449), .C2(new_n424), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n435), .A2(new_n450), .B1(new_n436), .B2(new_n437), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n446), .B1(new_n451), .B2(new_n445), .ZN(new_n452));
  INV_X1    g266(.A(new_n447), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n452), .A2(new_n453), .A3(new_n413), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT83), .B1(new_n448), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n452), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n447), .A2(new_n414), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n453), .B1(new_n433), .B2(new_n432), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n414), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n461), .A3(G469), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  INV_X1    g277(.A(G902), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n457), .A2(new_n434), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n413), .B1(new_n452), .B2(new_n453), .ZN(new_n467));
  AOI21_X1  g281(.A(G902), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n465), .B1(new_n468), .B2(new_n463), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT84), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n473));
  INV_X1    g287(.A(new_n471), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n473), .B(new_n474), .C1(new_n462), .C2(new_n469), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n311), .B(new_n410), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT25), .ZN(new_n478));
  NOR2_X1   g292(.A1(G119), .A2(G128), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n315), .A2(new_n316), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(G128), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT23), .ZN(new_n482));
  INV_X1    g296(.A(G110), .ZN(new_n483));
  AOI21_X1  g297(.A(G128), .B1(new_n315), .B2(new_n316), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n484), .A2(KEYINPUT23), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT78), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT24), .B(G110), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n486), .B2(new_n489), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n215), .B(new_n227), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT79), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n216), .B1(new_n481), .B2(new_n488), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n483), .B1(new_n482), .B2(new_n485), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n215), .A2(new_n227), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n486), .A2(new_n489), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n502), .B2(new_n490), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT79), .B1(new_n503), .B2(new_n497), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT22), .B(G137), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT80), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n499), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n493), .A2(new_n498), .A3(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n478), .B1(new_n512), .B2(G902), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n510), .A2(KEYINPUT25), .A3(new_n464), .A4(new_n511), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n299), .B1(G234), .B2(new_n464), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT77), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n192), .A2(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n268), .A2(G137), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n417), .A2(G134), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n422), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n374), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n362), .A2(new_n365), .A3(new_n368), .A4(new_n423), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n391), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT66), .B1(new_n440), .B2(new_n443), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT66), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n362), .A2(new_n539), .A3(new_n365), .A4(new_n368), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n540), .A3(new_n423), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n532), .A2(KEYINPUT67), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n422), .A2(new_n531), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n374), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n534), .A2(KEYINPUT30), .A3(new_n533), .ZN(new_n550));
  INV_X1    g364(.A(new_n391), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT71), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT30), .B1(new_n541), .B2(new_n546), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n551), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n537), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT31), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n542), .A2(new_n374), .A3(new_n545), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n446), .B1(new_n369), .B2(KEYINPUT66), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n562), .B2(new_n540), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n552), .B(KEYINPUT71), .C1(new_n563), .C2(KEYINPUT30), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n537), .ZN(new_n567));
  INV_X1    g381(.A(new_n528), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n535), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n391), .A2(KEYINPUT28), .A3(new_n533), .A4(new_n534), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n391), .B1(new_n541), .B2(new_n546), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT74), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT74), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n576), .B(new_n568), .C1(new_n572), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n559), .A2(new_n567), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(G472), .A2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT32), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n523), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI211_X1 g397(.A(KEYINPUT75), .B(KEYINPUT32), .C1(new_n579), .C2(new_n580), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G472), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n572), .A2(new_n573), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT29), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n568), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n534), .A2(new_n533), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n551), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n569), .B1(new_n591), .B2(new_n535), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT76), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n570), .A2(KEYINPUT76), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n594), .B(KEYINPUT29), .C1(new_n592), .C2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n589), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n565), .A2(new_n588), .A3(new_n535), .A4(new_n568), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n586), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n580), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n566), .B1(new_n565), .B2(new_n537), .ZN(new_n601));
  AOI211_X1 g415(.A(KEYINPUT31), .B(new_n536), .C1(new_n560), .C2(new_n564), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n603), .B2(new_n578), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n599), .B1(new_n604), .B2(KEYINPUT32), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n522), .B1(new_n585), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT75), .B1(new_n604), .B2(KEYINPUT32), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n581), .A2(new_n523), .A3(new_n582), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n522), .A2(new_n607), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n477), .B(new_n521), .C1(new_n606), .C2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  INV_X1    g425(.A(new_n472), .ZN(new_n612));
  INV_X1    g426(.A(new_n475), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n579), .A2(new_n464), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G472), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n581), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n521), .A3(new_n618), .ZN(new_n619));
  OR3_X1    g433(.A1(new_n304), .A2(KEYINPUT98), .A3(G478), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT98), .B1(new_n304), .B2(G478), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT33), .B1(new_n300), .B2(KEYINPUT96), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n301), .B2(new_n303), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n301), .A2(new_n303), .A3(new_n624), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n264), .A2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n622), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n255), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n394), .A2(new_n403), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n312), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n394), .A2(new_n403), .A3(new_n313), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n408), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT95), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT95), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n635), .A2(new_n639), .A3(new_n408), .A4(new_n636), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR4_X1   g455(.A1(new_n619), .A2(new_n263), .A3(new_n633), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT34), .B(G104), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(new_n310), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n255), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n263), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n619), .A2(new_n641), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND2_X1  g465(.A1(new_n499), .A2(new_n504), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT36), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n508), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT99), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n654), .B(KEYINPUT99), .Z(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n504), .A3(new_n499), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n656), .A2(new_n518), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n517), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n614), .A2(new_n311), .A3(new_n410), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n617), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT37), .B(G110), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  AND2_X1   g480(.A1(new_n661), .A2(new_n517), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n641), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n258), .B(KEYINPUT101), .Z(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n261), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n646), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n612), .B2(new_n613), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n668), .B(new_n675), .C1(new_n606), .C2(new_n609), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n672), .B(new_n678), .Z(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n472), .B2(new_n475), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n565), .A2(new_n535), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n528), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n591), .A2(new_n535), .ZN(new_n684));
  AOI21_X1  g498(.A(G902), .B1(new_n684), .B2(new_n568), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n586), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n604), .B2(KEYINPUT32), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n585), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT40), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n689), .B(new_n679), .C1(new_n472), .C2(new_n475), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n407), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n405), .A2(KEYINPUT38), .A3(new_n406), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n255), .A2(new_n310), .A3(new_n408), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n694), .A2(new_n662), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n681), .A2(new_n688), .A3(new_n690), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n696), .A2(new_n690), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(KEYINPUT103), .A3(new_n688), .A4(new_n681), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n266), .ZN(G45));
  NAND3_X1  g517(.A1(new_n255), .A2(new_n632), .A3(new_n673), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n612), .B2(new_n613), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n668), .B(new_n705), .C1(new_n606), .C2(new_n609), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  OR2_X1    g521(.A1(new_n468), .A2(new_n463), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n468), .A2(new_n463), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n471), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n638), .A3(new_n640), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n712), .A2(new_n263), .A3(new_n633), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n521), .B(new_n713), .C1(new_n606), .C2(new_n609), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT41), .B(G113), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT104), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n714), .B(new_n716), .ZN(G15));
  NOR2_X1   g531(.A1(new_n712), .A2(new_n648), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n521), .B(new_n718), .C1(new_n606), .C2(new_n609), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  INV_X1    g534(.A(new_n311), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n712), .A2(new_n721), .A3(new_n667), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n606), .B2(new_n609), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND4_X1  g538(.A1(new_n638), .A2(new_n255), .A3(new_n310), .A4(new_n640), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n263), .A3(new_n710), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n615), .A2(KEYINPUT106), .A3(G472), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n594), .B(new_n568), .C1(new_n592), .C2(new_n595), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n559), .A2(new_n567), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n580), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT105), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n732), .A3(new_n580), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT106), .B1(new_n615), .B2(G472), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n726), .A2(new_n521), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  INV_X1    g552(.A(new_n733), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n732), .B1(new_n729), .B2(new_n580), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n616), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n743), .A3(new_n662), .A4(new_n727), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n704), .A3(new_n712), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n209), .ZN(G27));
  NAND3_X1  g560(.A1(new_n607), .A2(new_n605), .A3(new_n608), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT77), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n585), .A2(new_n522), .A3(new_n605), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n704), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n465), .B(KEYINPUT107), .Z(new_n752));
  OAI21_X1  g566(.A(new_n458), .B1(new_n460), .B2(new_n414), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n709), .B(new_n752), .C1(new_n463), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n471), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n405), .A2(new_n408), .A3(new_n406), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n750), .A2(new_n521), .A3(new_n751), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n581), .A2(new_n582), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n605), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n751), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n766), .A3(new_n767), .A4(new_n521), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n521), .B1(new_n762), .B2(new_n763), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT109), .B1(new_n769), .B2(new_n765), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n758), .A2(new_n759), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT110), .B(G131), .Z(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G33));
  INV_X1    g587(.A(new_n674), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n750), .A2(new_n521), .A3(new_n774), .A4(new_n757), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n626), .A2(new_n627), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT97), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n628), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n780), .A2(new_n781), .B1(new_n621), .B2(new_n620), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT43), .B1(new_n255), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n248), .ZN(new_n784));
  INV_X1    g598(.A(new_n250), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  INV_X1    g601(.A(new_n236), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n464), .B1(new_n788), .B2(new_n251), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(G475), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n786), .A2(new_n632), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n662), .A2(new_n783), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n777), .B1(new_n792), .B2(new_n618), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n783), .A2(new_n791), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(KEYINPUT44), .A3(new_n617), .A4(new_n662), .ZN(new_n795));
  INV_X1    g609(.A(new_n406), .ZN(new_n796));
  INV_X1    g610(.A(new_n408), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n404), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n455), .B2(new_n461), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n803));
  OAI21_X1  g617(.A(G469), .B1(new_n753), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n752), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT46), .B(new_n752), .C1(new_n802), .C2(new_n804), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n709), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n471), .A3(new_n679), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n800), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NOR3_X1   g626(.A1(new_n521), .A2(new_n704), .A3(new_n756), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n809), .A2(KEYINPUT47), .A3(new_n471), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT47), .B1(new_n809), .B2(new_n471), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT111), .B1(new_n816), .B2(new_n750), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n809), .A2(new_n471), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT47), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n809), .A2(KEYINPUT47), .A3(new_n471), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n606), .A2(new_n609), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n813), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  XNOR2_X1  g641(.A(new_n468), .B(new_n463), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT49), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT49), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n474), .A2(new_n797), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n832), .A2(new_n255), .A3(new_n782), .ZN(new_n833));
  INV_X1    g647(.A(new_n688), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n521), .A4(new_n694), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n662), .B1(new_n472), .B2(new_n475), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n784), .A2(new_n785), .B1(G475), .B2(new_n789), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n308), .A2(new_n309), .A3(new_n673), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n798), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n840), .B(new_n790), .C1(new_n248), .C2(new_n250), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT114), .B1(new_n842), .B2(new_n756), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n837), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n734), .A2(new_n667), .A3(new_n704), .A4(new_n735), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n750), .A2(new_n844), .B1(new_n845), .B2(new_n757), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n775), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n714), .A2(new_n719), .A3(new_n723), .A4(new_n737), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n758), .A2(new_n759), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n768), .A2(new_n770), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n409), .A2(new_n633), .A3(new_n263), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n614), .A2(new_n521), .A3(new_n618), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n610), .A2(KEYINPUT112), .A3(new_n854), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n648), .A2(KEYINPUT113), .A3(new_n409), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT113), .B1(new_n648), .B2(new_n409), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n858), .A2(new_n619), .B1(new_n663), .B2(new_n617), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n610), .A2(new_n854), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n849), .A2(new_n852), .A3(new_n855), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n641), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n845), .A2(new_n864), .A3(new_n711), .ZN(new_n865));
  INV_X1    g679(.A(new_n725), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n662), .A2(new_n755), .A3(new_n672), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n688), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n676), .A2(new_n706), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT52), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n836), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n869), .B(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n862), .A2(new_n855), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n771), .A2(new_n847), .A3(new_n848), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n864), .A2(new_n662), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n748), .B2(new_n749), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n745), .B1(new_n878), .B2(new_n675), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n836), .B1(new_n880), .B2(KEYINPUT52), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n871), .A2(new_n872), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n836), .B1(new_n879), .B2(new_n873), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n872), .B1(new_n871), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n710), .A2(new_n756), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n794), .A2(new_n670), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n769), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT48), .ZN(new_n890));
  INV_X1    g704(.A(G952), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(G953), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n520), .A2(new_n258), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n585), .A3(new_n687), .A4(new_n887), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n736), .A2(new_n521), .A3(new_n670), .A4(new_n794), .ZN(new_n895));
  OAI221_X1 g709(.A(new_n892), .B1(new_n894), .B2(new_n633), .C1(new_n895), .C2(new_n712), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n783), .A2(new_n791), .A3(new_n670), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n897), .A2(new_n734), .A3(new_n520), .A4(new_n735), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n828), .A2(new_n471), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n798), .B(new_n898), .C1(new_n822), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NOR4_X1   g715(.A1(new_n520), .A2(new_n258), .A3(new_n710), .A4(new_n756), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n255), .A2(new_n632), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n834), .A2(new_n901), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n888), .A2(new_n744), .ZN(new_n905));
  INV_X1    g719(.A(new_n903), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT117), .B1(new_n894), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n900), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n910));
  NOR2_X1   g724(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n694), .A2(new_n797), .A3(new_n711), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n895), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n911), .ZN(new_n914));
  INV_X1    g728(.A(new_n912), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n898), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n910), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n890), .B(new_n896), .C1(new_n909), .C2(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n895), .A2(new_n911), .A3(new_n912), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n898), .B2(new_n915), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT116), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT116), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n913), .A2(new_n922), .A3(new_n916), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n921), .A2(new_n900), .A3(new_n923), .A4(new_n908), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT118), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n910), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n924), .B2(new_n910), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n883), .A2(new_n886), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n835), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT119), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n933), .B(new_n835), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(G75));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n464), .B1(new_n871), .B2(new_n882), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT56), .B1(new_n937), .B2(G210), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n399), .A2(new_n401), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n402), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT55), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n936), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n257), .A2(G952), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n938), .B2(new_n942), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n938), .A2(new_n936), .A3(new_n942), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(G51));
  XOR2_X1   g762(.A(new_n752), .B(KEYINPUT57), .Z(new_n949));
  AOI21_X1  g763(.A(new_n872), .B1(new_n871), .B2(new_n882), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n883), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n466), .A2(new_n467), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n937), .A2(new_n805), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(G54));
  NAND3_X1  g769(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .ZN(new_n956));
  INV_X1    g770(.A(new_n246), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n944), .ZN(G60));
  OR2_X1    g774(.A1(new_n883), .A2(new_n886), .ZN(new_n961));
  XOR2_X1   g775(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n264), .A2(new_n464), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n778), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n778), .B(new_n964), .C1(new_n883), .C2(new_n950), .ZN(new_n966));
  INV_X1    g780(.A(new_n944), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n965), .A2(new_n968), .ZN(G63));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT61), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT124), .Z(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n871), .A2(new_n882), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT122), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n656), .A2(new_n658), .ZN(new_n979));
  OAI221_X1 g793(.A(new_n967), .B1(new_n970), .B2(KEYINPUT61), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n512), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n973), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n978), .A2(new_n979), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n967), .B1(new_n970), .B2(KEYINPUT61), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n972), .A3(new_n981), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n987), .ZN(G66));
  INV_X1    g802(.A(new_n262), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n257), .B1(new_n989), .B2(G224), .ZN(new_n990));
  INV_X1    g804(.A(new_n875), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n991), .A2(new_n848), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n992), .B2(new_n257), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n939), .B1(G898), .B2(new_n257), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(G69));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n549), .A2(new_n550), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(new_n241), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n824), .A2(new_n520), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n646), .B1(new_n255), .B2(new_n632), .ZN(new_n1001));
  OR3_X1    g815(.A1(new_n680), .A2(new_n1001), .A3(new_n756), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI22_X1  g817(.A1(new_n1000), .A2(new_n1003), .B1(new_n800), .B2(new_n810), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n826), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n879), .A2(new_n706), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n702), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n879), .A2(new_n706), .ZN(new_n1009));
  INV_X1    g823(.A(new_n702), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT62), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1005), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n999), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  NAND2_X1  g828(.A1(G900), .A2(G953), .ZN(new_n1015));
  INV_X1    g829(.A(new_n775), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n799), .B1(new_n725), .B2(new_n769), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1016), .B1(new_n810), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n826), .A2(new_n1018), .A3(new_n852), .A4(new_n1009), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n998), .B(new_n1015), .C1(new_n1019), .C2(G953), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n257), .B1(G227), .B2(G900), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT125), .Z(new_n1022));
  NAND4_X1  g836(.A1(new_n1013), .A2(new_n1014), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1011), .A2(new_n1008), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n811), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n825), .B2(new_n817), .ZN(new_n1027));
  AOI21_X1  g841(.A(G953), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1020), .B(new_n1022), .C1(new_n1028), .C2(new_n998), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(KEYINPUT126), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1021), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n996), .B(new_n1023), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1008), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n1007), .A2(new_n702), .A3(new_n1006), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1027), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n998), .B1(new_n1037), .B2(new_n257), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n998), .A2(new_n1015), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1019), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1039), .B1(new_n1040), .B2(new_n257), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1021), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1042), .A2(KEYINPUT126), .A3(new_n1029), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n996), .B1(new_n1043), .B2(new_n1023), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1034), .A2(new_n1044), .ZN(G72));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  OAI21_X1  g861(.A(new_n1047), .B1(new_n992), .B2(new_n1019), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n682), .A2(new_n528), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n944), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OR2_X1    g864(.A1(new_n992), .A2(new_n1037), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n1051), .A2(new_n1047), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1050), .B1(new_n1052), .B2(new_n683), .ZN(new_n1053));
  INV_X1    g867(.A(new_n1049), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1054), .A2(new_n683), .A3(new_n1047), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1055), .B1(new_n871), .B2(new_n885), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n1053), .A2(new_n1056), .ZN(G57));
endmodule


