//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n465), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT66), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(new_n480), .A3(new_n472), .ZN(new_n484));
  OAI221_X1 g059(.A(new_n476), .B1(new_n481), .B2(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n472), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n479), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n462), .A2(new_n464), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n472), .B2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT67), .B1(new_n501), .B2(KEYINPUT68), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT5), .B1(new_n501), .B2(KEYINPUT67), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(KEYINPUT67), .B(KEYINPUT5), .C1(new_n501), .C2(KEYINPUT68), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n504), .A2(new_n505), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n510), .A2(G88), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n509), .A2(new_n514), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n504), .A2(G63), .A3(new_n505), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G51), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n515), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT70), .B(G89), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n504), .A2(new_n505), .A3(new_n513), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n522), .A2(new_n529), .ZN(G168));
  NAND3_X1  g105(.A1(new_n504), .A2(G64), .A3(new_n505), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n519), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n504), .A2(G90), .A3(new_n505), .A4(new_n513), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  NAND3_X1  g112(.A1(new_n504), .A2(G56), .A3(new_n505), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n519), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n504), .A2(G81), .A3(new_n505), .A4(new_n513), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n515), .A2(G43), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT71), .Z(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n515), .A2(G53), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(KEYINPUT72), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n552), .B(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G91), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT73), .B(G65), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n504), .A2(new_n505), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n558), .B1(new_n562), .B2(G651), .ZN(new_n563));
  AOI211_X1 g138(.A(KEYINPUT74), .B(new_n519), .C1(new_n560), .C2(new_n561), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n555), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(G299));
  INV_X1    g140(.A(new_n533), .ZN(new_n566));
  INV_X1    g141(.A(new_n536), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT75), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(new_n533), .B2(new_n536), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n519), .B1(new_n506), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(G49), .B2(new_n515), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n510), .A2(new_n513), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT76), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n556), .A2(new_n579), .A3(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n504), .A2(G61), .A3(new_n505), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT77), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n519), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n504), .A2(G86), .A3(new_n505), .A4(new_n513), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n515), .A2(G48), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n556), .A2(G85), .B1(G47), .B2(new_n515), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n519), .B2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  INV_X1    g169(.A(G79), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n506), .A2(new_n594), .B1(new_n595), .B2(new_n501), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  OAI221_X1 g173(.A(new_n598), .B1(new_n595), .B2(new_n501), .C1(new_n506), .C2(new_n594), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(G651), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n504), .A2(G92), .A3(new_n505), .A4(new_n513), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT10), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n515), .A2(G54), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT78), .B1(new_n605), .B2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  MUX2_X1   g182(.A(KEYINPUT78), .B(new_n606), .S(new_n607), .Z(G284));
  MUX2_X1   g183(.A(KEYINPUT78), .B(new_n606), .S(new_n607), .Z(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  XNOR2_X1  g187(.A(G280), .B(KEYINPUT80), .ZN(G297));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n605), .B1(new_n614), .B2(G860), .ZN(G148));
  OAI21_X1  g190(.A(KEYINPUT81), .B1(new_n544), .B2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n605), .A2(new_n614), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  MUX2_X1   g193(.A(KEYINPUT81), .B(new_n616), .S(new_n618), .Z(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g195(.A(G135), .ZN(new_n621));
  OR3_X1    g196(.A1(new_n484), .A2(KEYINPUT82), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n481), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G123), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT82), .B1(new_n484), .B2(new_n621), .ZN(new_n627));
  NAND4_X1  g202(.A1(new_n622), .A2(new_n624), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2438), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2451), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n646), .B(new_n647), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(KEYINPUT85), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(KEYINPUT85), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n654), .B(KEYINPUT17), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n657), .C1(new_n653), .C2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT86), .ZN(new_n661));
  INV_X1    g236(.A(new_n651), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n653), .A2(new_n654), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n651), .A3(new_n653), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n629), .ZN(new_n667));
  INV_X1    g242(.A(G2100), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n672), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n682), .C1(new_n680), .C2(new_n679), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT88), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n684), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  NOR2_X1   g267(.A1(G16), .A2(G21), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G168), .B2(G16), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G1966), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n696), .A2(G28), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(G28), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G5), .A2(G16), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G171), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G1961), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(G27), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G164), .B2(new_n699), .ZN(new_n707));
  AOI211_X1 g282(.A(new_n695), .B(new_n705), .C1(G2078), .C2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT24), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n699), .B1(new_n709), .B2(G34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT98), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(G34), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT98), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(new_n699), .C1(new_n709), .C2(G34), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n468), .A2(new_n473), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n699), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT100), .Z(new_n721));
  INV_X1    g296(.A(G2084), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n707), .A2(G2078), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n628), .A2(new_n699), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  NOR4_X1   g301(.A1(new_n723), .A2(new_n724), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2090), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n485), .A2(G29), .ZN(new_n729));
  INV_X1    g304(.A(G35), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(G29), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n729), .B(new_n733), .C1(G29), .C2(new_n730), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n484), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G139), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  NAND2_X1  g314(.A1(G115), .A2(G2104), .ZN(new_n740));
  INV_X1    g315(.A(G127), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n465), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT96), .B1(new_n742), .B2(G2105), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(G2105), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n737), .B(new_n739), .C1(new_n743), .C2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT97), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n744), .B(new_n745), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n750), .A2(KEYINPUT97), .A3(new_n737), .A4(new_n739), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n751), .A3(G29), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G29), .B2(G33), .ZN(new_n754));
  OR3_X1    g329(.A1(new_n753), .A2(G29), .A3(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G2072), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n752), .A2(new_n758), .A3(new_n754), .A4(new_n755), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n735), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n702), .A2(G1961), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AND4_X1   g337(.A1(new_n708), .A2(new_n727), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G32), .ZN(new_n764));
  AOI22_X1  g339(.A1(G129), .A2(new_n623), .B1(new_n736), .B2(G141), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT101), .Z(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT102), .B(KEYINPUT26), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n765), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n764), .B1(new_n772), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT27), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1996), .ZN(new_n775));
  NOR2_X1   g350(.A1(G104), .A2(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n778));
  INV_X1    g353(.A(G128), .ZN(new_n779));
  INV_X1    g354(.A(G140), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n778), .B1(new_n481), .B2(new_n779), .C1(new_n780), .C2(new_n484), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n699), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT28), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n782), .A2(G2067), .A3(new_n785), .ZN(new_n789));
  INV_X1    g364(.A(G16), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G19), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n544), .B2(new_n790), .ZN(new_n792));
  INV_X1    g367(.A(G1341), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n788), .A2(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n790), .A2(G4), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n604), .B2(G16), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(G1348), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(G1348), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT94), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n732), .A2(new_n728), .A3(new_n734), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n763), .A2(new_n775), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n790), .A2(G22), .ZN(new_n805));
  AOI211_X1 g380(.A(KEYINPUT91), .B(new_n805), .C1(G303), .C2(G16), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n508), .A2(G651), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n514), .A2(new_n516), .ZN(new_n809));
  OAI21_X1  g384(.A(G16), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n805), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n807), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G1971), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n806), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT91), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n810), .A2(new_n807), .A3(new_n811), .ZN(new_n817));
  AOI21_X1  g392(.A(G1971), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G1976), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n575), .A2(new_n578), .A3(new_n580), .A4(G16), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n822));
  OR2_X1    g397(.A1(G16), .A2(G23), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n821), .A2(new_n823), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT33), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n829), .A2(G1976), .A3(new_n824), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n790), .A2(G6), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n589), .B2(new_n790), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT32), .B(G1981), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT90), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n819), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n819), .A2(new_n831), .A3(KEYINPUT34), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G1986), .ZN(new_n842));
  NAND2_X1  g417(.A1(G290), .A2(G16), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT89), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n790), .A2(G24), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n842), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n848), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n850), .A2(G1986), .A3(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n699), .A2(G25), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n623), .A2(G119), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n736), .A2(G131), .ZN(new_n854));
  OR2_X1    g429(.A1(G95), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n852), .B1(new_n858), .B2(new_n699), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G1991), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n849), .A2(new_n851), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n841), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT36), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n841), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n804), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n721), .A2(new_n722), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n790), .A2(KEYINPUT23), .A3(G20), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT23), .ZN(new_n872));
  INV_X1    g447(.A(G20), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(G16), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n874), .C1(new_n611), .C2(new_n790), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(G1956), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n694), .A2(G1966), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n869), .A2(new_n870), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(G311));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI211_X1 g456(.A(new_n761), .B(new_n735), .C1(new_n757), .C2(new_n759), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n882), .A2(new_n803), .A3(new_n708), .A4(new_n727), .ZN(new_n883));
  INV_X1    g458(.A(G1996), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n774), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT94), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n801), .B(new_n886), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n867), .B1(new_n841), .B2(new_n864), .ZN(new_n889));
  AOI211_X1 g464(.A(KEYINPUT36), .B(new_n863), .C1(new_n839), .C2(new_n840), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n888), .B(new_n877), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(KEYINPUT103), .A3(new_n870), .A4(new_n876), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n881), .A2(new_n893), .ZN(G150));
  NAND2_X1  g469(.A1(G80), .A2(G543), .ZN(new_n895));
  INV_X1    g470(.A(G67), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n506), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G651), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n504), .A2(G93), .A3(new_n505), .A4(new_n513), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n515), .A2(G55), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G860), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT37), .Z(new_n904));
  NOR2_X1   g479(.A1(new_n604), .A2(new_n614), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT39), .ZN(new_n906));
  XNOR2_X1  g481(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n544), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n898), .B(new_n901), .C1(new_n540), .C2(new_n543), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n908), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n904), .B1(new_n912), .B2(G860), .ZN(G145));
  NAND3_X1  g488(.A1(new_n462), .A2(new_n464), .A3(new_n492), .ZN(new_n914));
  INV_X1    g489(.A(G102), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n472), .ZN(new_n916));
  INV_X1    g491(.A(G114), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G2105), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n918), .A3(G2104), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n914), .B2(new_n919), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n489), .B(new_n490), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n781), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(new_n772), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n749), .A2(new_n751), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n926), .A2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n924), .B(new_n771), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G142), .ZN(new_n935));
  NOR2_X1   g510(.A1(G106), .A2(G2105), .ZN(new_n936));
  OAI21_X1  g511(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n484), .A2(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(G130), .B2(new_n623), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(new_n632), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(new_n858), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n931), .A2(new_n943), .A3(new_n933), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n485), .B(KEYINPUT105), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(new_n719), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(new_n628), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n942), .A2(new_n948), .A3(new_n944), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g529(.A1(G305), .A2(KEYINPUT109), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n589), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(G303), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(G288), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n959), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT42), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n604), .B(G299), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n611), .A2(new_n604), .ZN(new_n971));
  NAND4_X1  g546(.A1(G299), .A2(new_n600), .A3(new_n603), .A4(new_n602), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(KEYINPUT108), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT41), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n611), .A2(new_n975), .A3(new_n604), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(KEYINPUT41), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n617), .B(new_n911), .ZN(new_n981));
  MUX2_X1   g556(.A(new_n970), .B(new_n980), .S(new_n981), .Z(new_n982));
  XNOR2_X1  g557(.A(new_n969), .B(new_n982), .ZN(new_n983));
  MUX2_X1   g558(.A(new_n902), .B(new_n983), .S(G868), .Z(G295));
  MUX2_X1   g559(.A(new_n902), .B(new_n983), .S(G868), .Z(G331));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n909), .A2(new_n910), .ZN(new_n987));
  NAND2_X1  g562(.A1(G301), .A2(G168), .ZN(new_n988));
  NOR3_X1   g563(.A1(G168), .A2(new_n533), .A3(new_n536), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G286), .B1(new_n568), .B2(new_n570), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n911), .B1(new_n992), .B2(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n979), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n991), .B2(new_n993), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n992), .A2(new_n989), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT112), .B1(new_n1000), .B2(new_n987), .ZN(new_n1001));
  OR3_X1    g576(.A1(new_n999), .A2(new_n970), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n979), .A2(new_n994), .A3(KEYINPUT111), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n997), .A2(new_n968), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n960), .B(new_n961), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n966), .B1(new_n1005), .B2(new_n959), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n973), .A2(KEYINPUT41), .A3(new_n976), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n999), .B2(new_n1001), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n970), .B1(new_n1008), .B2(new_n994), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1007), .B(KEYINPUT41), .C1(new_n999), .C2(new_n1001), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1004), .A2(new_n1012), .A3(new_n951), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1004), .A2(new_n1012), .A3(new_n1015), .A4(new_n951), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n986), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n997), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1006), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(new_n951), .A3(new_n1004), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1020), .A2(new_n986), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT44), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1013), .A2(KEYINPUT43), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1022), .A2(new_n1027), .ZN(G397));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n1029));
  AND2_X1   g604(.A1(G160), .A2(G40), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n489), .A2(new_n490), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT106), .B1(new_n493), .B2(new_n496), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT117), .B1(new_n1034), .B2(G1384), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n923), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1029), .B(new_n1030), .C1(new_n1039), .C2(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1041));
  AOI211_X1 g616(.A(KEYINPUT117), .B(G1384), .C1(new_n1041), .C2(new_n491), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1036), .B1(new_n923), .B2(new_n1037), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1030), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(KEYINPUT122), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n491), .B2(new_n497), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT45), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1040), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1966), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G160), .A2(G40), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n498), .A2(new_n1037), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1054), .B1(KEYINPUT50), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1057), .A2(G2084), .ZN(new_n1058));
  OAI21_X1  g633(.A(G286), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1058), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1060), .B1(new_n1061), .B2(G168), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1062), .A3(KEYINPUT51), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  AOI211_X1 g639(.A(G286), .B(new_n1058), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n1060), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT45), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1055), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n923), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1030), .A3(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT116), .B(G1971), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1057), .B2(G2090), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G303), .A2(G8), .ZN(new_n1078));
  XOR2_X1   g653(.A(new_n1078), .B(KEYINPUT55), .Z(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(G8), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1054), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n1060), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n582), .A2(new_n584), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G651), .ZN(new_n1085));
  INV_X1    g660(.A(new_n588), .ZN(new_n1086));
  INV_X1    g661(.A(G1981), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(G1981), .B1(new_n585), .B2(new_n588), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1083), .B1(new_n1090), .B2(KEYINPUT118), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1092), .B(KEYINPUT49), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1044), .B(G8), .C1(new_n820), .C2(G288), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1082), .A2(new_n1094), .B1(new_n1095), .B2(KEYINPUT52), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(G288), .B2(new_n820), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1082), .B(new_n1097), .C1(new_n820), .C2(G288), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1080), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT121), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1102), .B(new_n1030), .C1(new_n1039), .C2(new_n1052), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1030), .A2(new_n1052), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1044), .A2(KEYINPUT120), .A3(new_n1104), .ZN(new_n1105));
  AOI211_X1 g680(.A(G2090), .B(new_n1101), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1076), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1079), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1099), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G2078), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1040), .A2(new_n1046), .A3(new_n1048), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G2078), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1071), .A2(new_n1114), .A3(new_n1030), .A4(new_n1072), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1057), .A2(new_n704), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(G301), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1063), .A2(KEYINPUT62), .A3(new_n1066), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1069), .A2(new_n1110), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G299), .A2(KEYINPUT123), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT57), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1073), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT56), .B(G2072), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1101), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1121), .B(new_n1124), .C1(new_n1125), .C2(G1956), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1081), .A2(new_n787), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1057), .ZN(new_n1131));
  OAI221_X1 g706(.A(new_n1130), .B1(KEYINPUT60), .B2(new_n605), .C1(new_n1131), .C2(G1348), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT58), .B(G1341), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1073), .A2(G1996), .B1(new_n1081), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT124), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  OAI221_X1 g713(.A(new_n1138), .B1(new_n1081), .B2(new_n1135), .C1(G1996), .C2(new_n1073), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1139), .A3(new_n544), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1137), .A2(new_n1139), .A3(new_n1142), .A4(new_n544), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1129), .A2(new_n1134), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1130), .B1(new_n1131), .B2(G1348), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1126), .A2(new_n605), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1124), .B1(new_n1125), .B2(G1956), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1121), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1112), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1030), .A2(new_n1072), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT45), .B1(new_n923), .B2(new_n1037), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1116), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1158), .B2(G171), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1113), .A2(G301), .A3(new_n1116), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1113), .A2(KEYINPUT126), .A3(new_n1116), .A4(G301), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1063), .A2(new_n1066), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1146), .A2(new_n605), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1150), .A2(KEYINPUT61), .A3(new_n1126), .A4(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G301), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1158), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1153), .B1(new_n1169), .B2(new_n1117), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1110), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1152), .A2(new_n1165), .A3(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1061), .A2(new_n1060), .A3(G286), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1077), .A2(G8), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1176), .B1(new_n1177), .B2(new_n1109), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1173), .A2(new_n1080), .A3(new_n1175), .A4(new_n1178), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1110), .A2(new_n1173), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(KEYINPUT63), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1174), .A2(new_n1080), .ZN(new_n1182));
  NOR2_X1   g757(.A1(G288), .A2(G1976), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT119), .Z(new_n1184));
  OAI21_X1  g759(.A(new_n1088), .B1(new_n1184), .B2(new_n1094), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1182), .B1(new_n1082), .B2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1119), .A2(new_n1172), .A3(new_n1181), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1030), .A2(new_n1156), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n781), .B(G2067), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT115), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n771), .A2(G1996), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n772), .A2(new_n1188), .A3(new_n884), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1194), .A2(KEYINPUT114), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(KEYINPUT114), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OR2_X1    g772(.A1(new_n857), .A2(new_n860), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n857), .A2(new_n860), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1188), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(G290), .B(G1986), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1201), .B1(new_n1189), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1187), .A2(new_n1203), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n781), .A2(G2067), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1188), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1191), .A2(new_n771), .ZN(new_n1208));
  OAI21_X1  g783(.A(KEYINPUT46), .B1(new_n1188), .B2(G1996), .ZN(new_n1209));
  OR3_X1    g784(.A1(new_n1188), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1208), .A2(new_n1189), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT47), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1188), .A2(G290), .A3(G1986), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT127), .ZN(new_n1214));
  XNOR2_X1  g789(.A(new_n1214), .B(KEYINPUT48), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1201), .A2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1207), .A2(new_n1212), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1204), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g793(.A1(G319), .A2(new_n953), .A3(new_n649), .A4(new_n669), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n1220), .A2(new_n1025), .A3(new_n691), .ZN(G225));
  INV_X1    g795(.A(G225), .ZN(G308));
endmodule


