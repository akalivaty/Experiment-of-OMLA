//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT75), .A2(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(new_n188), .ZN(new_n194));
  NAND3_X1  g008(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n192), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n199));
  AOI21_X1  g013(.A(G140), .B1(KEYINPUT75), .B2(G125), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n197), .B(KEYINPUT16), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n187), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT16), .B1(new_n199), .B2(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT76), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n205), .A2(G146), .A3(new_n201), .A4(new_n192), .ZN(new_n206));
  NOR2_X1   g020(.A1(G237), .A2(G953), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G214), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(G143), .A3(G214), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT17), .A3(G131), .ZN(new_n213));
  INV_X1    g027(.A(new_n211), .ZN(new_n214));
  AOI21_X1  g028(.A(G143), .B1(new_n207), .B2(G214), .ZN(new_n215));
  OAI21_X1  g029(.A(G131), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(new_n217), .A3(new_n211), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n203), .A2(new_n206), .A3(new_n213), .A4(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n212), .A2(KEYINPUT18), .A3(G131), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT65), .B(G146), .ZN(new_n223));
  INV_X1    g037(.A(G125), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G140), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n189), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n194), .A2(G146), .A3(new_n195), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT18), .A2(G131), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n210), .A2(new_n211), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n222), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G113), .B(G122), .ZN(new_n232));
  INV_X1    g046(.A(G104), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n232), .B(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n221), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n206), .A2(KEYINPUT78), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n204), .A2(KEYINPUT76), .B1(new_n191), .B2(new_n190), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT78), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G146), .A4(new_n201), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n216), .A2(new_n218), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT19), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n189), .A2(new_n225), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT87), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n194), .A2(KEYINPUT19), .A3(new_n195), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n243), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n244), .A2(new_n223), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n236), .A2(new_n239), .A3(new_n240), .A4(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n248), .A2(new_n231), .ZN(new_n249));
  OAI211_X1 g063(.A(KEYINPUT88), .B(new_n235), .C1(new_n249), .C2(new_n234), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT88), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n234), .B1(new_n248), .B2(new_n231), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n221), .A2(new_n231), .A3(new_n234), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G475), .A2(G902), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT20), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n259), .A3(KEYINPUT20), .ZN(new_n260));
  NOR3_X1   g074(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n252), .B2(new_n253), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n234), .B1(new_n221), .B2(new_n231), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n253), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G475), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(G478), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT13), .B1(new_n272), .B2(G143), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G128), .B(G143), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G122), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G116), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G122), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G107), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n282), .B1(new_n279), .B2(new_n281), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n286), .ZN(new_n288));
  AOI21_X1  g102(.A(G107), .B1(new_n288), .B2(new_n283), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n277), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n276), .B(new_n274), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n293), .A2(new_n279), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n291), .B(new_n292), .C1(new_n295), .C2(new_n285), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(G953), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT91), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT91), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n290), .A2(new_n302), .A3(new_n296), .A4(new_n299), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n290), .A2(new_n296), .ZN(new_n304));
  INV_X1    g118(.A(new_n299), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT93), .A3(new_n264), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT93), .B1(new_n307), .B2(new_n264), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n271), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n270), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(G234), .A2(G237), .ZN(new_n314));
  INV_X1    g128(.A(G953), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n314), .A2(G952), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n314), .A2(G902), .A3(G953), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT21), .B(G898), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n268), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n187), .A2(KEYINPUT65), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n323), .A3(G143), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n187), .A2(G143), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n272), .B1(new_n324), .B2(KEYINPUT1), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n187), .A2(G143), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n321), .A2(new_n323), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(new_n209), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n328), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n274), .A2(G137), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n274), .A2(G137), .ZN(new_n337));
  OAI21_X1  g151(.A(G131), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n274), .B2(G137), .ZN(new_n340));
  INV_X1    g154(.A(G137), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT11), .A3(G134), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n340), .A2(new_n342), .A3(new_n217), .A4(new_n335), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n334), .A2(KEYINPUT67), .A3(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n340), .A2(new_n335), .A3(new_n342), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G131), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n343), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n330), .B1(new_n223), .B2(G143), .ZN(new_n352));
  XOR2_X1   g166(.A(KEYINPUT0), .B(G128), .Z(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n324), .A2(KEYINPUT0), .A3(G128), .A4(new_n326), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n351), .A2(new_n354), .A3(KEYINPUT66), .A4(new_n355), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n347), .A2(new_n348), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(G116), .B(G119), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT2), .B(G113), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(KEYINPUT68), .B2(new_n363), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n345), .A2(KEYINPUT30), .A3(new_n356), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n362), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n369), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n345), .A2(new_n356), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT26), .B(G101), .Z(new_n375));
  NAND2_X1  g189(.A1(new_n207), .A2(G210), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n373), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT70), .B1(new_n382), .B2(KEYINPUT28), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT70), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n373), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n382), .B1(new_n360), .B2(new_n369), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n387), .B(new_n379), .C1(new_n385), .C2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n372), .B1(new_n345), .B2(new_n356), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT28), .B1(new_n382), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n379), .A2(KEYINPUT29), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n383), .A2(new_n392), .A3(new_n386), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n264), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT71), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(KEYINPUT71), .A3(new_n264), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G472), .B1(new_n390), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n371), .A2(new_n379), .A3(new_n373), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT31), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n388), .A2(new_n385), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n383), .A2(new_n386), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n380), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT31), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n371), .A2(new_n406), .A3(new_n379), .A4(new_n373), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n409));
  NOR2_X1   g223(.A1(G472), .A2(G902), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n408), .B2(new_n410), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n400), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G140), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n315), .A2(G227), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n325), .B1(new_n223), .B2(G143), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n272), .B1(new_n330), .B2(KEYINPUT1), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n328), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT3), .B1(new_n233), .B2(G107), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n285), .A3(G104), .ZN(new_n425));
  INV_X1    g239(.A(G101), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n233), .A2(G107), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n423), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n233), .A2(G107), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n285), .A2(G104), .ZN(new_n430));
  OAI21_X1  g244(.A(G101), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n422), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G101), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n438), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n428), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(G101), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n439), .A2(new_n355), .A3(new_n354), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT81), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n428), .A2(new_n431), .A3(KEYINPUT10), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n334), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n334), .B2(new_n444), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n436), .B(new_n442), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n419), .B1(new_n447), .B2(new_n351), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n436), .A2(new_n442), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n334), .A2(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n334), .A2(new_n443), .A3(new_n444), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n350), .A2(new_n343), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n453), .A3(KEYINPUT82), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n447), .A2(new_n351), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n418), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n432), .B(new_n328), .C1(new_n329), .C2(new_n333), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n434), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT12), .B1(new_n460), .B2(new_n351), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT12), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n462), .B(new_n454), .C1(new_n434), .C2(new_n459), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n417), .B(new_n464), .C1(new_n448), .C2(new_n455), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n414), .B(new_n264), .C1(new_n458), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(G469), .A2(G902), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n456), .A2(new_n457), .A3(new_n418), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n448), .B2(new_n455), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(G469), .C1(new_n418), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT79), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G214), .B1(G237), .B2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n354), .A2(new_n355), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G125), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n224), .B(new_n328), .C1(new_n329), .C2(new_n333), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n315), .A2(G224), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n482), .B(new_n483), .Z(new_n484));
  NAND3_X1  g298(.A1(new_n439), .A2(new_n369), .A3(new_n441), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n363), .A2(KEYINPUT5), .ZN(new_n486));
  INV_X1    g300(.A(G119), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G116), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n486), .B(G113), .C1(KEYINPUT5), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n367), .A2(new_n363), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n433), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G122), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT83), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n494), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n485), .A2(new_n493), .A3(new_n491), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n495), .A3(KEYINPUT6), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n484), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n480), .A2(new_n481), .B1(KEYINPUT7), .B2(new_n483), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT84), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT85), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT7), .B1(new_n483), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n506), .B2(new_n483), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n480), .A2(new_n481), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n489), .A2(new_n490), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n432), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n491), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n493), .B(KEYINPUT8), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n480), .A2(KEYINPUT86), .A3(new_n481), .A4(new_n508), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n511), .A2(new_n516), .A3(new_n499), .A4(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n264), .B1(new_n505), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n478), .B1(new_n502), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n505), .A2(new_n518), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n521), .A2(new_n264), .A3(new_n477), .A4(new_n501), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n476), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n471), .A2(new_n474), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n487), .A2(G128), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT72), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n487), .B2(G128), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n526), .A2(new_n528), .B1(new_n487), .B2(G128), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT73), .B1(new_n487), .B2(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT23), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT73), .B(new_n534), .C1(new_n487), .C2(G128), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n535), .A3(new_n525), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n531), .B1(G110), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n236), .A2(new_n537), .A3(new_n239), .A4(new_n226), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n529), .A2(new_n530), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G110), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n536), .B2(new_n540), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n539), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n203), .A2(new_n206), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT77), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT77), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n538), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT22), .B(G137), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n315), .A2(G221), .A3(G234), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n538), .B(new_n551), .C1(new_n546), .C2(new_n547), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n264), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n553), .A2(KEYINPUT25), .A3(new_n264), .A4(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n298), .B1(G234), .B2(new_n264), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(G902), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n554), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n320), .A2(new_n413), .A3(new_n524), .A4(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  AND4_X1   g381(.A1(new_n561), .A2(new_n471), .A3(new_n563), .A4(new_n474), .ZN(new_n568));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n408), .B2(new_n264), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n410), .B2(new_n408), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n319), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n306), .A2(KEYINPUT33), .A3(new_n300), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(KEYINPUT94), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n307), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(KEYINPUT94), .ZN(new_n578));
  INV_X1    g392(.A(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G902), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n575), .A2(new_n577), .A3(new_n578), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n307), .A2(new_n264), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n579), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n268), .A2(new_n523), .A3(new_n573), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n572), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT34), .B(G104), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  INV_X1    g403(.A(new_n523), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n250), .A2(new_n254), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n261), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n258), .A2(new_n260), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n267), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n311), .B2(new_n312), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n573), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n590), .B1(new_n596), .B2(KEYINPUT95), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n595), .A3(new_n598), .A4(new_n573), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n597), .A2(KEYINPUT96), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT96), .B1(new_n597), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n572), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G107), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  OR2_X1    g418(.A1(new_n552), .A2(KEYINPUT36), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n548), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n548), .A2(new_n605), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n606), .A2(new_n562), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n559), .B2(new_n560), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n320), .A2(new_n524), .A3(new_n571), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  INV_X1    g427(.A(G900), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n316), .B1(new_n317), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n593), .A2(new_n595), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n593), .A2(new_n595), .A3(new_n619), .A4(new_n616), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n523), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n618), .A2(KEYINPUT98), .A3(new_n523), .A4(new_n620), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n471), .A2(new_n474), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n413), .A2(new_n625), .A3(new_n610), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT99), .B(G128), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G30));
  XOR2_X1   g443(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n615), .B(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT40), .Z(new_n633));
  OR2_X1    g447(.A1(new_n411), .A2(new_n412), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n380), .B1(new_n371), .B2(new_n373), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n382), .A2(new_n391), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n264), .B1(new_n636), .B2(new_n379), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n609), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n520), .A2(new_n522), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT38), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n642), .A2(new_n475), .A3(new_n268), .A4(new_n313), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n633), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n209), .ZN(G45));
  INV_X1    g459(.A(new_n584), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n615), .B(new_n646), .C1(new_n263), .C2(new_n267), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n413), .A2(new_n647), .A3(new_n524), .A4(new_n610), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G146), .ZN(G48));
  OAI21_X1  g463(.A(new_n264), .B1(new_n458), .B2(new_n465), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(KEYINPUT101), .A3(G469), .ZN(new_n651));
  NAND2_X1  g465(.A1(KEYINPUT101), .A2(G469), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n264), .B(new_n652), .C1(new_n458), .C2(new_n465), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n651), .A2(new_n472), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n586), .A2(new_n413), .A3(new_n565), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT41), .B(G113), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G15));
  NAND2_X1  g471(.A1(new_n413), .A2(new_n565), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n659), .B(new_n654), .C1(new_n600), .C2(new_n601), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G116), .ZN(G18));
  AND4_X1   g475(.A1(new_n472), .A2(new_n651), .A3(new_n523), .A4(new_n653), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n320), .A2(new_n413), .A3(new_n662), .A4(new_n610), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  AOI21_X1  g478(.A(new_n404), .B1(KEYINPUT28), .B2(new_n636), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n402), .B(new_n407), .C1(new_n665), .C2(new_n379), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(new_n410), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n667), .A2(new_n564), .A3(new_n570), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n268), .A2(new_n523), .A3(new_n313), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n573), .A4(new_n654), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G122), .ZN(G24));
  NOR3_X1   g485(.A1(new_n667), .A2(new_n570), .A3(new_n609), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n647), .A3(new_n662), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G125), .ZN(G27));
  AND2_X1   g488(.A1(new_n471), .A2(new_n472), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n641), .A2(new_n476), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n413), .A2(new_n565), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(KEYINPUT42), .A3(new_n647), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n680));
  INV_X1    g494(.A(new_n647), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n680), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G131), .ZN(G33));
  NAND2_X1  g498(.A1(new_n618), .A2(new_n620), .ZN(new_n685));
  OR3_X1    g499(.A1(new_n677), .A2(KEYINPUT102), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT102), .B1(new_n677), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G134), .ZN(G36));
  OAI21_X1  g503(.A(new_n468), .B1(new_n418), .B2(new_n469), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n414), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n691), .B2(new_n690), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n467), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n693), .A2(KEYINPUT46), .A3(new_n467), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n466), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n698), .A2(new_n472), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n631), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT103), .Z(new_n701));
  NOR2_X1   g515(.A1(new_n268), .A2(new_n646), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n702), .B2(new_n705), .ZN(new_n707));
  INV_X1    g521(.A(new_n571), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n610), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n676), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n710), .B2(new_n709), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n701), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G137), .ZN(G39));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n699), .B1(KEYINPUT105), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n716), .B1(new_n699), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n676), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n413), .A2(new_n565), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n647), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G140), .ZN(G42));
  AND2_X1   g537(.A1(new_n707), .A2(new_n316), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n654), .A2(new_n676), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n659), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n728), .B(KEYINPUT48), .Z(new_n729));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n730));
  INV_X1    g544(.A(new_n639), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n565), .A3(new_n316), .A4(new_n726), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT113), .Z(new_n733));
  AOI21_X1  g547(.A(new_n646), .B1(new_n263), .B2(new_n267), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n662), .A3(new_n668), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(G952), .A3(new_n315), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n729), .B1(new_n730), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n724), .A2(new_n668), .A3(new_n676), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n651), .A2(new_n653), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n474), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n739), .B1(new_n719), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n268), .A2(new_n584), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n733), .A2(new_n743), .B1(new_n672), .B2(new_n727), .ZN(new_n744));
  NOR2_X1   g558(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n642), .A2(new_n475), .A3(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n724), .A2(new_n654), .A3(new_n668), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n742), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n750), .A2(KEYINPUT114), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  OAI221_X1 g567(.A(new_n738), .B1(new_n730), .B2(new_n737), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n750), .A2(new_n751), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT115), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n648), .A2(new_n673), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n413), .A2(new_n625), .A3(new_n610), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n622), .B2(new_n621), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n762), .B2(new_n624), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n675), .A2(new_n616), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n639), .A3(new_n609), .A4(new_n669), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT108), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n648), .A2(new_n673), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n627), .A2(new_n767), .A3(KEYINPUT108), .A4(new_n765), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n759), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n627), .A2(new_n767), .A3(new_n765), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT52), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n758), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(new_n775), .B2(new_n768), .ZN(new_n776));
  INV_X1    g590(.A(new_n772), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n776), .A2(KEYINPUT109), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n672), .A2(new_n647), .A3(new_n675), .ZN(new_n780));
  INV_X1    g594(.A(new_n413), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n313), .A2(new_n594), .A3(new_n615), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n625), .A2(new_n593), .A3(new_n610), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n676), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n688), .A2(new_n683), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n655), .A2(new_n566), .A3(new_n611), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n268), .A2(new_n584), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT106), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n590), .A2(new_n319), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n734), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n789), .A2(new_n795), .A3(new_n790), .A4(new_n792), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n572), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n268), .B1(new_n311), .B2(new_n312), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n568), .A3(new_n790), .A4(new_n571), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n670), .A2(new_n799), .A3(new_n663), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n787), .A2(new_n797), .A3(new_n800), .A4(new_n660), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n779), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n786), .A2(new_n801), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n775), .A2(KEYINPUT52), .A3(new_n768), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n770), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT110), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT54), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(KEYINPUT53), .B(new_n805), .C1(new_n773), .C2(new_n778), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n807), .A2(new_n814), .A3(new_n808), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n807), .B2(new_n808), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n812), .B(new_n813), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n757), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(G952), .B2(G953), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n740), .B(KEYINPUT49), .Z(new_n820));
  NOR4_X1   g634(.A1(new_n642), .A2(new_n564), .A3(new_n473), .A4(new_n476), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n731), .A2(new_n820), .A3(new_n821), .A4(new_n702), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(G75));
  NOR2_X1   g637(.A1(new_n315), .A2(G952), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n264), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT56), .B1(new_n828), .B2(G210), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n500), .A2(new_n497), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(new_n484), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT55), .Z(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n825), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n829), .B2(new_n833), .ZN(G51));
  NAND2_X1  g649(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(KEYINPUT117), .A3(new_n817), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n826), .A2(new_n838), .A3(KEYINPUT54), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n467), .B(KEYINPUT57), .Z(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n458), .A2(new_n465), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n837), .A2(KEYINPUT118), .A3(new_n839), .A4(new_n840), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n827), .A2(new_n264), .A3(new_n693), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n824), .B1(new_n846), .B2(new_n847), .ZN(G54));
  NAND3_X1  g662(.A1(new_n828), .A2(KEYINPUT58), .A3(G475), .ZN(new_n849));
  INV_X1    g663(.A(new_n591), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n851), .A2(new_n852), .A3(new_n824), .ZN(G60));
  XNOR2_X1  g667(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n579), .A2(new_n264), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n854), .B(new_n855), .Z(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n811), .B2(new_n817), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT119), .Z(new_n859));
  OAI21_X1  g673(.A(new_n825), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n837), .A2(new_n839), .ZN(new_n861));
  INV_X1    g675(.A(new_n856), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(G63));
  AND2_X1   g678(.A1(new_n606), .A2(new_n607), .ZN(new_n865));
  NAND2_X1  g679(.A1(G217), .A2(G902), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT60), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n826), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n869), .A2(new_n825), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n553), .A2(new_n554), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n827), .B2(new_n867), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n873), .B(new_n876), .ZN(G66));
  NAND2_X1  g691(.A1(new_n801), .A2(new_n315), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT122), .ZN(new_n879));
  INV_X1    g693(.A(G224), .ZN(new_n880));
  OAI21_X1  g694(.A(G953), .B1(new_n318), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n830), .B1(G898), .B2(new_n315), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(G69));
  NAND2_X1  g698(.A1(new_n362), .A2(new_n370), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n614), .B2(new_n315), .ZN(new_n888));
  INV_X1    g702(.A(new_n763), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n701), .A2(new_n659), .A3(new_n669), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n713), .A2(new_n722), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n892), .B(new_n893), .C1(new_n891), .C2(new_n890), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n688), .A2(new_n683), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT126), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n888), .B1(new_n897), .B2(new_n315), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n887), .B(KEYINPUT123), .Z(new_n899));
  NOR2_X1   g713(.A1(new_n658), .A2(new_n720), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n789), .A2(new_n792), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n900), .B(new_n632), .C1(new_n901), .C2(new_n798), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n722), .B1(KEYINPUT124), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(KEYINPUT124), .B2(new_n902), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n644), .A2(new_n889), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT62), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(KEYINPUT62), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n904), .A2(new_n713), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n899), .B1(new_n908), .B2(new_n315), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n898), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n315), .B1(G227), .B2(G900), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n910), .B(new_n914), .ZN(G72));
  NAND2_X1  g729(.A1(G472), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT63), .Z(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n908), .B2(new_n801), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n824), .B1(new_n918), .B2(new_n635), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n374), .A2(new_n379), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n894), .A2(new_n801), .A3(new_n896), .ZN(new_n921));
  INV_X1    g735(.A(new_n917), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n804), .A2(new_n810), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n920), .A2(new_n635), .A3(new_n922), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(G57));
endmodule


