//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT69), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n457), .B2(new_n458), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G125), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n472), .B2(new_n462), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G101), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n471), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT71), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n477), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n477), .A2(new_n466), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT72), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n485), .A2(new_n492), .A3(new_n487), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(G162));
  NAND4_X1  g069(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT4), .A4(G138), .ZN(new_n495));
  NAND2_X1  g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n464), .B2(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n500), .B2(new_n466), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n464), .A2(G138), .A3(new_n466), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT73), .A3(G50), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n504), .A2(new_n513), .A3(new_n515), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n511), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT74), .B(G51), .Z(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n505), .B2(new_n524), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT75), .Z(new_n526));
  INV_X1    g101(.A(new_n520), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT7), .Z(new_n530));
  NOR3_X1   g105(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n516), .A2(G64), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n518), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n520), .A2(new_n535), .B1(new_n505), .B2(new_n536), .ZN(new_n537));
  OR3_X1    g112(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT76), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT76), .B1(new_n534), .B2(new_n537), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G171));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n520), .A2(new_n541), .B1(new_n505), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n513), .A2(new_n515), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n551), .A3(G651), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n544), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n546), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n516), .A2(G91), .A3(new_n504), .ZN(new_n565));
  XOR2_X1   g140(.A(KEYINPUT6), .B(G651), .Z(new_n566));
  AND2_X1   g141(.A1(G53), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n568), .B2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n566), .A2(new_n569), .B1(KEYINPUT78), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(KEYINPUT78), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n504), .A2(new_n568), .A3(new_n572), .A4(new_n567), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n564), .A2(new_n565), .A3(new_n571), .A4(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  OR2_X1    g151(.A1(new_n511), .A2(new_n521), .ZN(G303));
  NAND2_X1  g152(.A1(new_n527), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n506), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n520), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n513), .A2(new_n515), .A3(G61), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n518), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT81), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n584), .A2(new_n589), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n527), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n506), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n597), .B(new_n598), .C1(new_n518), .C2(new_n599), .ZN(G290));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n520), .A2(KEYINPUT82), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT82), .B1(new_n520), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n546), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(G54), .A2(new_n506), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n603), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(G171), .ZN(G284));
  OAI21_X1  g190(.A(new_n614), .B1(new_n613), .B2(G171), .ZN(G321));
  NAND2_X1  g191(.A1(G299), .A2(new_n613), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G168), .B2(new_n613), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(G168), .B2(new_n613), .ZN(G280));
  INV_X1    g194(.A(new_n612), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT83), .B(G559), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(G860), .B2(new_n622), .ZN(G148));
  NAND2_X1  g198(.A1(new_n620), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n486), .A2(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n488), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n486), .A2(G135), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT85), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2435), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2438), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2451), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2454), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n649), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n650), .B2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n641), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n640), .A3(new_n654), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n659), .A3(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n666), .B1(new_n671), .B2(new_n665), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT87), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n681), .A2(new_n682), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  OR3_X1    g259(.A1(new_n678), .A2(new_n683), .A3(new_n680), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n684), .B(new_n685), .C1(new_n682), .C2(new_n681), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT88), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1991), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G29), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(G29), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n491), .B2(new_n493), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT29), .B1(new_n701), .B2(new_n696), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(G2090), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G20), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G299), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  INV_X1    g285(.A(G1956), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT100), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n699), .A2(new_n713), .A3(G2090), .A4(new_n702), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n704), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(KEYINPUT102), .ZN(new_n716));
  NOR2_X1   g291(.A1(G5), .A2(G16), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G171), .B2(G16), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT97), .B(G1961), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT28), .ZN(new_n721));
  INV_X1    g296(.A(G26), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n488), .A2(G128), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n486), .A2(G140), .ZN(new_n728));
  OR2_X1    g303(.A1(G104), .A2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n729), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n488), .A2(KEYINPUT94), .A3(G128), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n727), .A2(new_n728), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n723), .B1(new_n733), .B2(new_n721), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2067), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n486), .A2(G139), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n737), .B(new_n738), .C1(new_n466), .C2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  MUX2_X1   g316(.A(G33), .B(new_n741), .S(G29), .Z(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(G2072), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n720), .A2(new_n735), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G168), .A2(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G16), .B2(G21), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G1341), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n554), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G16), .B2(G19), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n746), .A2(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n716), .A2(new_n744), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n715), .A2(KEYINPUT102), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n706), .A2(G4), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n620), .B2(new_n706), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1348), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n488), .A2(G129), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT26), .Z(new_n760));
  AOI22_X1  g335(.A1(new_n464), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n758), .B(new_n760), .C1(G2105), .C2(new_n761), .ZN(new_n762));
  MUX2_X1   g337(.A(G32), .B(new_n762), .S(G29), .Z(new_n763));
  XOR2_X1   g338(.A(KEYINPUT27), .B(G1996), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n636), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  AND2_X1   g343(.A1(KEYINPUT24), .A2(G34), .ZN(new_n769));
  NOR2_X1   g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n700), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n481), .B2(new_n700), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT30), .B(G28), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n772), .A2(new_n773), .B1(new_n700), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n757), .A2(new_n766), .A3(new_n768), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n742), .A2(G2072), .ZN(new_n777));
  NOR2_X1   g352(.A1(G27), .A2(G29), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G164), .B2(G29), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT98), .B(G2078), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n777), .B(new_n781), .C1(new_n749), .C2(new_n751), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n753), .A2(new_n754), .A3(new_n776), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G11), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT36), .ZN(new_n785));
  NOR2_X1   g360(.A1(G6), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n595), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI211_X1 g364(.A(KEYINPUT32), .B(new_n786), .C1(new_n595), .C2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1981), .ZN(new_n791));
  OR3_X1    g366(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n706), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n706), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT33), .B(G1976), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT92), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n795), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n799));
  INV_X1    g374(.A(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G303), .B2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n801), .B1(new_n803), .B2(new_n799), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g381(.A(G1971), .B(new_n801), .C1(new_n803), .C2(new_n799), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n798), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n791), .B1(new_n789), .B2(new_n790), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n792), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n792), .A2(new_n808), .A3(KEYINPUT34), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT90), .Z(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n486), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n488), .A2(G119), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G29), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G25), .B2(G29), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT91), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(KEYINPUT91), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT35), .B(G1991), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n826), .A3(new_n824), .ZN(new_n829));
  MUX2_X1   g404(.A(G24), .B(G290), .S(G16), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G1986), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(G1986), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n828), .A2(new_n829), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n785), .B1(new_n814), .B2(new_n834), .ZN(new_n835));
  AOI211_X1 g410(.A(KEYINPUT36), .B(new_n833), .C1(new_n812), .C2(new_n813), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n783), .B(new_n784), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n772), .A2(new_n773), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT96), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n699), .A2(new_n702), .ZN(new_n840));
  INV_X1    g415(.A(G2090), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT99), .Z(new_n843));
  NOR3_X1   g418(.A1(new_n837), .A2(new_n839), .A3(new_n843), .ZN(G311));
  NOR2_X1   g419(.A1(new_n835), .A2(new_n836), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n753), .A2(new_n776), .A3(new_n782), .ZN(new_n846));
  INV_X1    g421(.A(new_n754), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n839), .ZN(new_n850));
  INV_X1    g425(.A(new_n843), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n784), .ZN(G150));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n520), .A2(new_n853), .B1(new_n505), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n516), .A2(G67), .ZN(new_n857));
  NAND2_X1  g432(.A1(G80), .A2(G543), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G651), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT103), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n518), .B1(new_n857), .B2(new_n858), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n855), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(G860), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n620), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n861), .A2(new_n864), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n553), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n550), .A2(new_n552), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(new_n544), .C1(new_n863), .C2(new_n855), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT39), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n868), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n866), .B1(new_n875), .B2(G860), .ZN(G145));
  NAND2_X1  g451(.A1(new_n488), .A2(G130), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(KEYINPUT104), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT104), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n486), .A2(G142), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(new_n629), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n820), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n469), .A2(new_n471), .A3(G126), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n466), .B1(new_n887), .B2(new_n498), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT4), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n502), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n497), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n762), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n732), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n894), .A2(new_n741), .ZN(new_n895));
  NOR2_X1   g470(.A1(G162), .A2(G160), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n481), .B1(new_n491), .B2(new_n493), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n896), .A2(new_n636), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n636), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n740), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n895), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n895), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n886), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(new_n885), .A3(new_n902), .ZN(new_n907));
  XOR2_X1   g482(.A(KEYINPUT105), .B(G37), .Z(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n869), .A2(G868), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n591), .A2(new_n794), .A3(new_n594), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n794), .B1(new_n591), .B2(new_n594), .ZN(new_n915));
  OAI21_X1  g490(.A(G166), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n595), .A2(G288), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n591), .A2(new_n794), .A3(new_n594), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(G303), .A3(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(G290), .B(KEYINPUT108), .Z(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n916), .B2(new_n919), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n924), .A2(KEYINPUT109), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(KEYINPUT109), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n921), .A2(new_n922), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT109), .A3(new_n924), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n624), .B(new_n873), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n620), .A2(KEYINPUT106), .A3(new_n709), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n612), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(KEYINPUT41), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n612), .A2(new_n934), .A3(new_n935), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n935), .B1(new_n612), .B2(new_n934), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n931), .A2(new_n932), .A3(new_n937), .A4(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n931), .A2(new_n937), .A3(new_n941), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n939), .A2(new_n940), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n931), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n942), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n930), .B(new_n947), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n911), .B(new_n913), .C1(new_n948), .C2(new_n613), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n943), .A2(new_n946), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n930), .A2(new_n950), .A3(new_n942), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n927), .A3(new_n929), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n613), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT110), .B1(new_n953), .B2(new_n912), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n954), .ZN(G295));
  OAI21_X1  g530(.A(new_n913), .B1(new_n948), .B2(new_n613), .ZN(G331));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n871), .A2(new_n544), .B1(new_n861), .B2(new_n864), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n553), .B1(new_n860), .B2(new_n856), .ZN(new_n959));
  OAI21_X1  g534(.A(G301), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n870), .A2(new_n872), .A3(G171), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n960), .A2(G168), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G168), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n944), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n870), .A2(G171), .A3(new_n872), .ZN(new_n965));
  AOI21_X1  g540(.A(G171), .B1(new_n870), .B2(new_n872), .ZN(new_n966));
  OAI21_X1  g541(.A(G286), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(G168), .A3(new_n961), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n941), .A3(new_n937), .A4(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n928), .A2(new_n964), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT111), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n928), .A2(new_n964), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n964), .A2(new_n969), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n923), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n975), .A3(new_n908), .A4(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n971), .B2(new_n973), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n980), .B2(new_n977), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n957), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AND4_X1   g557(.A1(KEYINPUT43), .A2(new_n974), .A3(new_n908), .A4(new_n977), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n980), .B2(new_n977), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(G397));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(G1384), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n892), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G40), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n479), .B2(new_n466), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n472), .A2(new_n462), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT70), .B1(new_n993), .B2(G2105), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n461), .B(new_n466), .C1(new_n472), .C2(new_n462), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n992), .B(KEYINPUT114), .C1(new_n994), .C2(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n990), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n732), .B(G2067), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n762), .B(G1996), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n827), .A3(new_n820), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n732), .A2(G2067), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n1008));
  OR3_X1    g583(.A1(new_n1001), .A2(new_n1008), .A3(G1996), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1001), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n762), .B2(new_n1002), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1001), .B2(G1996), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  OR2_X1    g589(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n820), .B(new_n827), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1001), .A2(G1986), .A3(G290), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT48), .Z(new_n1019));
  AOI211_X1 g594(.A(new_n1007), .B(new_n1014), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT50), .B1(new_n892), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  AOI211_X1 g598(.A(new_n1023), .B(G1384), .C1(new_n890), .C2(new_n891), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1000), .B(new_n773), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(G164), .B2(G1384), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n892), .A2(new_n1021), .A3(new_n989), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1000), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n747), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1023), .B1(G164), .B2(G1384), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n892), .A2(KEYINPUT50), .A3(new_n1021), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1035), .A2(KEYINPUT120), .A3(new_n773), .A4(new_n1000), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1027), .A2(new_n1032), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G286), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(KEYINPUT121), .A3(new_n1039), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G288), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G164), .A2(G1384), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1038), .B(new_n1046), .C1(new_n1000), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT117), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT118), .B1(new_n592), .B2(new_n791), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  NOR4_X1   g627(.A1(new_n584), .A2(new_n589), .A3(new_n1052), .A4(G1981), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1051), .A2(new_n1053), .B1(new_n791), .B2(new_n592), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1038), .B1(new_n1000), .B2(new_n1047), .ZN(new_n1057));
  OAI221_X1 g632(.A(KEYINPUT49), .B1(new_n791), .B2(new_n592), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(G288), .A2(new_n1045), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1046), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1057), .A2(new_n1049), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n999), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT114), .B1(new_n475), .B2(new_n992), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1047), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(G8), .A3(new_n1061), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT52), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1050), .A2(new_n1059), .A3(new_n1062), .A4(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G166), .A2(new_n1038), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n989), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(G164), .B2(G1384), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n892), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1000), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n805), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1022), .A2(new_n1024), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(G2090), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1072), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT122), .B1(new_n1069), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(G8), .A3(new_n1072), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT52), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1067), .B1(new_n1066), .B2(KEYINPUT52), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1072), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1033), .A2(new_n1034), .B1(new_n998), .B2(new_n999), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n805), .A2(new_n1076), .B1(new_n1088), .B2(new_n841), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1087), .B1(new_n1089), .B2(new_n1038), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1062), .A2(new_n1059), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1085), .A2(new_n1086), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1044), .A2(new_n1081), .A3(new_n1082), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT63), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1069), .A2(new_n1082), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1059), .A2(new_n1045), .A3(new_n794), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1095), .B1(new_n1057), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1961), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1078), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1078), .A2(KEYINPUT125), .A3(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n991), .B(new_n473), .C1(new_n466), .C2(new_n479), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n988), .B2(new_n989), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1108), .B1(new_n1110), .B2(KEYINPUT126), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1112), .B(new_n1109), .C1(new_n988), .C2(new_n989), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(new_n1075), .A3(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(G171), .B(KEYINPUT54), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1106), .B1(new_n1076), .B2(G2078), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1105), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1116), .B(new_n1101), .C1(new_n1031), .C2(new_n1108), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1027), .A2(G168), .A3(new_n1032), .A4(new_n1036), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(G8), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1037), .A2(G286), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(G8), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT51), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1121), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1000), .A2(new_n1074), .A3(new_n1075), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n564), .A2(KEYINPUT123), .A3(new_n565), .ZN(new_n1133));
  AOI21_X1  g708(.A(G299), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(G299), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1131), .B(new_n1137), .C1(new_n1088), .C2(G1956), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n612), .ZN(new_n1140));
  INV_X1    g715(.A(G2067), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1000), .A2(new_n1141), .A3(new_n1047), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1088), .B2(G1348), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1078), .A2(new_n711), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1131), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1135), .A2(new_n1146), .A3(new_n1136), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1136), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n1148), .B2(new_n1134), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1140), .A2(new_n1143), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1137), .B1(new_n1144), .B2(new_n1131), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1139), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1142), .B(KEYINPUT60), .C1(new_n1088), .C2(G1348), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n620), .A3(new_n1157), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1157), .A2(new_n620), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1131), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1956), .B1(new_n1035), .B2(new_n1000), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1150), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT61), .A3(new_n1138), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .A4(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1076), .A2(G1996), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT58), .B(G1341), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1000), .B2(new_n1047), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n554), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1151), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1129), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1125), .B1(new_n1037), .B2(G286), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1173), .A2(new_n1127), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1125), .B1(new_n1122), .B2(G8), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT62), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1118), .A2(G171), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1128), .B(new_n1178), .C1(new_n1127), .C2(new_n1173), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1044), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1172), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1079), .A2(G8), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1072), .B1(KEYINPUT119), .B2(G8), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1186), .A2(new_n1069), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1099), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(G290), .B(G1986), .Z(new_n1189));
  OAI21_X1  g764(.A(new_n1017), .B1(new_n1001), .B2(new_n1189), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT115), .Z(new_n1191));
  OAI21_X1  g766(.A(new_n1020), .B1(new_n1188), .B2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g767(.A1(new_n660), .A2(G319), .A3(new_n673), .ZN(new_n1194));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g770(.A1(new_n660), .A2(G319), .A3(KEYINPUT127), .A4(new_n673), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n909), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n980), .A2(new_n977), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1200), .A2(KEYINPUT43), .ZN(new_n1201));
  AOI211_X1 g775(.A(G229), .B(new_n1199), .C1(new_n1201), .C2(new_n978), .ZN(G308));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n978), .ZN(new_n1203));
  NAND4_X1  g777(.A1(new_n1203), .A2(new_n694), .A3(new_n909), .A4(new_n1198), .ZN(G225));
endmodule


