//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT78), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(G107), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n202));
  OAI211_X1 g016(.A(G104), .B(new_n198), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n197), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n194), .A2(new_n196), .A3(G107), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n200), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT67), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(new_n211), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n213), .A2(new_n215), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n217), .A2(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT80), .B1(new_n209), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n219), .B1(new_n218), .B2(new_n211), .ZN(new_n227));
  AND4_X1   g041(.A1(new_n219), .A2(new_n211), .A3(new_n213), .A4(new_n215), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT78), .B(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(new_n231), .B2(G107), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n232), .A2(new_n207), .A3(new_n203), .A4(new_n206), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n229), .A2(new_n230), .A3(new_n233), .A4(new_n200), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT10), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G137), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n239), .A2(new_n241), .A3(KEYINPUT11), .A4(G134), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT65), .A2(G134), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(G137), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(G137), .B1(new_n245), .B2(new_n246), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n242), .B(new_n247), .C1(new_n248), .C2(KEYINPUT11), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT65), .A2(G134), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT65), .A2(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n238), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(new_n247), .A4(new_n242), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n203), .B(new_n206), .C1(new_n197), .C2(new_n204), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G101), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n218), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n214), .A2(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n212), .B2(G143), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n214), .A2(KEYINPUT64), .A3(G146), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT0), .B(G128), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n260), .A2(G101), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n233), .A3(KEYINPUT4), .ZN(new_n275));
  OAI211_X1 g089(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n214), .C2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G128), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT68), .B1(new_n213), .B2(KEYINPUT1), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT69), .B1(new_n279), .B2(new_n269), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n217), .A2(new_n220), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n267), .A2(new_n268), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n213), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n283), .B(new_n284), .C1(new_n278), .C2(new_n277), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(KEYINPUT10), .B(new_n200), .C1(new_n205), .C2(new_n208), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n273), .A2(new_n275), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n237), .A2(new_n259), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G140), .ZN(new_n291));
  INV_X1    g105(.A(G953), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n292), .A2(G227), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n291), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n286), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n296), .A2(new_n209), .B1(new_n225), .B2(new_n234), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT12), .B1(new_n258), .B2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n297), .A2(new_n259), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n299), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(G143), .B2(new_n212), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n210), .B1(new_n303), .B2(KEYINPUT68), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n221), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n269), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n307), .A2(new_n284), .B1(new_n220), .B2(new_n217), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n280), .A3(new_n209), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n235), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n301), .B1(new_n310), .B2(new_n258), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n290), .B(new_n295), .C1(new_n300), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n286), .A2(new_n288), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n260), .A2(G101), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT4), .B1(new_n205), .B2(new_n208), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n272), .B(new_n262), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT10), .B1(new_n225), .B2(new_n234), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n258), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n290), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n294), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G469), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n191), .ZN(new_n324));
  NAND2_X1  g138(.A1(G469), .A2(G902), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n317), .A2(new_n318), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n294), .B1(new_n327), .B2(new_n259), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n319), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n299), .B1(new_n297), .B2(new_n259), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n310), .A2(new_n258), .A3(new_n301), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n330), .A2(new_n331), .B1(new_n259), .B2(new_n327), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n329), .B1(new_n332), .B2(new_n295), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT82), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n329), .B(new_n335), .C1(new_n332), .C2(new_n295), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(G469), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n192), .B1(new_n326), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G214), .B1(G237), .B2(G902), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G116), .B(G119), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT5), .ZN(new_n342));
  INV_X1    g156(.A(G116), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n343), .A2(KEYINPUT5), .A3(G119), .ZN(new_n344));
  INV_X1    g158(.A(G113), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT2), .B(G113), .Z(new_n347));
  AOI22_X1  g161(.A1(new_n342), .A2(new_n346), .B1(new_n347), .B2(new_n341), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n233), .A2(new_n200), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n314), .A2(new_n315), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n347), .B(new_n341), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n262), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n349), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G122), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n354), .B(new_n349), .C1(new_n350), .C2(new_n352), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n359), .A3(new_n355), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n264), .B(G125), .C1(new_n269), .C2(new_n270), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G125), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n286), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G224), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n366), .B(new_n362), .C1(new_n286), .C2(new_n363), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n360), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT83), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n358), .A2(new_n370), .A3(new_n373), .A4(new_n360), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n367), .A2(KEYINPUT7), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n209), .B(new_n348), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n354), .B(KEYINPUT8), .Z(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n357), .B1(new_n364), .B2(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n191), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT84), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n382), .B1(new_n372), .B2(new_n374), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n387), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n340), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n292), .A3(G214), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(G143), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n256), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n394), .B(new_n214), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT18), .A3(G131), .ZN(new_n399));
  XNOR2_X1  g213(.A(G125), .B(G140), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n212), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n400), .A2(KEYINPUT16), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n363), .A2(KEYINPUT16), .A3(G140), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(G146), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n398), .A2(KEYINPUT17), .A3(G131), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n398), .A2(G131), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n395), .A2(new_n256), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n415), .A2(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n193), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n420), .A2(KEYINPUT87), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n406), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n191), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n405), .A2(new_n404), .B1(new_n412), .B2(new_n416), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT88), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n406), .A2(new_n417), .ZN(new_n427));
  INV_X1    g241(.A(new_n421), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n191), .A4(new_n422), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n426), .A2(G475), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n407), .A2(G146), .A3(new_n408), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n415), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n400), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(KEYINPUT19), .Z(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n212), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n419), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n406), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n440), .B(new_n441), .C1(new_n424), .C2(new_n420), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT20), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n427), .A2(new_n419), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n440), .A4(new_n441), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n432), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n214), .A2(KEYINPUT13), .A3(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT90), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n210), .A2(G143), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n210), .A2(G143), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n450), .B(new_n451), .C1(KEYINPUT13), .C2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n449), .A2(KEYINPUT90), .ZN(new_n454));
  OAI21_X1  g268(.A(G134), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n245), .A2(new_n246), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n214), .A2(G128), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n451), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n343), .A2(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT89), .B(G122), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(new_n343), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(G107), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(G107), .ZN(new_n463));
  OAI221_X1 g277(.A(new_n455), .B1(new_n456), .B2(new_n458), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n459), .B(KEYINPUT14), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n460), .A2(new_n343), .ZN(new_n466));
  OAI21_X1  g280(.A(G107), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n458), .B(new_n456), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n467), .B(new_n468), .C1(G107), .C2(new_n461), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n190), .A2(G217), .A3(new_n292), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n471), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n478), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G952), .ZN(new_n482));
  AOI211_X1 g296(.A(G953), .B(new_n482), .C1(G234), .C2(G237), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n191), .B(new_n292), .C1(G234), .C2(G237), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(G898), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n448), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n338), .A2(new_n392), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G234), .ZN(new_n489));
  OAI21_X1  g303(.A(G217), .B1(new_n489), .B2(G902), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT74), .ZN(new_n491));
  INV_X1    g305(.A(G119), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G128), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n210), .A2(G119), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT24), .B(G110), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT76), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n500));
  INV_X1    g314(.A(new_n494), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n493), .B(new_n500), .C1(new_n501), .C2(KEYINPUT23), .ZN(new_n502));
  OR3_X1    g316(.A1(new_n502), .A2(KEYINPUT75), .A3(G110), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT75), .B1(new_n502), .B2(G110), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n499), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n400), .A2(new_n212), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n433), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n502), .A2(G110), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n495), .B2(new_n496), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n410), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT22), .B(G137), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n187), .A2(new_n489), .A3(G953), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n511), .B(new_n512), .Z(new_n513));
  XNOR2_X1  g327(.A(new_n510), .B(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n514), .A2(KEYINPUT25), .A3(new_n191), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT25), .B1(new_n514), .B2(new_n191), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n491), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n491), .A2(G902), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n521));
  INV_X1    g335(.A(G472), .ZN(new_n522));
  AOI21_X1  g336(.A(G134), .B1(new_n239), .B2(new_n241), .ZN(new_n523));
  OAI21_X1  g337(.A(G131), .B1(new_n523), .B2(new_n248), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n257), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(new_n308), .B2(new_n280), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n271), .B1(new_n250), .B2(new_n257), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n526), .A2(new_n351), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n351), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n257), .A2(new_n524), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n286), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n527), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT28), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n535));
  NAND3_X1  g349(.A1(new_n393), .A2(new_n292), .A3(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(new_n532), .A3(new_n529), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT29), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n258), .B2(new_n272), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n531), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT70), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT70), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n531), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n286), .A2(new_n530), .B1(new_n258), .B2(new_n272), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n351), .B1(new_n552), .B2(KEYINPUT30), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n528), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n544), .B1(new_n555), .B2(new_n539), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n351), .B1(new_n526), .B2(new_n527), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n541), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT28), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT29), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n562), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI211_X1 g378(.A(new_n521), .B(new_n522), .C1(new_n556), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n531), .A2(new_n532), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n545), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n546), .A2(new_n531), .A3(new_n549), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n549), .B1(new_n546), .B2(new_n531), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n568), .B(new_n351), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n539), .B1(new_n571), .B2(new_n541), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n541), .A2(new_n542), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n539), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n542), .B1(new_n557), .B2(new_n541), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n562), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n191), .B(new_n566), .C1(new_n572), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT73), .B1(new_n577), .B2(G472), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n565), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n553), .B1(new_n550), .B2(new_n548), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n541), .A2(new_n539), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT31), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n573), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n540), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT31), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n571), .A2(new_n585), .A3(new_n539), .A4(new_n541), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G472), .A2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT32), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT32), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n591), .A3(new_n588), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n520), .B1(new_n579), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n488), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  INV_X1    g410(.A(new_n520), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n338), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n589), .A2(KEYINPUT92), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n587), .A2(new_n191), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n522), .B1(new_n600), .B2(KEYINPUT91), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n587), .A2(new_n602), .A3(new_n191), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n601), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n598), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n384), .A2(KEYINPUT93), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT93), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n390), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n386), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n476), .A2(G902), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n472), .B2(new_n474), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n472), .A2(new_n615), .A3(new_n474), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT94), .B1(new_n475), .B2(G478), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n618), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT94), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n613), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n448), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n486), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n610), .B1(new_n375), .B2(new_n383), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n340), .B1(new_n628), .B2(new_n385), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n612), .A2(new_n626), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n193), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n612), .A2(new_n629), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n443), .A2(new_n446), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n442), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n432), .A2(new_n639), .A3(new_n481), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n486), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n636), .B1(new_n637), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n612), .A2(new_n642), .A3(new_n629), .A4(KEYINPUT97), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n608), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n198), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(new_n607), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n604), .ZN(new_n652));
  INV_X1    g466(.A(new_n513), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n510), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n518), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n517), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n338), .A2(new_n392), .A3(new_n487), .A4(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NAND2_X1  g475(.A1(new_n577), .A2(G472), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n521), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n577), .A2(KEYINPUT73), .A3(G472), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n591), .B1(new_n587), .B2(new_n588), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n587), .A2(new_n591), .A3(new_n588), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n338), .A3(new_n657), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n484), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n483), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n641), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n612), .A2(new_n629), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n210), .ZN(G30));
  XNOR2_X1  g491(.A(new_n672), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n338), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT40), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n679), .B(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n389), .A2(new_n391), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT38), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n559), .A2(new_n560), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n191), .B1(new_n689), .B2(new_n539), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n555), .A2(new_n540), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n666), .B2(new_n665), .ZN(new_n693));
  INV_X1    g507(.A(new_n657), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n448), .A2(new_n481), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n339), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n683), .A2(new_n685), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n214), .ZN(G45));
  NAND4_X1  g513(.A1(new_n448), .A2(new_n621), .A3(new_n624), .A4(new_n672), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n612), .A3(new_n629), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n668), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n212), .ZN(G48));
  NAND2_X1  g518(.A1(new_n330), .A2(new_n331), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n705), .A2(new_n328), .B1(new_n320), .B2(new_n294), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT100), .ZN(new_n708));
  INV_X1    g522(.A(new_n192), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n324), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n707), .A2(new_n324), .A3(new_n709), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n667), .A2(new_n597), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n630), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT41), .B(G113), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  AOI21_X1  g530(.A(new_n713), .B1(new_n644), .B2(new_n645), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT101), .B(G116), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G18));
  NAND3_X1  g533(.A1(new_n667), .A2(new_n487), .A3(new_n657), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n612), .A2(new_n712), .A3(new_n629), .A4(new_n710), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n492), .ZN(G21));
  AND3_X1   g537(.A1(new_n612), .A2(new_n629), .A3(new_n695), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n712), .A2(new_n627), .A3(new_n710), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n522), .B1(new_n587), .B2(new_n191), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n561), .A2(new_n573), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n582), .B(new_n586), .C1(new_n729), .C2(new_n539), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n728), .A2(KEYINPUT102), .B1(new_n730), .B2(new_n588), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n597), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(KEYINPUT103), .A3(new_n597), .A4(new_n733), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n726), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n738), .B(G122), .Z(G24));
  NAND4_X1  g553(.A1(new_n731), .A2(new_n701), .A3(new_n657), .A4(new_n733), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n721), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n363), .ZN(G27));
  OR2_X1    g556(.A1(new_n594), .A2(KEYINPUT107), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n329), .B(G469), .C1(new_n332), .C2(new_n295), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n325), .B(KEYINPUT104), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n324), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT105), .B1(new_n746), .B2(new_n709), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n389), .A2(new_n339), .A3(new_n391), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n746), .A2(new_n709), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT105), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n594), .A2(KEYINPUT107), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n700), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n743), .A2(new_n752), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n594), .A2(new_n749), .A3(new_n701), .A4(new_n751), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(KEYINPUT106), .A3(new_n754), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT106), .B1(new_n757), .B2(new_n754), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  NAND4_X1  g575(.A1(new_n594), .A2(new_n749), .A3(new_n674), .A4(new_n751), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  INV_X1    g577(.A(new_n448), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n621), .A3(new_n624), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n765), .B2(KEYINPUT108), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n767), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n652), .A3(new_n657), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n334), .B2(new_n336), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  OAI21_X1  g592(.A(G469), .B1(new_n333), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n745), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT46), .B(new_n745), .C1(new_n777), .C2(new_n779), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n324), .A3(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(new_n709), .A3(new_n678), .ZN(new_n785));
  INV_X1    g599(.A(new_n748), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n773), .A2(new_n774), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XOR2_X1   g602(.A(KEYINPUT110), .B(G137), .Z(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(G39));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n709), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n784), .A2(new_n709), .A3(new_n792), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n748), .A2(new_n597), .A3(new_n700), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n593), .A3(new_n579), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NAND2_X1  g613(.A1(new_n736), .A2(new_n737), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n772), .A3(new_n483), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT50), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n712), .A2(new_n710), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n340), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n807), .B2(new_n687), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n688), .A2(KEYINPUT117), .A3(new_n340), .A4(new_n806), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n802), .A2(new_n804), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n808), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(new_n801), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n806), .A2(new_n786), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n766), .A2(KEYINPUT109), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n671), .B(new_n814), .C1(new_n817), .C2(new_n767), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n730), .A2(new_n588), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n727), .B2(new_n732), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n727), .A2(new_n732), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n694), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n814), .A2(new_n520), .A3(new_n671), .A4(new_n693), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n448), .B1(new_n621), .B2(new_n624), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n818), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n810), .A2(new_n813), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n801), .A2(new_n748), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n707), .A2(new_n324), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n794), .B(new_n795), .C1(new_n709), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT116), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n829), .A3(KEYINPUT116), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n743), .A2(new_n753), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n818), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT48), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(KEYINPUT119), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n801), .A2(new_n721), .ZN(new_n838));
  AOI211_X1 g652(.A(new_n482), .B(G953), .C1(new_n823), .C2(new_n626), .ZN(new_n839));
  XNOR2_X1  g653(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n818), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n827), .A2(new_n829), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT51), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n845), .B2(new_n826), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT120), .B1(new_n833), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n826), .A2(new_n845), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n842), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n850));
  INV_X1    g664(.A(new_n832), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n826), .A2(new_n851), .A3(new_n830), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n849), .B(new_n850), .C1(KEYINPUT51), .C2(new_n852), .ZN(new_n853));
  OAI22_X1  g667(.A1(new_n713), .A2(new_n630), .B1(new_n720), .B2(new_n721), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n738), .A2(new_n717), .A3(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n481), .A2(new_n432), .A3(new_n447), .A4(new_n627), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n686), .A2(new_n339), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n392), .A2(KEYINPUT112), .A3(new_n856), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n392), .A2(new_n627), .A3(new_n626), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n608), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n595), .B1(new_n658), .B2(new_n652), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n740), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n752), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n667), .A2(new_n338), .A3(new_n657), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n481), .A2(new_n673), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n432), .A2(new_n869), .A3(new_n639), .A4(new_n640), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n339), .A3(new_n391), .A4(new_n389), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT113), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n786), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n867), .A2(new_n875), .A3(new_n762), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n760), .A2(new_n855), .A3(new_n865), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n740), .A2(new_n721), .B1(new_n668), .B2(new_n675), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n750), .A2(new_n693), .A3(new_n694), .A4(new_n672), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n612), .A2(new_n629), .A3(new_n695), .ZN(new_n883));
  OAI22_X1  g697(.A1(new_n668), .A2(new_n702), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT52), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n880), .B2(new_n884), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n879), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n879), .A3(new_n888), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n878), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT53), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n886), .A2(new_n888), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n878), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(KEYINPUT54), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n717), .A2(new_n854), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n738), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n855), .A2(KEYINPUT115), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n760), .A2(new_n876), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n862), .A2(new_n608), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n659), .A2(new_n905), .A3(KEYINPUT53), .A4(new_n595), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n886), .B2(new_n888), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n895), .A2(KEYINPUT114), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n877), .B1(new_n909), .B2(new_n890), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n898), .B(new_n908), .C1(new_n910), .C2(KEYINPUT53), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n847), .A2(new_n853), .A3(new_n897), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(G952), .B2(G953), .ZN(new_n913));
  NOR4_X1   g727(.A1(new_n765), .A2(new_n520), .A3(new_n340), .A4(new_n192), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n828), .A2(KEYINPUT49), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n828), .A2(KEYINPUT49), .ZN(new_n917));
  OR4_X1    g731(.A1(new_n687), .A2(new_n916), .A3(new_n693), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n913), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n292), .A2(G952), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n358), .A2(new_n360), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n370), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n908), .B1(new_n910), .B2(KEYINPUT53), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(G210), .A3(G902), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n923), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT121), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n925), .A2(new_n930), .A3(new_n926), .A4(new_n923), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n920), .B(new_n927), .C1(new_n929), .C2(new_n931), .ZN(G51));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n911), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n891), .A2(new_n889), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n894), .B1(new_n935), .B2(new_n877), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n936), .A2(KEYINPUT122), .A3(new_n898), .A4(new_n908), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n924), .A2(KEYINPUT54), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n745), .B(KEYINPUT57), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n322), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n924), .A2(G902), .A3(new_n780), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n920), .B1(new_n942), .B2(new_n943), .ZN(G54));
  AND2_X1   g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n924), .A2(G902), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n444), .A2(new_n440), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n920), .ZN(new_n949));
  INV_X1    g763(.A(new_n947), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n924), .A2(G902), .A3(new_n950), .A4(new_n945), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT123), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n948), .A2(new_n954), .A3(new_n949), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G60));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT59), .Z(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n897), .B2(new_n911), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n949), .B1(new_n959), .B2(new_n622), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n617), .B2(new_n618), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n939), .B2(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT124), .Z(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT60), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n924), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n514), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n924), .A2(new_n655), .A3(new_n965), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n949), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G66));
  OAI21_X1  g786(.A(G953), .B1(new_n485), .B2(new_n365), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n855), .A2(new_n865), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n921), .B1(G898), .B2(new_n292), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  NAND2_X1  g791(.A1(new_n551), .A2(new_n568), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n437), .ZN(new_n979));
  INV_X1    g793(.A(new_n703), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n881), .A2(new_n980), .ZN(new_n981));
  OR3_X1    g795(.A1(new_n698), .A2(KEYINPUT62), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n626), .B1(new_n481), .B2(new_n764), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n983), .A2(new_n679), .A3(new_n748), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n594), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n982), .A2(new_n788), .A3(new_n798), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT62), .B1(new_n698), .B2(new_n981), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n987), .A2(KEYINPUT125), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(KEYINPUT125), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n979), .B1(new_n990), .B2(G953), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n292), .B1(G227), .B2(G900), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n788), .A2(new_n798), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n834), .A2(new_n785), .A3(new_n724), .ZN(new_n996));
  AND4_X1   g810(.A1(new_n980), .A2(new_n996), .A3(new_n762), .A4(new_n881), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n995), .A2(new_n292), .A3(new_n760), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n979), .B1(G900), .B2(G953), .ZN(new_n999));
  AOI22_X1  g813(.A1(new_n998), .A2(new_n999), .B1(new_n993), .B2(new_n992), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n991), .A2(new_n994), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n994), .B1(new_n991), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(G72));
  NOR3_X1   g817(.A1(new_n580), .A2(new_n539), .A3(new_n528), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n691), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  AND4_X1   g821(.A1(new_n893), .A2(new_n896), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1007), .B(KEYINPUT127), .Z(new_n1009));
  OAI21_X1  g823(.A(new_n949), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n990), .A2(new_n691), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n995), .A2(new_n760), .A3(new_n997), .A4(new_n1004), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n1008), .B(new_n1010), .C1(new_n1013), .C2(new_n974), .ZN(G57));
endmodule


