//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT95), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n203), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n212));
  AOI21_X1  g011(.A(G36gat), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n210), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n214));
  OR3_X1    g013(.A1(new_n213), .A2(KEYINPUT15), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT15), .B1(new_n213), .B2(new_n214), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT17), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n208), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n206), .B(G8gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n220), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n220), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT96), .B1(new_n208), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n224), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n226), .B(KEYINPUT13), .Z(new_n231));
  NAND3_X1  g030(.A1(new_n223), .A2(KEYINPUT96), .A3(new_n220), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n224), .A2(new_n222), .A3(new_n226), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n227), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G197gat), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT11), .B(G169gat), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n241), .B(KEYINPUT12), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT97), .ZN(new_n244));
  INV_X1    g043(.A(new_n242), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n227), .A2(new_n233), .A3(new_n245), .A4(new_n236), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n237), .A2(KEYINPUT97), .A3(new_n242), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G141gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G148gat), .ZN(new_n251));
  INV_X1    g050(.A(G148gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G141gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT2), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G155gat), .ZN(new_n258));
  INV_X1    g057(.A(G162gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT79), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n260), .A2(new_n263), .A3(new_n255), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n257), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT82), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT80), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n252), .A2(G141gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n270), .A3(new_n261), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n258), .A2(KEYINPUT81), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G155gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n272), .B1(new_n276), .B2(G162gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n266), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT81), .B(G155gat), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT2), .B1(new_n279), .B2(new_n259), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n269), .A2(new_n268), .B1(new_n260), .B2(new_n255), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n280), .A2(KEYINPUT82), .A3(new_n267), .A4(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n265), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G120gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(new_n284), .B2(new_n285), .ZN(new_n287));
  OR2_X1    g086(.A1(G127gat), .A2(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(G127gat), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT70), .B(G134gat), .Z(new_n290));
  OAI211_X1 g089(.A(new_n287), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT71), .B(G113gat), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n286), .B(new_n292), .C1(new_n293), .C2(new_n285), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n283), .A2(KEYINPUT4), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT4), .B1(new_n283), .B2(new_n296), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n282), .ZN(new_n300));
  INV_X1    g099(.A(new_n265), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT3), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT83), .B1(new_n283), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n296), .B1(new_n283), .B2(new_n305), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n299), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n295), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n283), .A2(new_n296), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n309), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n283), .A2(KEYINPUT4), .A3(new_n296), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n318), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n322), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n297), .A2(new_n298), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT84), .B1(new_n327), .B2(new_n308), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n317), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT0), .ZN(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n324), .B1(new_n318), .B2(new_n323), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(KEYINPUT84), .A3(new_n308), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n336), .A2(new_n337), .B1(new_n310), .B2(new_n316), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n333), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n337), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n333), .B1(new_n343), .B2(new_n317), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n344), .B2(KEYINPUT6), .ZN(new_n345));
  NOR4_X1   g144(.A1(new_n338), .A2(KEYINPUT85), .A3(new_n340), .A4(new_n333), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n352), .B(KEYINPUT75), .Z(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT26), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n354), .B(new_n357), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT27), .B(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(G190gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT68), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n364), .B2(new_n365), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n363), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT65), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n354), .A2(KEYINPUT24), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT24), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(G183gat), .A3(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n372), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI211_X1 g178(.A(KEYINPUT65), .B(new_n377), .C1(new_n373), .C2(new_n375), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT66), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n358), .B1(new_n361), .B2(KEYINPUT23), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n384), .A2(G169gat), .A3(G176gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n382), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n361), .A2(KEYINPUT23), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n384), .B1(G169gat), .B2(G176gat), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(KEYINPUT66), .A3(new_n388), .A4(new_n358), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT25), .B1(new_n381), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n387), .A2(KEYINPUT25), .A3(new_n388), .A4(new_n358), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT67), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n376), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n371), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n353), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G197gat), .B(G204gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(G211gat), .A2(G218gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G211gat), .B(G218gat), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(G197gat), .A2(G204gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n406), .A2(new_n407), .B1(new_n400), .B2(new_n399), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n403), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n353), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n376), .A2(new_n378), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT65), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n376), .A2(new_n372), .A3(new_n378), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n386), .A4(new_n389), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT25), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n394), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G183gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT27), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT27), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G183gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n424), .A3(new_n365), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(KEYINPUT68), .A3(new_n366), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n362), .B1(new_n426), .B2(new_n368), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT69), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI211_X1 g228(.A(KEYINPUT69), .B(new_n362), .C1(new_n426), .C2(new_n368), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n412), .B1(new_n420), .B2(new_n431), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n397), .A2(new_n411), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n420), .A2(new_n353), .A3(new_n371), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n353), .A2(KEYINPUT29), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n371), .A2(KEYINPUT69), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n428), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n394), .B1(new_n416), .B2(new_n417), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(new_n440), .A3(new_n411), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n351), .B1(new_n433), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n353), .B1(new_n438), .B2(new_n439), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n420), .B2(new_n371), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n410), .B(new_n444), .C1(new_n445), .C2(new_n353), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n446), .A2(KEYINPUT30), .A3(new_n441), .A4(new_n350), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n446), .A2(new_n441), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT76), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT30), .A4(new_n350), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT77), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT77), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n457));
  NAND2_X1  g256(.A1(new_n446), .A2(new_n441), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(new_n351), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n347), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G78gat), .B(G106gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G22gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G228gat), .ZN(new_n464));
  INV_X1    g263(.A(G233gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT29), .B1(new_n405), .B2(new_n409), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT3), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n402), .A2(new_n404), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n408), .A2(new_n403), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n396), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT88), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n302), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n300), .A2(new_n305), .A3(new_n301), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n396), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n476), .A2(KEYINPUT89), .B1(new_n478), .B2(new_n411), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n283), .B1(new_n470), .B2(new_n474), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n467), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n405), .A2(KEYINPUT87), .ZN(new_n484));
  OR3_X1    g283(.A1(new_n408), .A2(KEYINPUT87), .A3(new_n403), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n409), .A2(KEYINPUT86), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n408), .A2(new_n487), .A3(new_n403), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT3), .B1(new_n489), .B2(new_n396), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n467), .B1(new_n490), .B2(new_n283), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT29), .B1(new_n283), .B2(new_n305), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(new_n410), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n483), .A2(KEYINPUT90), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n480), .A2(new_n481), .B1(new_n492), .B2(new_n410), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n476), .A2(KEYINPUT89), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n466), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n494), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G50gat), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n495), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n502), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT90), .B1(new_n483), .B2(new_n494), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n496), .A3(new_n500), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n463), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n420), .A2(new_n295), .A3(new_n431), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n296), .B1(new_n438), .B2(new_n439), .ZN(new_n510));
  NAND2_X1  g309(.A1(G227gat), .A2(G233gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n511), .B(KEYINPUT64), .Z(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT72), .A4(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT32), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n512), .B1(new_n509), .B2(new_n510), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT34), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT33), .B1(new_n515), .B2(new_n516), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G15gat), .B(G43gat), .Z(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G71gat), .B(G99gat), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  AOI21_X1  g327(.A(new_n521), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n519), .B(KEYINPUT34), .ZN(new_n530));
  INV_X1    g329(.A(new_n528), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n530), .A2(new_n522), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n518), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n502), .B1(new_n495), .B2(new_n501), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n505), .A2(new_n506), .A3(new_n504), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n462), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n523), .A2(new_n521), .A3(new_n528), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n530), .B1(new_n522), .B2(new_n531), .ZN(new_n538));
  INV_X1    g337(.A(new_n518), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n508), .A2(new_n533), .A3(new_n536), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n460), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT94), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n544), .B(KEYINPUT35), .C1(new_n460), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n539), .B1(new_n537), .B2(new_n538), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n533), .A2(KEYINPUT93), .A3(new_n540), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n347), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n452), .A2(new_n459), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n508), .A2(new_n553), .A3(new_n554), .A4(new_n536), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n299), .A2(new_n308), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n315), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT39), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(new_n334), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n560), .B(KEYINPUT39), .C1(new_n315), .C2(new_n314), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(KEYINPUT40), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n335), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n536), .B(new_n508), .C1(new_n568), .C2(new_n553), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n434), .A2(new_n440), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(new_n410), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n411), .B(new_n444), .C1(new_n445), .C2(new_n353), .ZN(new_n574));
  AOI211_X1 g373(.A(KEYINPUT38), .B(new_n350), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n449), .A2(new_n571), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n575), .A2(new_n576), .B1(new_n449), .B2(new_n350), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n341), .C1(new_n345), .C2(new_n346), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT85), .B1(new_n335), .B2(new_n340), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n344), .A2(new_n342), .A3(KEYINPUT6), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n583), .A2(KEYINPUT91), .A3(new_n341), .A4(new_n577), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n350), .B1(new_n458), .B2(KEYINPUT37), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n585), .A2(KEYINPUT92), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(KEYINPUT92), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n576), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT38), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n580), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n508), .A2(new_n536), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(new_n548), .B2(new_n549), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n533), .A2(KEYINPUT36), .A3(new_n540), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n460), .A2(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n249), .B1(new_n558), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n347), .ZN(new_n599));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT98), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT9), .ZN(new_n602));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603));
  INV_X1    g402(.A(G71gat), .ZN(new_n604));
  INV_X1    g403(.A(G78gat), .ZN(new_n605));
  OAI221_X1 g404(.A(new_n601), .B1(new_n602), .B2(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT99), .ZN(new_n607));
  AND2_X1   g406(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(G64gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(G64gat), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n602), .A2(G71gat), .A3(G78gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n604), .A2(new_n605), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n289), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n607), .A2(new_n613), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n223), .B1(KEYINPUT21), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n618), .B(G127gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n258), .ZN(new_n628));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n622), .A2(new_n625), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n637));
  INV_X1    g436(.A(G85gat), .ZN(new_n638));
  INV_X1    g437(.A(G92gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(KEYINPUT8), .A2(new_n643), .B1(new_n638), .B2(new_n639), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G99gat), .B(G106gat), .Z(new_n646));
  OR2_X1    g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n645), .A2(KEYINPUT103), .A3(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n221), .ZN(new_n654));
  AND2_X1   g453(.A1(G232gat), .A2(G233gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n652), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(KEYINPUT104), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(KEYINPUT104), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n636), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n655), .A2(KEYINPUT41), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT101), .ZN(new_n664));
  XOR2_X1   g463(.A(G134gat), .B(G162gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n658), .A2(new_n636), .A3(new_n659), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n661), .A2(new_n662), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n666), .B(KEYINPUT105), .ZN(new_n669));
  INV_X1    g468(.A(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n660), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n649), .A2(KEYINPUT106), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n647), .B1(KEYINPUT106), .B2(new_n649), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n620), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n652), .A2(new_n614), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT10), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n620), .A2(KEYINPUT10), .A3(new_n652), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n673), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  INV_X1    g481(.A(new_n673), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(G120gat), .B(G148gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(G176gat), .B(G204gat), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n686), .B(new_n687), .Z(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n681), .A2(new_n684), .A3(new_n688), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n634), .A2(new_n672), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n598), .A2(new_n599), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G1gat), .ZN(G1324gat));
  INV_X1    g495(.A(new_n553), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n598), .A2(new_n697), .A3(new_n694), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(G8gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT16), .B(G8gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT42), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(KEYINPUT42), .B2(new_n701), .ZN(G1325gat));
  NAND2_X1  g502(.A1(new_n598), .A2(new_n694), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n594), .A2(new_n595), .ZN(new_n705));
  OAI21_X1  g504(.A(G15gat), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n550), .A2(new_n551), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(G15gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n704), .B2(new_n708), .ZN(G1326gat));
  INV_X1    g508(.A(new_n592), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n578), .A2(new_n579), .B1(KEYINPUT38), .B2(new_n588), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n569), .B1(new_n715), .B2(new_n584), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n460), .A2(new_n592), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n705), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n716), .A2(new_n718), .A3(KEYINPUT109), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n591), .B2(new_n596), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n558), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n672), .A2(KEYINPUT44), .ZN(new_n723));
  INV_X1    g522(.A(new_n672), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n556), .B1(new_n543), .B2(new_n545), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n716), .A2(new_n718), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n722), .A2(new_n723), .B1(new_n727), .B2(KEYINPUT44), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n692), .B(KEYINPUT108), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n249), .A3(new_n634), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n714), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n558), .A2(new_n597), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n724), .ZN(new_n736));
  INV_X1    g535(.A(new_n723), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n716), .B2(new_n718), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n591), .A2(new_n720), .A3(new_n596), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n737), .B1(new_n740), .B2(new_n558), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT110), .B(new_n731), .C1(new_n736), .C2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n733), .A2(new_n599), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n210), .B1(new_n743), .B2(KEYINPUT111), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT111), .B2(new_n743), .ZN(new_n745));
  INV_X1    g544(.A(new_n692), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n634), .A2(new_n672), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n598), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n599), .A2(new_n210), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n748), .A2(KEYINPUT107), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n745), .A2(new_n753), .ZN(G1328gat));
  NAND3_X1  g553(.A1(new_n733), .A2(new_n697), .A3(new_n742), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G36gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n748), .A2(G36gat), .A3(new_n553), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(G1329gat));
  INV_X1    g559(.A(new_n705), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n733), .A2(new_n761), .A3(new_n742), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n707), .A2(G43gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n598), .A2(new_n747), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n761), .B(new_n731), .C1(new_n736), .C2(new_n741), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G43gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n766), .B1(new_n772), .B2(new_n765), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n769), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n767), .B1(new_n762), .B2(G43gat), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT113), .B1(new_n776), .B2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1330gat));
  NOR3_X1   g577(.A1(new_n748), .A2(G50gat), .A3(new_n710), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n733), .A2(new_n592), .A3(new_n742), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(G50gat), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n782));
  NAND2_X1  g581(.A1(new_n727), .A2(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n725), .B1(new_n738), .B2(new_n739), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n737), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n592), .A3(new_n731), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n786), .A2(G50gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n779), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n781), .A2(new_n782), .B1(new_n787), .B2(new_n789), .ZN(G1331gat));
  NAND4_X1  g589(.A1(new_n730), .A2(new_n249), .A3(new_n634), .A4(new_n672), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n784), .A2(KEYINPUT115), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT115), .B1(new_n784), .B2(new_n791), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n599), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G57gat), .ZN(G1332gat));
  OAI22_X1  g596(.A1(new_n794), .A2(new_n553), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n697), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT49), .B(G64gat), .Z(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT116), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n798), .B(new_n803), .C1(new_n799), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1333gat));
  OAI21_X1  g604(.A(G71gat), .B1(new_n794), .B2(new_n705), .ZN(new_n806));
  INV_X1    g605(.A(new_n707), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n604), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n794), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(G1334gat));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n710), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(new_n605), .ZN(G1335gat));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  INV_X1    g613(.A(new_n249), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n634), .A2(new_n815), .A3(new_n692), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n785), .A2(new_n599), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n785), .A2(new_n819), .A3(new_n599), .A4(new_n816), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n818), .A2(new_n820), .A3(G85gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n746), .A2(new_n599), .A3(new_n638), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT118), .B1(new_n784), .B2(new_n672), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n722), .A2(new_n824), .A3(new_n724), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n634), .A2(new_n815), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n823), .A2(new_n825), .A3(KEYINPUT51), .A4(new_n826), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n822), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n814), .B1(new_n821), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n818), .A2(new_n820), .A3(G85gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n830), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n833), .B(KEYINPUT119), .C1(new_n835), .C2(new_n822), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n836), .ZN(G1336gat));
  NOR2_X1   g636(.A1(new_n553), .A2(G92gat), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n729), .B(new_n839), .C1(new_n829), .C2(new_n830), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n785), .A2(new_n816), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n639), .B1(new_n841), .B2(new_n697), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT52), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n834), .A2(new_n730), .A3(new_n838), .ZN(new_n844));
  INV_X1    g643(.A(new_n842), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(G1337gat));
  INV_X1    g647(.A(G99gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n807), .A2(new_n849), .A3(new_n746), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n841), .A2(new_n761), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n835), .A2(new_n850), .B1(new_n851), .B2(new_n849), .ZN(G1338gat));
  NOR2_X1   g651(.A1(new_n710), .A2(G106gat), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI211_X1 g653(.A(new_n729), .B(new_n854), .C1(new_n829), .C2(new_n830), .ZN(new_n855));
  INV_X1    g654(.A(G106gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n841), .B2(new_n592), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT53), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n834), .A2(new_n730), .A3(new_n853), .ZN(new_n859));
  INV_X1    g658(.A(new_n857), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(G1339gat));
  NOR2_X1   g662(.A1(new_n693), .A2(new_n815), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n673), .C1(new_n678), .C2(new_n680), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(new_n689), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n683), .B(new_n679), .C1(new_n682), .C2(KEYINPUT10), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(KEYINPUT54), .A3(new_n681), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n867), .A2(KEYINPUT55), .A3(new_n869), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n691), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n225), .A2(new_n226), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n241), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n246), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n668), .A2(new_n878), .A3(new_n671), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT120), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n873), .A2(new_n691), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT55), .B1(new_n867), .B2(new_n869), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n883), .A2(new_n724), .A3(new_n884), .A4(new_n878), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n883), .A2(new_n815), .B1(new_n746), .B2(new_n878), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n880), .B(new_n885), .C1(new_n886), .C2(new_n724), .ZN(new_n887));
  INV_X1    g686(.A(new_n634), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n864), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n592), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n890), .A2(new_n599), .A3(new_n553), .A4(new_n807), .ZN(new_n891));
  OAI21_X1  g690(.A(G113gat), .B1(new_n891), .B2(new_n249), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n599), .A2(new_n553), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n889), .A2(new_n541), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n293), .A3(new_n815), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1340gat));
  NOR3_X1   g695(.A1(new_n891), .A2(new_n285), .A3(new_n729), .ZN(new_n897));
  AOI21_X1  g696(.A(G120gat), .B1(new_n894), .B2(new_n746), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1341gat));
  OAI21_X1  g698(.A(G127gat), .B1(new_n891), .B2(new_n888), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n289), .A3(new_n634), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1342gat));
  NAND3_X1  g701(.A1(new_n894), .A2(new_n290), .A3(new_n724), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT56), .ZN(new_n904));
  OAI21_X1  g703(.A(G134gat), .B1(new_n891), .B2(new_n672), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(KEYINPUT56), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G1343gat));
  NOR2_X1   g706(.A1(new_n889), .A2(new_n893), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n761), .A2(new_n710), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n250), .B1(new_n910), .B2(new_n249), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n761), .A2(new_n893), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n883), .A2(new_n815), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n746), .A2(new_n878), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n724), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n885), .A2(new_n880), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n888), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n864), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n710), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n867), .A2(KEYINPUT121), .A3(new_n869), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT121), .B1(new_n867), .B2(new_n869), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT55), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n247), .A2(new_n873), .A3(new_n248), .A4(new_n691), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n915), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n672), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n880), .A3(new_n885), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n864), .B1(new_n929), .B2(new_n888), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT57), .B1(new_n930), .B2(new_n710), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n922), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n815), .A2(G141gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n911), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT58), .Z(G1344gat));
  OAI21_X1  g734(.A(KEYINPUT57), .B1(new_n889), .B2(new_n710), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n874), .A2(new_n879), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n927), .B2(new_n672), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n919), .B1(new_n938), .B2(new_n634), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n710), .A2(KEYINPUT57), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n761), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n893), .A2(new_n692), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n936), .A2(new_n941), .A3(new_n945), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G148gat), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT59), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT124), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n922), .A2(new_n931), .A3(new_n746), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n252), .A2(KEYINPUT59), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n950), .A2(KEYINPUT122), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT122), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n955), .B(KEYINPUT59), .C1(new_n944), .C2(new_n947), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n949), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n910), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n252), .A3(new_n746), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1345gat));
  OAI21_X1  g759(.A(new_n276), .B1(new_n932), .B2(new_n888), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n958), .A2(new_n279), .A3(new_n634), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1346gat));
  NOR3_X1   g762(.A1(new_n932), .A2(new_n259), .A3(new_n672), .ZN(new_n964));
  AOI21_X1  g763(.A(G162gat), .B1(new_n958), .B2(new_n724), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(new_n965), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n552), .A2(new_n553), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n890), .A2(new_n967), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(new_n355), .A3(new_n249), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n889), .A2(new_n599), .A3(new_n553), .ZN(new_n970));
  INV_X1    g769(.A(new_n541), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n815), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n969), .B1(new_n974), .B2(new_n355), .ZN(G1348gat));
  OAI21_X1  g774(.A(G176gat), .B1(new_n968), .B2(new_n729), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n746), .A2(new_n356), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n972), .B2(new_n977), .ZN(G1349gat));
  OAI21_X1  g777(.A(G183gat), .B1(new_n968), .B2(new_n888), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n634), .A2(new_n364), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n972), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n981), .B(new_n982), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n973), .A2(new_n365), .A3(new_n724), .ZN(new_n984));
  OAI21_X1  g783(.A(G190gat), .B1(new_n968), .B2(new_n672), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n985), .A2(KEYINPUT61), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(KEYINPUT61), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1351gat));
  AND2_X1   g787(.A1(new_n970), .A2(new_n909), .ZN(new_n989));
  XNOR2_X1  g788(.A(KEYINPUT126), .B(G197gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(new_n815), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n936), .A2(new_n941), .A3(new_n347), .A4(new_n697), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n992), .A2(new_n249), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n991), .B1(new_n993), .B2(new_n990), .ZN(G1352gat));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  AOI21_X1  g794(.A(G204gat), .B1(new_n995), .B2(KEYINPUT62), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n989), .A2(new_n746), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n997), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(G204gat), .B1(new_n992), .B2(new_n729), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1353gat));
  INV_X1    g800(.A(G211gat), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n989), .A2(new_n1002), .A3(new_n634), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n992), .A2(new_n888), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  INV_X1    g806(.A(G218gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n989), .A2(new_n1008), .A3(new_n724), .ZN(new_n1009));
  OAI21_X1  g808(.A(G218gat), .B1(new_n992), .B2(new_n672), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1355gat));
endmodule


