//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G140), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT88), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G140), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(G146), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT89), .ZN(new_n197));
  XNOR2_X1  g011(.A(G125), .B(G140), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n191), .A2(new_n197), .A3(G146), .A4(new_n195), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT18), .A2(G131), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(G237), .A2(G953), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n206), .A2(G143), .A3(G214), .ZN(new_n207));
  AOI21_X1  g021(.A(G143), .B1(new_n206), .B2(G214), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT86), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G237), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G214), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(G143), .A3(G214), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT86), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n205), .B1(new_n210), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT87), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(KEYINPUT87), .B(new_n205), .C1(new_n210), .C2(new_n217), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n216), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT90), .A3(new_n204), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT90), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n222), .B2(new_n205), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n203), .A2(new_n220), .A3(new_n221), .A4(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(G131), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT72), .B1(new_n192), .B2(KEYINPUT16), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT72), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT16), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n188), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT71), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n198), .A2(new_n244), .A3(KEYINPUT16), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n199), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n243), .A3(new_n245), .A4(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n222), .A2(KEYINPUT17), .A3(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n236), .A2(new_n247), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n228), .A2(new_n231), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT92), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n233), .A2(new_n234), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT19), .ZN(new_n254));
  OR2_X1    g068(.A1(new_n254), .A2(KEYINPUT91), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n191), .A2(KEYINPUT19), .A3(new_n195), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT19), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n198), .A2(KEYINPUT91), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n253), .B(new_n248), .C1(new_n259), .C2(G146), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n228), .A2(new_n252), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n231), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n252), .B1(new_n228), .B2(new_n260), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n251), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n266));
  NOR2_X1   g080(.A1(G475), .A2(G902), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT93), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n267), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT20), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT93), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n265), .A2(new_n272), .A3(new_n266), .A4(new_n267), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n228), .A2(new_n231), .A3(new_n250), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n231), .B1(new_n228), .B2(new_n250), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT94), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT94), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(G475), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G478), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT15), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT70), .B(G902), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G107), .ZN(new_n287));
  INV_X1    g101(.A(G122), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G116), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n287), .B1(new_n289), .B2(KEYINPUT14), .ZN(new_n290));
  XNOR2_X1  g104(.A(G116), .B(G122), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n214), .A2(G128), .ZN(new_n293));
  INV_X1    g107(.A(G128), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G143), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT96), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G128), .B(G143), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(KEYINPUT96), .ZN(new_n300));
  INV_X1    g114(.A(G134), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(KEYINPUT96), .ZN(new_n304));
  AOI21_X1  g118(.A(G134), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n292), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n301), .B1(new_n298), .B2(new_n300), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G122), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n289), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT95), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT95), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n291), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n287), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n299), .A2(KEYINPUT13), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n315), .B(G134), .C1(KEYINPUT13), .C2(new_n293), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(KEYINPUT95), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n291), .A2(new_n312), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G107), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n307), .A2(new_n314), .A3(new_n316), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n306), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT9), .B(G234), .ZN(new_n322));
  INV_X1    g136(.A(G217), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n322), .A2(new_n323), .A3(G953), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n306), .A2(new_n320), .A3(new_n324), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n286), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT97), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI211_X1 g144(.A(KEYINPUT97), .B(new_n286), .C1(new_n326), .C2(new_n327), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n284), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI22_X1  g146(.A1(new_n328), .A2(new_n329), .B1(KEYINPUT15), .B2(new_n283), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(G234), .A2(G237), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n335), .A2(G952), .A3(new_n212), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n286), .A2(G953), .A3(new_n335), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT21), .B(G898), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n274), .A2(new_n282), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT11), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n301), .B2(G137), .ZN(new_n344));
  INV_X1    g158(.A(G137), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT11), .A3(G134), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n301), .A2(G137), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n232), .A4(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n301), .A2(G137), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n345), .A2(G134), .ZN(new_n350));
  OAI21_X1  g164(.A(G131), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n348), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n214), .A2(KEYINPUT1), .A3(G146), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n199), .A2(G143), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n214), .A2(G146), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n356), .B1(new_n359), .B2(new_n294), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n294), .A2(KEYINPUT1), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n357), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n355), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G131), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n348), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT0), .A2(G128), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT0), .A2(G128), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n359), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G143), .B(G146), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n368), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n364), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT66), .ZN(new_n377));
  INV_X1    g191(.A(G119), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(G116), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n308), .A2(KEYINPUT66), .A3(G119), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT2), .A2(G113), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT65), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT2), .A3(G113), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT2), .A2(G113), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n381), .A2(new_n388), .A3(new_n389), .A4(new_n382), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n366), .A2(new_n348), .B1(new_n371), .B2(new_n373), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT64), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n352), .A2(new_n395), .B1(new_n360), .B2(new_n362), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n348), .A2(new_n351), .A3(KEYINPUT64), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n376), .B(new_n393), .C1(KEYINPUT30), .C2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n211), .A2(new_n212), .A3(G210), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G101), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n352), .A2(KEYINPUT67), .B1(new_n360), .B2(new_n362), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n394), .B1(new_n405), .B2(new_n355), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n391), .A2(new_n392), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT31), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n364), .A2(new_n407), .A3(new_n375), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT28), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n406), .A2(KEYINPUT28), .A3(new_n407), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n352), .A2(new_n395), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n363), .A3(new_n397), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n375), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n393), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n404), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT31), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n399), .A2(new_n408), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n410), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(G472), .A2(G902), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT32), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT32), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  INV_X1    g242(.A(new_n413), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n411), .A2(KEYINPUT69), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n364), .A2(new_n375), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n393), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n364), .A2(new_n407), .A3(new_n433), .A4(new_n375), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n429), .B1(new_n435), .B2(KEYINPUT28), .ZN(new_n436));
  INV_X1    g250(.A(new_n404), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT29), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n419), .A2(new_n437), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n399), .A2(new_n404), .A3(new_n411), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n438), .B(new_n285), .C1(new_n441), .C2(KEYINPUT29), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n426), .A2(new_n428), .B1(new_n442), .B2(G472), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n294), .A2(G119), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT23), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n378), .A2(G128), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n294), .A2(KEYINPUT23), .A3(G119), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G110), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n444), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT24), .B(G110), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n244), .B1(new_n198), .B2(KEYINPUT16), .ZN(new_n455));
  AND4_X1   g269(.A1(new_n244), .A2(new_n192), .A3(new_n193), .A4(KEYINPUT16), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(G146), .B1(new_n457), .B2(new_n241), .ZN(new_n458));
  INV_X1    g272(.A(new_n248), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT73), .B(G110), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n461), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n451), .A2(new_n452), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n199), .B2(new_n198), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n248), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n345), .A2(KEYINPUT22), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT22), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G137), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT74), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT74), .B1(new_n466), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT75), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT74), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n467), .A2(G137), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n345), .A2(KEYINPUT22), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT74), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n471), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n473), .B1(new_n471), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n460), .A2(new_n465), .A3(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT75), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n472), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n471), .A2(new_n480), .A3(new_n473), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n453), .B1(new_n247), .B2(new_n248), .ZN(new_n490));
  INV_X1    g304(.A(new_n465), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n492), .A3(new_n285), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT25), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n484), .A2(new_n492), .A3(KEYINPUT25), .A4(new_n285), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n323), .B1(new_n285), .B2(G234), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n484), .A2(new_n492), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(KEYINPUT76), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(KEYINPUT76), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n498), .A2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n443), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G221), .B1(new_n322), .B2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT77), .ZN(new_n509));
  INV_X1    g323(.A(G469), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(new_n275), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT81), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n362), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n372), .A2(KEYINPUT81), .A3(new_n361), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n360), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT3), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n230), .B2(G107), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n287), .A2(KEYINPUT3), .A3(G104), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n517), .A2(new_n518), .B1(new_n230), .B2(G107), .ZN(new_n519));
  AND2_X1   g333(.A1(KEYINPUT78), .A2(G101), .ZN(new_n520));
  NOR2_X1   g334(.A1(KEYINPUT78), .A2(G101), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT80), .B1(new_n287), .B2(G104), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT80), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n230), .A3(G107), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n287), .A2(G104), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n519), .A2(new_n522), .B1(new_n527), .B2(G101), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n515), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT10), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n367), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n518), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n230), .A2(G107), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n522), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G101), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n535), .B(KEYINPUT4), .C1(new_n536), .C2(new_n519), .ZN(new_n537));
  INV_X1    g351(.A(new_n519), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(G101), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n374), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n530), .B1(new_n360), .B2(new_n362), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n528), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n531), .A2(new_n532), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n363), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n527), .A2(G101), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n535), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n529), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT12), .B1(new_n549), .B2(new_n367), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n551), .B(new_n532), .C1(new_n548), .C2(new_n529), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n544), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(G110), .B(G140), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n212), .A2(G227), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n544), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n529), .A2(new_n530), .B1(new_n528), .B2(new_n542), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n532), .B1(new_n559), .B2(new_n541), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n553), .A2(new_n556), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n511), .B1(new_n562), .B2(G469), .ZN(new_n563));
  INV_X1    g377(.A(new_n544), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n556), .B1(new_n564), .B2(new_n560), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n544), .B(new_n557), .C1(new_n550), .C2(new_n552), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n510), .A3(new_n285), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n509), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G122), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT82), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n393), .A2(new_n537), .A3(new_n574), .A4(new_n540), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT5), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n378), .A3(G116), .ZN(new_n577));
  OAI211_X1 g391(.A(G113), .B(new_n577), .C1(new_n383), .C2(new_n576), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n392), .A3(new_n528), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n519), .A2(new_n536), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n391), .A2(new_n392), .B1(new_n581), .B2(new_n539), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n574), .B1(new_n582), .B2(new_n537), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n573), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n393), .A2(new_n537), .A3(new_n540), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT82), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n586), .A2(new_n572), .A3(new_n579), .A4(new_n575), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(KEYINPUT6), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT6), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n589), .B(new_n573), .C1(new_n580), .C2(new_n583), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n545), .A2(new_n187), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n371), .A2(G125), .A3(new_n373), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT83), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n371), .A2(KEYINPUT83), .A3(G125), .A4(new_n373), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G224), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G953), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n588), .A2(new_n590), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n572), .B(KEYINPUT8), .Z(new_n601));
  NAND2_X1  g415(.A1(new_n578), .A2(new_n392), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n547), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n603), .B2(new_n579), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT84), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n594), .A2(new_n605), .A3(new_n595), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT7), .B1(new_n597), .B2(G953), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n596), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n594), .A2(new_n595), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(KEYINPUT84), .A3(new_n591), .A4(new_n607), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n604), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n612), .B2(new_n587), .ZN(new_n613));
  OAI21_X1  g427(.A(G210), .B1(G237), .B2(G902), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT85), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n600), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n600), .B2(new_n613), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n571), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n570), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n342), .A2(new_n507), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(new_n522), .Z(G3));
  NAND2_X1  g436(.A1(new_n274), .A2(new_n282), .ZN(new_n623));
  INV_X1    g437(.A(new_n327), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n324), .B1(new_n306), .B2(new_n320), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(KEYINPUT98), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n627), .A2(KEYINPUT98), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n626), .B1(new_n630), .B2(new_n628), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n286), .A2(new_n283), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n283), .B1(new_n626), .B2(new_n286), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT99), .B1(new_n623), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  INV_X1    g451(.A(new_n635), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n637), .B(new_n638), .C1(new_n274), .C2(new_n282), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n339), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n641), .B(new_n571), .C1(new_n617), .C2(new_n618), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n399), .A2(new_n421), .A3(new_n408), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n411), .A2(new_n412), .B1(new_n417), .B2(new_n393), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n437), .B1(new_n645), .B2(new_n414), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n421), .B1(new_n399), .B2(new_n408), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n648), .B2(new_n286), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n649), .A2(new_n425), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n570), .A2(new_n506), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n640), .A2(new_n643), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n652), .B(new_n654), .ZN(G6));
  AND3_X1   g469(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n334), .B(new_n282), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n643), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(KEYINPUT101), .B1(new_n642), .B2(new_n658), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n650), .A3(new_n651), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n287), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT102), .B(KEYINPUT35), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n460), .A2(new_n483), .A3(new_n668), .A4(new_n465), .ZN(new_n669));
  OAI22_X1  g483(.A1(new_n490), .A2(new_n491), .B1(new_n489), .B2(KEYINPUT36), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n504), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n499), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n649), .A2(new_n425), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n342), .A2(new_n620), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(new_n673), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n426), .A2(new_n428), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n442), .A2(G472), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n336), .B1(new_n337), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n658), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n620), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n683), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n569), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n678), .A2(new_n334), .A3(new_n571), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n600), .A2(new_n613), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n615), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n600), .A2(new_n613), .A3(new_n616), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n275), .B1(new_n435), .B2(new_n437), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n404), .B1(new_n399), .B2(new_n411), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n679), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n697), .A2(new_n623), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n692), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT104), .B(G143), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G45));
  AOI21_X1  g519(.A(new_n638), .B1(new_n274), .B2(new_n282), .ZN(new_n706));
  INV_X1    g520(.A(new_n683), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n706), .A2(new_n620), .A3(new_n681), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  INV_X1    g523(.A(new_n428), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n427), .B1(new_n423), .B2(new_n424), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT29), .B1(new_n439), .B2(new_n440), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n437), .A2(KEYINPUT29), .ZN(new_n713));
  AOI211_X1 g527(.A(new_n713), .B(new_n429), .C1(new_n435), .C2(KEYINPUT28), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n712), .A2(new_n714), .A3(new_n286), .ZN(new_n715));
  INV_X1    g529(.A(G472), .ZN(new_n716));
  OAI22_X1  g530(.A1(new_n710), .A2(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n506), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n510), .B1(new_n567), .B2(new_n285), .ZN(new_n719));
  AOI211_X1 g533(.A(G469), .B(new_n286), .C1(new_n565), .C2(new_n566), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n509), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n643), .B(new_n723), .C1(new_n636), .C2(new_n639), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  AOI211_X1 g540(.A(KEYINPUT105), .B(new_n722), .C1(new_n661), .C2(new_n662), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n663), .B2(new_n723), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n308), .ZN(G18));
  INV_X1    g545(.A(new_n721), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n619), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n342), .A2(new_n681), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  OAI211_X1 g551(.A(new_n410), .B(new_n422), .C1(new_n436), .C2(new_n437), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n424), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n649), .A2(new_n739), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n732), .A2(new_n740), .A3(new_n506), .A4(new_n339), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n334), .B(new_n571), .C1(new_n617), .C2(new_n618), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n623), .A2(KEYINPUT107), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT107), .B1(new_n623), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT108), .B(G122), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G24));
  NAND3_X1  g562(.A1(new_n649), .A2(new_n673), .A3(new_n739), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n649), .A2(new_n673), .A3(new_n739), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n706), .A3(new_n707), .A4(new_n733), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n706), .A2(new_n707), .ZN(new_n757));
  INV_X1    g571(.A(new_n571), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n617), .A2(new_n618), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n717), .A2(new_n718), .A3(new_n569), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n756), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n638), .B(new_n683), .C1(new_n274), .C2(new_n282), .ZN(new_n762));
  INV_X1    g576(.A(new_n759), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n570), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(KEYINPUT42), .A3(new_n764), .A4(new_n507), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n507), .A3(new_n684), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  NOR2_X1   g583(.A1(new_n623), .A2(new_n638), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT43), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n650), .A2(new_n678), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(KEYINPUT44), .A3(new_n772), .ZN(new_n776));
  INV_X1    g590(.A(new_n509), .ZN(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n562), .B2(KEYINPUT45), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n562), .A2(KEYINPUT45), .ZN(new_n779));
  OAI22_X1  g593(.A1(new_n778), .A2(new_n779), .B1(new_n510), .B2(new_n275), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n780), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n568), .B1(new_n784), .B2(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n777), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n687), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n775), .A2(new_n759), .A3(new_n776), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  OAI21_X1  g604(.A(new_n786), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n791));
  XOR2_X1   g605(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n777), .B(new_n793), .C1(new_n783), .C2(new_n785), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n443), .A2(new_n506), .A3(new_n759), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n757), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  AND2_X1   g614(.A1(new_n771), .A2(new_n336), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n763), .A2(new_n732), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n507), .ZN(new_n804));
  NOR2_X1   g618(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n807));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n507), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n740), .A2(new_n506), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n733), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n212), .A2(G952), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n718), .A2(new_n679), .A3(new_n336), .A4(new_n700), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n802), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n812), .B1(new_n640), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n806), .A2(new_n808), .A3(new_n811), .A4(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n815), .A2(new_n623), .A3(new_n635), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n803), .B2(new_n753), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n801), .A2(new_n809), .A3(new_n759), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n791), .A2(new_n794), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n719), .A2(new_n720), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n777), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n821), .A2(new_n822), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n697), .A2(new_n571), .A3(new_n732), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT50), .B1(new_n810), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n810), .A2(KEYINPUT50), .A3(new_n830), .ZN(new_n832));
  OAI221_X1 g646(.A(new_n820), .B1(new_n828), .B2(new_n829), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n818), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  AND4_X1   g650(.A1(KEYINPUT106), .A2(new_n342), .A3(new_n681), .A4(new_n733), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n721), .A2(new_n696), .A3(new_n571), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n341), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT106), .B1(new_n839), .B2(new_n681), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n724), .B(new_n746), .C1(new_n837), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n836), .B1(new_n730), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n663), .A2(new_n723), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT105), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n663), .A2(new_n728), .A3(new_n723), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n724), .A2(new_n746), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n736), .A4(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n271), .A2(new_n268), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n334), .A2(new_n683), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n681), .A2(new_n282), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n753), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(new_n757), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n764), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n855), .A2(new_n766), .A3(new_n768), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n342), .B(new_n620), .C1(new_n507), .C2(new_n674), .ZN(new_n857));
  INV_X1    g671(.A(new_n623), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n706), .B1(new_n858), .B2(new_n334), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n651), .A2(new_n643), .A3(new_n650), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n857), .B(KEYINPUT112), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n754), .A2(new_n685), .A3(new_n708), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n701), .A2(new_n569), .A3(new_n678), .A4(new_n707), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n623), .A2(new_n743), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT107), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n623), .A2(new_n743), .A3(KEYINPUT107), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n868), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n570), .A2(new_n673), .A3(new_n683), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n701), .B(new_n877), .C1(new_n744), .C2(new_n745), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n620), .B(new_n681), .C1(new_n762), .C2(new_n684), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT52), .A4(new_n754), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n867), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n849), .A2(new_n866), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n730), .A2(new_n841), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n876), .A2(new_n880), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n865), .A4(new_n856), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n867), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n882), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(KEYINPUT113), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT113), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n885), .A2(new_n890), .A3(new_n867), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n885), .A2(new_n867), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n888), .B1(new_n893), .B2(KEYINPUT54), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n835), .B(new_n894), .C1(new_n834), .C2(new_n833), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n826), .A2(KEYINPUT49), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n638), .A2(new_n758), .A3(new_n509), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n897), .A2(new_n718), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  OR4_X1    g714(.A1(new_n623), .A2(new_n900), .A3(new_n697), .A4(new_n701), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n212), .A2(G952), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n882), .A2(new_n886), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n285), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT56), .B1(new_n906), .B2(new_n615), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n588), .A2(new_n590), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n599), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n904), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(KEYINPUT117), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n907), .A2(KEYINPUT118), .A3(new_n912), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(G51));
  XNOR2_X1  g731(.A(new_n511), .B(KEYINPUT57), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n887), .B1(new_n882), .B2(new_n886), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n888), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n567), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n779), .A2(new_n778), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT119), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n906), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n903), .B1(new_n921), .B2(new_n924), .ZN(G54));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n882), .A2(new_n886), .ZN(new_n927));
  AND4_X1   g741(.A1(KEYINPUT58), .A2(new_n927), .A3(G475), .A4(new_n286), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n265), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n904), .B1(new_n928), .B2(new_n265), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n928), .A2(new_n265), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(KEYINPUT120), .A3(new_n904), .A4(new_n929), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(G60));
  NAND2_X1  g749(.A1(new_n629), .A2(new_n631), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n894), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n936), .A2(new_n938), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n927), .A2(KEYINPUT54), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n882), .A2(new_n886), .A3(new_n887), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n941), .B1(new_n946), .B2(new_n903), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n942), .B1(new_n888), .B2(new_n919), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(KEYINPUT121), .A3(new_n904), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n951), .B(new_n936), .C1(new_n894), .C2(new_n938), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n940), .A2(new_n950), .A3(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n905), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n669), .A3(new_n670), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n503), .B1(new_n905), .B2(new_n955), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n904), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G66));
  OAI21_X1  g775(.A(G953), .B1(new_n338), .B2(new_n597), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT123), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n883), .A2(new_n865), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n212), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n908), .B1(G898), .B2(new_n212), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n965), .B(new_n966), .Z(G69));
  AOI21_X1  g781(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n788), .B(new_n507), .C1(new_n745), .C2(new_n744), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT125), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n754), .A2(new_n766), .A3(new_n768), .A4(new_n879), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n970), .A2(new_n799), .A3(new_n789), .A4(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n376), .B1(new_n398), .B2(KEYINPUT30), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT124), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(new_n259), .Z(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n212), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n869), .A2(new_n703), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT62), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n859), .A2(new_n787), .A3(new_n760), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n799), .A2(new_n978), .A3(new_n789), .A4(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n212), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n982), .B2(new_n975), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n968), .B1(new_n983), .B2(new_n682), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n968), .B2(new_n983), .ZN(G72));
  INV_X1    g799(.A(new_n893), .ZN(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  NAND2_X1  g802(.A1(new_n440), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n986), .A2(new_n699), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n978), .A2(new_n980), .ZN(new_n993));
  INV_X1    g807(.A(new_n964), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n993), .A2(new_n789), .A3(new_n799), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n992), .B1(new_n995), .B2(new_n988), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n992), .B(new_n988), .C1(new_n981), .C2(new_n964), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n699), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n988), .B1(new_n972), .B2(new_n964), .ZN(new_n1000));
  INV_X1    g814(.A(new_n440), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n903), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n991), .A2(new_n999), .A3(KEYINPUT127), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1002), .B1(new_n998), .B2(new_n996), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(new_n990), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1003), .A2(new_n1006), .ZN(G57));
endmodule


