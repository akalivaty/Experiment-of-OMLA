//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n191), .B1(G119), .B2(new_n190), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT23), .B1(new_n190), .B2(G119), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G119), .B(G128), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT24), .B(G110), .Z(new_n196));
  AOI22_X1  g010(.A1(new_n194), .A2(G110), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G125), .B(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n200), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(G146), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(G146), .B1(new_n199), .B2(new_n201), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n197), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI22_X1  g019(.A1(new_n194), .A2(G110), .B1(new_n195), .B2(new_n196), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT64), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT64), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n198), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n202), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT22), .B(G137), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT74), .ZN(new_n214));
  OR2_X1    g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n214), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n215), .B2(new_n218), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n205), .A2(new_n211), .A3(new_n221), .ZN(new_n224));
  AOI21_X1  g038(.A(G902), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n189), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI211_X1 g041(.A(KEYINPUT25), .B(G902), .C1(new_n223), .C2(new_n224), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT75), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n224), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n188), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT75), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n225), .A2(new_n226), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .A4(new_n189), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n189), .A2(G902), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT76), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n229), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT73), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n242));
  NOR2_X1   g056(.A1(G472), .A2(G902), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT64), .A2(G146), .ZN(new_n251));
  AOI21_X1  g065(.A(G143), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n247), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(G137), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT66), .B(G131), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n265), .A2(new_n259), .A3(new_n260), .A4(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n268), .B(new_n247), .C1(new_n252), .C2(new_n254), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n250), .A2(G143), .A3(new_n251), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G146), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n245), .A3(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n256), .A2(new_n267), .A3(new_n269), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n275));
  AND4_X1   g089(.A1(new_n275), .A2(new_n270), .A3(G128), .A4(new_n272), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n207), .A2(new_n208), .A3(new_n271), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT67), .B1(new_n277), .B2(new_n275), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n270), .A2(new_n279), .A3(KEYINPUT1), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(G128), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n252), .A2(new_n254), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n276), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n266), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n261), .A2(G134), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n260), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n274), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n190), .B1(new_n294), .B2(KEYINPUT67), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n282), .B1(new_n295), .B2(new_n280), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n289), .B1(new_n296), .B2(new_n276), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n270), .A2(new_n272), .ZN(new_n299));
  AOI22_X1  g113(.A1(KEYINPUT65), .A2(new_n255), .B1(new_n299), .B2(new_n245), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n267), .A4(new_n269), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n297), .A2(new_n298), .A3(KEYINPUT30), .A4(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G116), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G116), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n307), .A3(G119), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT68), .B(G116), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT69), .A3(G119), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n304), .A2(G119), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT2), .B(G113), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n313), .B1(new_n308), .B2(new_n309), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n316), .A3(new_n312), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n293), .A2(new_n303), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G210), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n323), .A2(G237), .A3(G953), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT27), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT26), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n297), .A2(new_n298), .A3(new_n302), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n319), .A2(new_n316), .A3(new_n312), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n316), .B1(new_n319), .B2(new_n312), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT71), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n318), .A2(new_n333), .A3(new_n320), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n328), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n322), .A2(KEYINPUT31), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT31), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n326), .B(G101), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n297), .A2(new_n298), .A3(new_n302), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT71), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n333), .B1(new_n318), .B2(new_n320), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n293), .A2(new_n303), .A3(new_n321), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n343), .A2(new_n297), .A3(new_n298), .A4(new_n302), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n291), .A2(new_n321), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n348), .B1(new_n291), .B2(new_n335), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n339), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n244), .B1(new_n347), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n242), .B1(new_n355), .B2(KEYINPUT32), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT31), .B1(new_n322), .B2(new_n336), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n338), .A3(new_n345), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT32), .B1(new_n359), .B2(new_n243), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n329), .A2(new_n335), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n322), .A2(new_n363), .A3(new_n328), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n328), .B1(new_n351), .B2(new_n353), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n329), .A2(new_n335), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n349), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n353), .B1(new_n369), .B2(KEYINPUT28), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n339), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(G902), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G472), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n357), .A2(new_n358), .ZN(new_n376));
  INV_X1    g190(.A(new_n350), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT28), .B1(new_n363), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n328), .B1(new_n378), .B2(new_n352), .ZN(new_n379));
  OAI211_X1 g193(.A(KEYINPUT32), .B(new_n243), .C1(new_n376), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n241), .B1(new_n362), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n359), .A2(new_n243), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT32), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT72), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI211_X1 g199(.A(new_n242), .B(KEYINPUT32), .C1(new_n359), .C2(new_n243), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G472), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n339), .B1(new_n378), .B2(new_n352), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n371), .B1(new_n389), .B2(new_n364), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n390), .B2(new_n373), .ZN(new_n391));
  INV_X1    g205(.A(new_n380), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(KEYINPUT73), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n240), .B1(new_n382), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G469), .ZN(new_n396));
  INV_X1    g210(.A(new_n284), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(G104), .ZN(new_n400));
  OR2_X1    g214(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n403));
  NOR2_X1   g217(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n404));
  OAI211_X1 g218(.A(G104), .B(new_n398), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n327), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT80), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n402), .A2(KEYINPUT80), .A3(new_n405), .A4(new_n327), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G104), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G107), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n327), .B1(new_n400), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT81), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n410), .A2(KEYINPUT84), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT84), .B1(new_n410), .B2(new_n414), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT10), .B(new_n397), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n190), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n299), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n270), .B2(new_n272), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT82), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n299), .A2(new_n275), .A3(G128), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n410), .A3(new_n414), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n426));
  NAND2_X1  g240(.A1(new_n402), .A2(new_n405), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(G101), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n269), .A2(new_n429), .A3(new_n256), .A4(new_n273), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n428), .B1(new_n427), .B2(G101), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n410), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n425), .A2(new_n426), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n267), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n417), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(G110), .B(G140), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n216), .A2(G227), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT12), .ZN(new_n441));
  INV_X1    g255(.A(new_n425), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n415), .A2(new_n416), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n284), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(new_n434), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n415), .A2(new_n416), .A3(new_n397), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT12), .B(new_n267), .C1(new_n446), .C2(new_n442), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n440), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n417), .A2(new_n433), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n267), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n439), .B1(new_n450), .B2(new_n435), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n396), .B(new_n188), .C1(new_n448), .C2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n396), .A2(new_n188), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n440), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n450), .ZN(new_n456));
  INV_X1    g270(.A(new_n435), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n445), .B2(new_n447), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n458), .B2(new_n439), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n452), .B(new_n454), .C1(new_n459), .C2(new_n396), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT9), .B(G234), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT77), .ZN(new_n462));
  OAI21_X1  g276(.A(G221), .B1(new_n462), .B2(G902), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n463), .B(KEYINPUT78), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G214), .B1(G237), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n313), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(G113), .B(new_n470), .C1(new_n315), .C2(new_n469), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n320), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n415), .B2(new_n416), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n432), .A2(new_n475), .A3(new_n321), .A4(new_n429), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n410), .A2(new_n431), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n429), .B1(new_n330), .B2(new_n331), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G122), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n474), .A2(new_n479), .A3(new_n481), .A4(new_n476), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n300), .A2(new_n269), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G125), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n284), .A2(new_n200), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n216), .A2(G224), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n489), .B(new_n490), .Z(new_n491));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n492), .A3(new_n482), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n487), .A2(new_n488), .B1(new_n495), .B2(new_n490), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n490), .A2(KEYINPUT7), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n410), .A2(new_n414), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n472), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT86), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n472), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n474), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n481), .B(KEYINPUT8), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n498), .A2(new_n484), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n188), .ZN(new_n508));
  OAI21_X1  g322(.A(G210), .B1(G237), .B2(G902), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n494), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n506), .A2(new_n484), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n512), .B2(new_n498), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n468), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n203), .A2(new_n204), .ZN(new_n518));
  NOR2_X1   g332(.A1(G237), .A2(G953), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(G143), .A3(G214), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(G143), .B1(new_n519), .B2(G214), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT88), .B1(new_n523), .B2(new_n265), .ZN(new_n524));
  INV_X1    g338(.A(new_n522), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n520), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT88), .ZN(new_n527));
  INV_X1    g341(.A(new_n265), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT90), .B(new_n518), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT90), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n524), .B2(new_n529), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n203), .A2(new_n204), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n523), .A2(new_n265), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n530), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(G113), .B(G122), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(new_n411), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n523), .B1(new_n542), .B2(new_n286), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n526), .A2(KEYINPUT18), .A3(G131), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n210), .B1(new_n249), .B2(new_n198), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n524), .A2(new_n537), .A3(new_n529), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT19), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n198), .B1(KEYINPUT89), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(KEYINPUT89), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n209), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n548), .B(new_n202), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n546), .ZN(new_n555));
  INV_X1    g369(.A(new_n541), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n547), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(G475), .A2(G902), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n517), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT20), .B(new_n561), .C1(new_n547), .C2(new_n557), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n539), .A2(new_n546), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n556), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n564), .B2(new_n547), .ZN(new_n565));
  INV_X1    g379(.A(G475), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n560), .A2(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G128), .B(G143), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n258), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n311), .A2(G122), .ZN(new_n570));
  AND2_X1   g384(.A1(KEYINPUT91), .A2(G122), .ZN(new_n571));
  NOR2_X1   g385(.A1(KEYINPUT91), .A2(G122), .ZN(new_n572));
  OAI21_X1  g386(.A(G116), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n573), .A3(new_n398), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT92), .ZN(new_n576));
  OR3_X1    g390(.A1(new_n570), .A2(new_n576), .A3(KEYINPUT14), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n570), .B2(KEYINPUT14), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n570), .A2(KEYINPUT14), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n573), .A4(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n580), .B2(G107), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n570), .A2(new_n573), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G107), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n584), .A2(new_n574), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n568), .A2(new_n258), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n568), .A2(KEYINPUT13), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n271), .A2(G128), .ZN(new_n588));
  OAI21_X1  g402(.A(G134), .B1(new_n588), .B2(KEYINPUT13), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n586), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n462), .A2(new_n187), .A3(G953), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n582), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n595));
  INV_X1    g409(.A(new_n593), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n581), .B2(new_n591), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(KEYINPUT93), .B(new_n596), .C1(new_n581), .C2(new_n591), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n188), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G478), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n602), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n598), .A2(new_n599), .A3(new_n188), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n216), .A2(G952), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(G234), .B2(G237), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n188), .B(new_n216), .C1(G234), .C2(G237), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT21), .B(G898), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OR3_X1    g425(.A1(new_n567), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n516), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n395), .A2(new_n467), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  OR2_X1    g429(.A1(new_n516), .A2(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n600), .A2(new_n601), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n598), .A2(new_n618), .A3(new_n599), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n594), .A2(KEYINPUT33), .A3(new_n597), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n188), .A2(G478), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n617), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n567), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n388), .B1(new_n359), .B2(new_n188), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n627), .A2(new_n355), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n466), .A2(new_n240), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT94), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G6));
  INV_X1    g447(.A(KEYINPUT95), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n562), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n558), .A2(new_n517), .A3(new_n559), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT95), .ZN(new_n637));
  INV_X1    g451(.A(new_n560), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n565), .A2(new_n566), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n606), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n616), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n629), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n221), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n212), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n237), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n229), .A2(new_n235), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT96), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n628), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n613), .A2(new_n467), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT97), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n608), .B1(new_n609), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n639), .A2(new_n640), .A3(new_n606), .A4(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n656), .B1(new_n516), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n641), .ZN(new_n662));
  INV_X1    g476(.A(new_n468), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n510), .B1(new_n494), .B2(new_n508), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n513), .A2(new_n514), .A3(new_n509), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n662), .A2(new_n666), .A3(KEYINPUT98), .A4(new_n659), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n382), .A2(new_n394), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n649), .B(KEYINPUT96), .Z(new_n670));
  NAND4_X1  g484(.A1(new_n668), .A2(new_n669), .A3(new_n467), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XOR2_X1   g486(.A(new_n658), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n467), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n188), .B1(new_n369), .B2(new_n328), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n339), .B1(new_n345), .B2(new_n349), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n380), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n356), .A2(new_n679), .A3(new_n361), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n356), .A2(new_n679), .A3(KEYINPUT99), .A4(new_n361), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n664), .A2(new_n665), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(KEYINPUT38), .Z(new_n687));
  AND3_X1   g501(.A1(new_n567), .A2(new_n606), .A3(new_n468), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n650), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT100), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n675), .A2(new_n685), .A3(new_n687), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n271), .ZN(G45));
  NAND3_X1  g506(.A1(new_n624), .A2(new_n567), .A3(new_n659), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n516), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n669), .A2(new_n467), .A3(new_n670), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  OAI21_X1  g510(.A(new_n188), .B1(new_n448), .B2(new_n451), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(G469), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n452), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n464), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n395), .A2(new_n626), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND3_X1  g517(.A1(new_n395), .A2(new_n642), .A3(new_n700), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT101), .B(G116), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G18));
  NOR4_X1   g520(.A1(new_n516), .A2(new_n612), .A3(new_n699), .A4(new_n464), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n669), .A2(new_n670), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  NAND2_X1  g523(.A1(new_n686), .A2(new_n688), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n699), .A2(new_n464), .A3(new_n611), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n357), .B(new_n358), .C1(new_n370), .C2(new_n328), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(KEYINPUT102), .A3(new_n243), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT102), .B1(new_n713), .B2(new_n243), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n714), .A2(new_n715), .A3(new_n627), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n711), .A2(new_n712), .A3(new_n239), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AND2_X1   g532(.A1(new_n670), .A2(new_n716), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n516), .A2(new_n464), .A3(new_n699), .ZN(new_n720));
  INV_X1    g534(.A(new_n693), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n664), .A2(new_n665), .A3(new_n468), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n466), .A2(new_n693), .A3(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n362), .A2(new_n381), .A3(new_n241), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT73), .B1(new_n387), .B2(new_n393), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n239), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT103), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n395), .A2(new_n733), .A3(new_n728), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n726), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n360), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT105), .A3(new_n380), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n392), .B2(new_n360), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n739), .A3(new_n375), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n239), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT106), .A3(KEYINPUT42), .A4(new_n728), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  INV_X1    g558(.A(new_n727), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n467), .A2(new_n745), .A3(new_n721), .A4(KEYINPUT42), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n746), .B2(new_n741), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n724), .B1(new_n735), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n731), .A2(KEYINPUT103), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n733), .B1(new_n395), .B2(new_n728), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n725), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n743), .A2(new_n747), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(KEYINPUT107), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  NOR3_X1   g570(.A1(new_n466), .A2(new_n660), .A3(new_n727), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n239), .B(new_n757), .C1(new_n729), .C2(new_n730), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n395), .A2(new_n760), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n459), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n396), .B1(new_n459), .B2(new_n764), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n453), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n452), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n464), .ZN(new_n772));
  INV_X1    g586(.A(new_n567), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n624), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT43), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT43), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n624), .A2(new_n776), .A3(new_n773), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n670), .A2(new_n628), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(new_n778), .B2(new_n779), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n745), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n772), .A2(new_n673), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  OR3_X1    g599(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n464), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT47), .B1(new_n771), .B2(new_n464), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n669), .A2(new_n239), .A3(new_n693), .A4(new_n727), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n791));
  NOR2_X1   g605(.A1(G952), .A2(G953), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n606), .A2(new_n658), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n639), .A2(new_n793), .A3(new_n640), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n466), .A2(new_n727), .A3(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n670), .B(new_n795), .C1(new_n729), .C2(new_n730), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n669), .A2(KEYINPUT111), .A3(new_n670), .A4(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n719), .A2(new_n467), .A3(new_n721), .A4(new_n745), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n762), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n395), .B(new_n700), .C1(new_n626), .C2(new_n642), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n516), .A2(new_n611), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n773), .A2(new_n606), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n625), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n629), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n807), .A2(new_n652), .A3(new_n717), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n803), .A2(new_n808), .A3(new_n614), .A4(new_n708), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n802), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n671), .A2(new_n695), .A3(new_n722), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n649), .A2(new_n658), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n460), .A2(new_n465), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n710), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n684), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n813), .B1(new_n684), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n811), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n466), .B(new_n650), .C1(new_n382), .C2(new_n394), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n668), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT99), .B1(new_n387), .B2(new_n679), .ZN(new_n824));
  AND4_X1   g638(.A1(KEYINPUT99), .A2(new_n356), .A3(new_n679), .A4(new_n361), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n816), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT112), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n684), .A2(new_n813), .A3(new_n816), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n823), .A2(KEYINPUT52), .A3(new_n695), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n820), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n810), .A2(new_n831), .A3(new_n749), .A4(new_n754), .ZN(new_n832));
  XOR2_X1   g646(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n752), .B2(new_n753), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n838), .B(new_n839), .C1(new_n812), .C2(new_n819), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n829), .A2(new_n671), .A3(new_n695), .A4(new_n722), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n839), .B1(new_n842), .B2(new_n838), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n810), .B(new_n837), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n834), .A2(new_n835), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n841), .A2(new_n843), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n762), .A2(new_n800), .A3(new_n801), .ZN(new_n847));
  INV_X1    g661(.A(new_n809), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n749), .A2(new_n754), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n836), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n833), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n755), .A2(new_n810), .A3(new_n851), .A4(new_n831), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n835), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n727), .A2(new_n699), .A3(new_n464), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n608), .A2(new_n855), .A3(new_n775), .A4(new_n777), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n742), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT48), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n607), .B(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n716), .A2(new_n239), .ZN(new_n860));
  INV_X1    g674(.A(new_n608), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n778), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n862), .B2(new_n720), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n685), .A2(new_n239), .A3(new_n608), .A4(new_n855), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n858), .B(new_n863), .C1(new_n625), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n700), .A2(new_n663), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n862), .A3(new_n687), .A4(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n856), .A2(new_n719), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n864), .A2(new_n567), .A3(new_n624), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n699), .A2(new_n465), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n786), .B2(new_n787), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n745), .B(new_n862), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT51), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n862), .A2(new_n745), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n875), .B(new_n883), .C1(new_n877), .C2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n865), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n792), .B1(new_n854), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n699), .A2(KEYINPUT49), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT109), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n239), .A2(new_n465), .A3(new_n468), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n890), .B(new_n774), .C1(KEYINPUT49), .C2(new_n699), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n685), .A2(new_n889), .A3(new_n687), .A4(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT110), .Z(new_n893));
  OAI21_X1  g707(.A(new_n791), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n850), .A2(new_n852), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT54), .ZN(new_n896));
  INV_X1    g710(.A(new_n846), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n810), .A2(new_n837), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n897), .A2(new_n898), .B1(new_n832), .B2(new_n833), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n835), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n886), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n792), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n893), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(KEYINPUT120), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n894), .A2(new_n905), .ZN(G75));
  NAND2_X1  g720(.A1(new_n485), .A2(new_n493), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(new_n491), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n899), .A2(new_n323), .A3(new_n188), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n910), .B2(KEYINPUT56), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n216), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n910), .A2(KEYINPUT56), .A3(new_n909), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(G51));
  NOR2_X1   g730(.A1(new_n899), .A2(new_n835), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n845), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n453), .B(KEYINPUT57), .Z(new_n919));
  OAI22_X1  g733(.A1(new_n918), .A2(new_n919), .B1(new_n451), .B2(new_n448), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n899), .A2(new_n188), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n766), .A3(new_n767), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n912), .B1(new_n920), .B2(new_n922), .ZN(G54));
  AND2_X1   g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n921), .A2(new_n558), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n558), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n912), .ZN(G60));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  OR2_X1    g743(.A1(new_n622), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n913), .B1(new_n918), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n854), .A2(new_n929), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n622), .B2(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n834), .B2(new_n844), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n912), .B1(new_n936), .B2(new_n647), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT122), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n230), .B(KEYINPUT121), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n899), .B2(new_n935), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n941), .A3(KEYINPUT61), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n937), .B(new_n940), .C1(KEYINPUT122), .C2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(G66));
  XNOR2_X1  g759(.A(new_n809), .B(KEYINPUT123), .ZN(new_n946));
  NAND2_X1  g760(.A1(G224), .A2(G953), .ZN(new_n947));
  OAI22_X1  g761(.A1(new_n946), .A2(G953), .B1(new_n610), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n907), .B1(G898), .B2(new_n216), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  OR2_X1    g766(.A1(new_n691), .A2(new_n812), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n955));
  AOI211_X1 g769(.A(new_n727), .B(new_n674), .C1(new_n625), .C2(new_n805), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n395), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n789), .A2(new_n784), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n216), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n293), .A2(new_n303), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(new_n552), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n772), .A2(new_n673), .A3(new_n711), .A4(new_n742), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n762), .A2(new_n789), .A3(new_n784), .A4(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n812), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n755), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n968), .B2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n216), .B1(G227), .B2(G900), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G72));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n968), .B2(new_n946), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n365), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n974), .B1(new_n959), .B2(new_n946), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n912), .B1(new_n979), .B2(new_n677), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n974), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n364), .A2(new_n677), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n895), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n984), .A2(KEYINPUT127), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(KEYINPUT127), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(G57));
endmodule


