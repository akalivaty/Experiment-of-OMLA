//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  AND2_X1   g0008(.A1(G107), .A2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n209), .B(new_n215), .C1(G97), .C2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT68), .B(G77), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(new_n204), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT67), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n208), .B(new_n223), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n212), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n214), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT70), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(new_n250), .A3(new_n229), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n249), .B2(new_n229), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G68), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n211), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G58), .A2(G68), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G159), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT66), .B(G20), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n224), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT78), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT78), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n264), .A2(KEYINPUT7), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n261), .B1(new_n275), .B2(G68), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n254), .B1(new_n276), .B2(KEYINPUT16), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n278), .A2(new_n279), .A3(G20), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT79), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n228), .A2(new_n283), .A3(KEYINPUT7), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT79), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n269), .A2(new_n285), .A3(new_n274), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n261), .B1(new_n287), .B2(G68), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n277), .B1(KEYINPUT16), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n291), .B1(G223), .B2(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G87), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n292), .A2(KEYINPUT80), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT80), .B1(new_n292), .B2(new_n293), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT69), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G1), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n296), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G232), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n299), .A3(G274), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(G200), .B1(new_n298), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n295), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n292), .A2(KEYINPUT80), .A3(new_n293), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n296), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n310), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(G190), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT69), .B(G1), .ZN(new_n317));
  INV_X1    g0117(.A(G13), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n317), .A2(new_n318), .A3(new_n224), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT8), .B(G58), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n249), .A2(new_n229), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n251), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n317), .A2(new_n224), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n322), .B1(new_n328), .B2(new_n321), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n289), .A2(new_n311), .A3(new_n316), .A4(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT17), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n287), .A2(G68), .ZN(new_n334));
  INV_X1    g0134(.A(new_n261), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT16), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT7), .B1(new_n228), .B2(new_n283), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n269), .A2(new_n274), .ZN(new_n338));
  OAI21_X1  g0138(.A(G68), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(KEYINPUT16), .A3(new_n335), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n325), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n330), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n343), .A2(KEYINPUT17), .A3(new_n311), .A4(new_n316), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n333), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G169), .B1(new_n298), .B2(new_n310), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n314), .A2(new_n315), .A3(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n342), .A2(new_n348), .A3(KEYINPUT18), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT18), .B1(new_n342), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT81), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n342), .A2(new_n348), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT81), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n342), .A2(new_n348), .A3(KEYINPUT18), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n345), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G1698), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G222), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G223), .A2(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n263), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n220), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n296), .C1(new_n363), .C2(new_n263), .ZN(new_n364));
  INV_X1    g0164(.A(new_n307), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n364), .B(new_n309), .C1(new_n365), .C2(new_n290), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G200), .ZN(new_n367));
  XOR2_X1   g0167(.A(new_n367), .B(KEYINPUT74), .Z(new_n368));
  INV_X1    g0168(.A(G50), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n257), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n228), .A2(G33), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n320), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n327), .A2(G50), .B1(new_n373), .B2(new_n325), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n303), .A2(G13), .A3(G20), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(G50), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT9), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n366), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n368), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT10), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT10), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n368), .A2(new_n377), .A3(new_n382), .A4(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G169), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n366), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT71), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n366), .A2(G179), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n372), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT73), .ZN(new_n394));
  INV_X1    g0194(.A(new_n259), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n228), .A2(new_n220), .B1(new_n320), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT72), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n325), .B1(new_n220), .B2(new_n319), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n327), .A2(G77), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G238), .A2(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n263), .B(new_n402), .C1(new_n212), .C2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n296), .C1(G107), .C2(new_n263), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(new_n309), .C1(new_n219), .C2(new_n365), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(G179), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n385), .B2(new_n405), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n358), .A2(new_n384), .A3(new_n391), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n263), .A2(G226), .A3(new_n359), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G97), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT76), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT76), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(G33), .A3(G97), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n263), .A2(G232), .A3(G1698), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n263), .A2(KEYINPUT75), .A3(G226), .A4(new_n359), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n412), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n296), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n307), .A2(G238), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n309), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n420), .A2(new_n296), .B1(G238), .B2(new_n307), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n309), .ZN(new_n427));
  OAI21_X1  g0227(.A(G200), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n319), .A2(new_n255), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT12), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n255), .A2(G20), .ZN(new_n431));
  INV_X1    g0231(.A(G77), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n431), .B1(new_n369), .B2(new_n395), .C1(new_n372), .C2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n433), .A2(new_n325), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n430), .B1(new_n255), .B2(new_n328), .C1(new_n434), .C2(KEYINPUT11), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(KEYINPUT11), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n426), .A2(new_n425), .A3(new_n309), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(G190), .A3(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n428), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n405), .A2(G200), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n405), .A2(new_n378), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n401), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n439), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT14), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n447), .A2(G169), .B1(KEYINPUT77), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(KEYINPUT77), .ZN(new_n450));
  AOI211_X1 g0250(.A(new_n385), .B(new_n450), .C1(new_n438), .C2(new_n439), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n438), .A2(G179), .A3(new_n439), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n448), .A2(KEYINPUT77), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n449), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n442), .B(new_n446), .C1(new_n456), .C2(new_n437), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n409), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n303), .A2(G33), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n254), .A2(new_n375), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n375), .A2(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT25), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT23), .A2(G107), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n225), .A2(new_n227), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT23), .A2(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(G20), .C2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT22), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n225), .A2(new_n227), .B1(new_n267), .B2(new_n268), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G87), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n228), .A2(new_n263), .A3(new_n473), .A4(G87), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n472), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n228), .A2(new_n263), .A3(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT22), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n476), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n479), .A3(new_n472), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n466), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n462), .B(new_n464), .C1(new_n486), .C2(new_n254), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n278), .A2(new_n279), .B1(G250), .B2(G1698), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n359), .A2(G257), .ZN(new_n489));
  INV_X1    g0289(.A(G294), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n488), .A2(new_n489), .B1(new_n266), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n296), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT5), .B(G41), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n303), .A2(new_n493), .A3(G45), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(G264), .A3(new_n297), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n305), .B1(new_n300), .B2(new_n302), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n297), .A2(new_n496), .A3(G274), .A4(new_n493), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G179), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n385), .B2(new_n498), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n480), .B(new_n471), .C1(new_n483), .C2(new_n476), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n479), .B1(new_n484), .B2(new_n472), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(KEYINPUT87), .B2(new_n465), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n325), .ZN(new_n505));
  INV_X1    g0305(.A(G200), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT88), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n492), .A2(new_n495), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n378), .A3(new_n497), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT88), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n498), .A2(new_n511), .A3(new_n506), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n505), .A2(new_n513), .A3(new_n462), .A4(new_n464), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n228), .A2(G33), .A3(G97), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n515), .A2(new_n516), .B1(new_n474), .B2(G68), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n414), .A2(new_n416), .A3(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n228), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n217), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n254), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n392), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n375), .A2(new_n524), .ZN(new_n525));
  AND4_X1   g0325(.A1(G87), .A2(new_n254), .A3(new_n375), .A4(new_n459), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n263), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n263), .A2(G238), .A3(new_n359), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n296), .ZN(new_n535));
  INV_X1    g0335(.A(G274), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n296), .B1(new_n496), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n218), .B1(new_n317), .B2(new_n305), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n534), .A2(new_n296), .B1(new_n538), .B2(new_n537), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n527), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n385), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n228), .A2(new_n263), .A3(G68), .ZN(new_n546));
  INV_X1    g0346(.A(G97), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n262), .A2(new_n266), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n548), .B2(KEYINPUT19), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n518), .A2(new_n228), .B1(new_n217), .B2(new_n520), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n325), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n525), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n254), .A2(new_n375), .A3(new_n524), .A4(new_n459), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(G179), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n542), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n545), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n544), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n501), .A2(new_n514), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n218), .B1(new_n267), .B2(new_n268), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT4), .ZN(new_n561));
  OAI21_X1  g0361(.A(G1698), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G283), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n266), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(G244), .B1(new_n278), .B2(new_n279), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(new_n561), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n359), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n296), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n494), .A2(G257), .A3(new_n297), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n497), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n378), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n319), .A2(new_n547), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n460), .A2(new_n547), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n259), .A2(G77), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT6), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n576), .A2(new_n547), .A3(G107), .ZN(new_n577));
  XNOR2_X1  g0377(.A(G97), .B(G107), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n575), .B1(new_n579), .B2(new_n228), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n287), .B2(G107), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n573), .B(new_n574), .C1(new_n581), .C2(new_n254), .ZN(new_n582));
  INV_X1    g0382(.A(new_n497), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n568), .B2(new_n296), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n506), .B1(new_n584), .B2(new_n570), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n572), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n571), .A2(new_n385), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n555), .A3(new_n570), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(KEYINPUT82), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT82), .ZN(new_n592));
  INV_X1    g0392(.A(new_n585), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n378), .B2(new_n571), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n591), .B(new_n592), .C1(new_n594), .C2(new_n582), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n254), .A2(G116), .A3(new_n375), .A4(new_n459), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n375), .A2(G116), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n547), .A2(G33), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n228), .B(new_n601), .C1(new_n266), .C2(new_n563), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n249), .A2(new_n229), .B1(G20), .B2(new_n213), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n597), .B(new_n599), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n359), .A2(G257), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G264), .A2(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n263), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G303), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n283), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n613), .A3(new_n296), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n494), .A2(G270), .A3(new_n297), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT84), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n615), .A2(new_n616), .A3(new_n497), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n615), .B2(new_n497), .ZN(new_n618));
  OAI211_X1 g0418(.A(G179), .B(new_n614), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT85), .B1(new_n608), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n614), .ZN(new_n621));
  INV_X1    g0421(.A(new_n618), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n615), .A2(new_n616), .A3(new_n497), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT85), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n624), .A2(new_n625), .A3(G179), .A4(new_n607), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT20), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n262), .A2(new_n564), .A3(new_n600), .ZN(new_n628));
  INV_X1    g0428(.A(new_n603), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n598), .B1(new_n630), .B2(new_n604), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n385), .B1(new_n631), .B2(new_n597), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT21), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n632), .B2(new_n634), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n620), .B(new_n626), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n634), .A2(G200), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT86), .B1(new_n638), .B2(new_n608), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT86), .ZN(new_n640));
  AOI211_X1 g0440(.A(new_n640), .B(new_n607), .C1(new_n634), .C2(G200), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n624), .A2(G190), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n637), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n458), .A2(new_n559), .A3(new_n596), .A4(new_n644), .ZN(G372));
  OAI21_X1  g0445(.A(new_n408), .B1(new_n456), .B2(new_n437), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n333), .A2(new_n344), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n442), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n354), .A2(new_n356), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n390), .B1(new_n650), .B2(new_n384), .ZN(new_n651));
  INV_X1    g0451(.A(new_n458), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n516), .A2(new_n515), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n522), .A2(new_n546), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n525), .B1(new_n654), .B2(new_n325), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n655), .A2(new_n553), .B1(new_n555), .B2(new_n542), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n535), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n534), .A2(KEYINPUT89), .A3(new_n296), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n658), .A2(new_n659), .B1(new_n538), .B2(new_n537), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n656), .B1(new_n660), .B2(G169), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n543), .B(new_n527), .C1(new_n660), .C2(new_n506), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n514), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n586), .A2(new_n589), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n635), .A2(new_n636), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n620), .A2(new_n626), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n501), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n664), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n589), .A2(new_n662), .A3(new_n661), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n544), .A2(new_n557), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n673), .B2(new_n591), .ZN(new_n674));
  AND4_X1   g0474(.A1(new_n670), .A2(new_n672), .A3(new_n674), .A4(new_n661), .ZN(new_n675));
  INV_X1    g0475(.A(new_n661), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n584), .A2(new_n555), .A3(new_n570), .ZN(new_n677));
  AOI21_X1  g0477(.A(G169), .B1(new_n584), .B2(new_n570), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(new_n544), .A3(new_n557), .A4(new_n582), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n680), .B2(KEYINPUT26), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n670), .B1(new_n681), .B2(new_n672), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n669), .B1(new_n675), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n651), .B1(new_n652), .B2(new_n684), .ZN(G369));
  NAND2_X1  g0485(.A1(new_n228), .A2(G13), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .A3(new_n317), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT27), .B1(new_n686), .B2(new_n317), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n644), .B1(new_n608), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n637), .A2(new_n607), .A3(new_n691), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n487), .A2(new_n691), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n698), .A2(new_n514), .B1(new_n487), .B2(new_n500), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n501), .A2(new_n691), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n691), .B1(new_n666), .B2(new_n667), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n700), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n205), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G41), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n521), .A2(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n231), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g0511(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n712));
  XNOR2_X1  g0512(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n665), .A2(KEYINPUT95), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT95), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n586), .B2(new_n589), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n664), .A3(new_n668), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n671), .B1(new_n673), .B2(new_n591), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n662), .A2(new_n661), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT26), .A3(new_n589), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n661), .B(KEYINPUT93), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n718), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n692), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n672), .A2(new_n674), .A3(new_n661), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n681), .A2(new_n670), .A3(new_n672), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n691), .B1(new_n733), .B2(new_n669), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n619), .A2(new_n540), .ZN(new_n738));
  INV_X1    g0538(.A(new_n571), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n509), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n738), .A2(KEYINPUT30), .A3(new_n509), .A4(new_n739), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n660), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(new_n555), .A3(new_n498), .A4(new_n634), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n739), .ZN(new_n747));
  OAI211_X1 g0547(.A(KEYINPUT31), .B(new_n691), .C1(new_n744), .C2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT92), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n742), .A2(new_n743), .ZN(new_n751));
  INV_X1    g0551(.A(new_n747), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n692), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n644), .A2(new_n596), .A3(new_n559), .A4(new_n692), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(KEYINPUT31), .ZN(new_n755));
  OAI21_X1  g0555(.A(G330), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n737), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n713), .B1(new_n757), .B2(G1), .ZN(G364));
  AOI21_X1  g0558(.A(new_n229), .B1(G20), .B2(new_n385), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n262), .A2(G179), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT98), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n263), .B1(new_n765), .B2(G326), .ZN(new_n766));
  NOR4_X1   g0566(.A1(new_n228), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G329), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n506), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n262), .A2(new_n378), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n768), .B1(new_n563), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT100), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(KEYINPUT100), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n766), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n763), .A2(new_n378), .A3(new_n506), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n774), .B1(G311), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n763), .A2(new_n378), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n506), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI21_X1  g0581(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n763), .A2(G190), .A3(new_n506), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n782), .B1(G322), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n378), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n228), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n769), .A2(G20), .A3(G190), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n785), .B1(new_n490), .B2(new_n787), .C1(new_n612), .C2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n783), .A2(new_n211), .B1(new_n547), .B2(new_n787), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n283), .B1(new_n791), .B2(G87), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n792), .B1(new_n461), .B2(new_n770), .C1(new_n764), .C2(new_n369), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n790), .B(new_n793), .C1(G68), .C2(new_n779), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n767), .A2(G159), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT32), .Z(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(new_n220), .C2(new_n775), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT99), .Z(new_n798));
  AOI21_X1  g0598(.A(new_n760), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n686), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n299), .B1(new_n800), .B2(G45), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n707), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n759), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n205), .A2(new_n263), .ZN(new_n810));
  INV_X1    g0610(.A(G355), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n811), .B1(G116), .B2(new_n205), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT97), .Z(new_n813));
  NOR2_X1   g0613(.A1(new_n706), .A2(new_n263), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n232), .A2(new_n305), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n305), .C2(new_n244), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n809), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n799), .A2(new_n804), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n807), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n695), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G330), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n693), .A2(new_n821), .A3(new_n694), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n696), .A2(new_n804), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT96), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(KEYINPUT96), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n820), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT101), .ZN(G396));
  INV_X1    g0627(.A(KEYINPUT104), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n692), .B1(new_n399), .B2(new_n400), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n408), .B1(new_n445), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n408), .A2(new_n691), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT103), .B1(new_n734), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n734), .B2(new_n834), .ZN(new_n836));
  OAI211_X1 g0636(.A(KEYINPUT103), .B(new_n833), .C1(new_n684), .C2(new_n691), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n748), .B(KEYINPUT92), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n754), .A2(KEYINPUT31), .ZN(new_n840));
  INV_X1    g0640(.A(new_n753), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n821), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n828), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n803), .B1(new_n838), .B2(new_n843), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n836), .A2(KEYINPUT104), .A3(new_n756), .A4(new_n837), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n780), .A2(new_n563), .B1(new_n490), .B2(new_n783), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(G116), .B2(new_n776), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n765), .A2(G303), .ZN(new_n850));
  INV_X1    g0650(.A(new_n767), .ZN(new_n851));
  INV_X1    g0651(.A(G311), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n851), .A2(new_n852), .B1(new_n217), .B2(new_n770), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT102), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n283), .B1(new_n788), .B2(new_n461), .ZN(new_n855));
  INV_X1    g0655(.A(new_n787), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(G97), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n849), .A2(new_n850), .A3(new_n854), .A4(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G150), .A2(new_n779), .B1(new_n784), .B2(G143), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  INV_X1    g0660(.A(G159), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n859), .B1(new_n860), .B2(new_n764), .C1(new_n861), .C2(new_n775), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT34), .Z(new_n863));
  INV_X1    g0663(.A(new_n770), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G58), .A2(new_n856), .B1(new_n864), .B2(G68), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n283), .B1(new_n791), .B2(G50), .ZN(new_n866));
  INV_X1    g0666(.A(G132), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n865), .B(new_n866), .C1(new_n867), .C2(new_n851), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n858), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n804), .B1(new_n869), .B2(new_n759), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n759), .A2(new_n805), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(G77), .B2(new_n872), .C1(new_n806), .C2(new_n834), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n847), .A2(new_n873), .ZN(G384));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  INV_X1    g0675(.A(new_n689), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n342), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n647), .B2(new_n649), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n342), .B1(new_n348), .B2(new_n876), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n331), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n880), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n875), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n276), .A2(KEYINPUT16), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n330), .B1(new_n884), .B2(new_n341), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n876), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n348), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n331), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n331), .A2(new_n879), .A3(new_n881), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(KEYINPUT38), .B(new_n891), .C1(new_n358), .C2(new_n886), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n456), .A2(new_n437), .A3(new_n691), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n351), .A2(new_n357), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n886), .B1(new_n897), .B2(new_n647), .ZN(new_n898));
  INV_X1    g0698(.A(new_n891), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n875), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n892), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n895), .B(new_n896), .C1(new_n894), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n354), .A2(new_n356), .A3(new_n689), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n437), .A2(new_n692), .ZN(new_n904));
  OAI21_X1  g0704(.A(G169), .B1(new_n424), .B2(new_n427), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n450), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n447), .A2(KEYINPUT77), .A3(new_n448), .A4(G169), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n454), .A4(new_n452), .ZN(new_n908));
  INV_X1    g0708(.A(new_n437), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n904), .B(new_n441), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n691), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n683), .A2(new_n692), .A3(new_n834), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(new_n832), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n901), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n902), .A2(new_n903), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n652), .B1(new_n729), .B2(new_n736), .ZN(new_n918));
  INV_X1    g0718(.A(new_n651), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n917), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n842), .A2(new_n748), .ZN(new_n922));
  INV_X1    g0722(.A(new_n904), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n442), .B(new_n923), .C1(new_n456), .C2(new_n437), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n833), .B1(new_n924), .B2(new_n911), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n901), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT40), .ZN(new_n927));
  INV_X1    g0727(.A(new_n748), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n925), .B1(new_n755), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n883), .B2(new_n892), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n926), .A2(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n458), .A3(new_n922), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n900), .A2(new_n892), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n927), .B1(new_n934), .B2(new_n929), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n922), .A3(new_n925), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(G330), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n458), .B(G330), .C1(new_n755), .C2(new_n928), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n933), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n921), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n303), .B2(new_n800), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n579), .B(KEYINPUT105), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n213), .B1(new_n944), .B2(KEYINPUT35), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n945), .B(new_n230), .C1(KEYINPUT35), .C2(new_n944), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n256), .A2(new_n231), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n948), .A2(new_n220), .B1(G50), .B2(new_n255), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n318), .A3(new_n317), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  INV_X1    g0751(.A(G317), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n283), .B1(new_n547), .B2(new_n770), .C1(new_n851), .C2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT110), .Z(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G311), .B2(new_n765), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n780), .A2(new_n490), .B1(new_n612), .B2(new_n783), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G283), .B2(new_n776), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n856), .A2(G107), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n791), .A2(G116), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT46), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n955), .A2(new_n957), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n775), .A2(new_n369), .ZN(new_n962));
  INV_X1    g0762(.A(G150), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n783), .A2(new_n963), .B1(new_n220), .B2(new_n770), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n962), .B(new_n964), .C1(G137), .C2(new_n767), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n779), .A2(G159), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n856), .A2(G68), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n283), .B1(new_n791), .B2(G58), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n765), .A2(G143), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n961), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT47), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n759), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n692), .A2(new_n527), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n722), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n661), .A2(new_n974), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n807), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n814), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n808), .B1(new_n205), .B2(new_n392), .C1(new_n240), .C2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n973), .A2(new_n803), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n582), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n717), .B1(new_n981), .B2(new_n692), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n701), .A2(new_n703), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n591), .B1(new_n982), .B2(new_n501), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n692), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n984), .A2(new_n986), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n975), .A2(new_n976), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT107), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n589), .A2(new_n691), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n982), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n998), .B1(new_n702), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n702), .A2(new_n1001), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n995), .A2(new_n1003), .A3(new_n997), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1002), .A2(new_n1006), .A3(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n701), .B(new_n703), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n697), .B1(KEYINPUT109), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(KEYINPUT109), .B2(new_n1011), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1013), .A2(new_n702), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1000), .A2(new_n704), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT45), .Z(new_n1016));
  OR3_X1    g0816(.A1(new_n1000), .A2(KEYINPUT44), .A3(new_n704), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT44), .B1(new_n1000), .B2(new_n704), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1014), .A2(new_n757), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n757), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n707), .B(KEYINPUT41), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n802), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n980), .B1(new_n1010), .B2(new_n1025), .ZN(G387));
  AOI22_X1  g0826(.A1(G311), .A2(new_n779), .B1(new_n784), .B2(G317), .ZN(new_n1027));
  INV_X1    g0827(.A(G322), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1027), .B1(new_n612), .B2(new_n775), .C1(new_n1028), .C2(new_n764), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n563), .B2(new_n787), .C1(new_n490), .C2(new_n788), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n864), .A2(G116), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n263), .B1(new_n767), .B2(G326), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n780), .A2(new_n320), .B1(new_n255), .B2(new_n775), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n787), .A2(new_n392), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n791), .A2(new_n363), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n547), .B2(new_n770), .C1(new_n783), .C2(new_n369), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1036), .A2(new_n283), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n963), .B2(new_n851), .C1(new_n861), .C2(new_n764), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1035), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(KEYINPUT113), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1035), .A2(new_n1044), .A3(new_n1041), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n759), .A3(new_n1045), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n320), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1047), .A2(G116), .A3(new_n521), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT50), .B1(new_n320), .B2(G50), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n305), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G68), .B2(G77), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n978), .B(new_n1051), .C1(G45), .C2(new_n237), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n810), .A2(new_n709), .B1(G107), .B2(new_n205), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT112), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n808), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n807), .B1(new_n699), .B2(new_n700), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1046), .A2(new_n803), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n708), .B1(new_n1014), .B2(new_n757), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n757), .B2(new_n1014), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1013), .A2(new_n702), .A3(new_n802), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT111), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .ZN(G393));
  AOI21_X1  g0862(.A(new_n1021), .B1(new_n697), .B2(new_n701), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n702), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1063), .A2(new_n801), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n852), .A2(new_n783), .B1(new_n764), .B2(new_n952), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT52), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n851), .A2(new_n1028), .B1(new_n563), .B2(new_n788), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT116), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1068), .A2(new_n1069), .B1(new_n461), .B2(new_n770), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1067), .A2(new_n263), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n856), .A2(G116), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G303), .A2(new_n779), .B1(new_n776), .B2(G294), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G159), .A2(new_n784), .B1(new_n765), .B2(G150), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n856), .A2(G77), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n767), .A2(G143), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n864), .A2(G87), .B1(G68), .B2(new_n791), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n263), .B1(new_n369), .B2(new_n780), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n320), .B2(new_n775), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n760), .B1(new_n1075), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n814), .A2(new_n247), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n809), .B1(new_n706), .B2(G97), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n804), .B(new_n1086), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1000), .A2(new_n819), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT114), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1065), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1014), .A2(new_n757), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n707), .A3(new_n1022), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(G390));
  OAI211_X1 g0896(.A(new_n651), .B(new_n939), .C1(new_n737), .C2(new_n652), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n913), .B1(new_n756), .B2(new_n833), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n922), .A2(G330), .A3(new_n925), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n831), .B1(new_n734), .B2(new_n834), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n913), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n843), .A2(new_n834), .A3(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n727), .A2(new_n692), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n831), .B1(new_n1106), .B2(new_n830), .ZN(new_n1107));
  OAI211_X1 g0907(.A(G330), .B(new_n834), .C1(new_n755), .C2(new_n928), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n913), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1105), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1097), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n915), .B2(new_n896), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n896), .ZN(new_n1114));
  OAI211_X1 g0914(.A(KEYINPUT117), .B(new_n1114), .C1(new_n1101), .C2(new_n913), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n895), .B1(new_n894), .B2(new_n901), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1105), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n893), .B(new_n1114), .C1(new_n1107), .C2(new_n913), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1099), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1111), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1099), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n918), .A2(new_n940), .A3(new_n919), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1105), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1101), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1123), .A2(new_n1131), .A3(new_n707), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n801), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1116), .A2(new_n805), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n851), .A2(new_n490), .B1(new_n255), .B2(new_n770), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n783), .B2(new_n213), .C1(new_n547), .C2(new_n775), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G87), .B2(new_n791), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1079), .B1(new_n764), .B2(new_n563), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n263), .B(new_n1140), .C1(G107), .C2(new_n779), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n1136), .C2(new_n1135), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT119), .Z(new_n1143));
  NAND2_X1  g0943(.A1(new_n856), .A2(G159), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n283), .B1(new_n765), .B2(G128), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n788), .A2(new_n963), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT53), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(new_n369), .C2(new_n770), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT54), .B(G143), .Z(new_n1149));
  AOI22_X1  g0949(.A1(G137), .A2(new_n779), .B1(new_n776), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n867), .B2(new_n783), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1148), .B(new_n1151), .C1(G125), .C2(new_n767), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1143), .B1(new_n1144), .B2(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n803), .B1(new_n321), .B2(new_n872), .C1(new_n1153), .C2(new_n760), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1134), .A2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1133), .A2(KEYINPUT120), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n802), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1155), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1132), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT121), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT121), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1163), .B(new_n1132), .C1(new_n1156), .C2(new_n1160), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(G378));
  NAND2_X1  g0965(.A1(new_n384), .A2(new_n391), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  OR2_X1    g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n376), .A2(new_n876), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n376), .A3(new_n876), .A4(new_n1169), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n937), .A2(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n902), .A2(new_n903), .A3(new_n916), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n935), .A2(new_n1174), .A3(G330), .A4(new_n936), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1177), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1174), .A2(new_n805), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n803), .B1(G50), .B2(new_n872), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n369), .B1(new_n278), .B2(G41), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n770), .A2(new_n211), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n776), .B2(new_n524), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n213), .B2(new_n764), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1038), .B1(new_n783), .B2(new_n461), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n304), .B1(new_n851), .B2(new_n563), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n779), .A2(G97), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1190), .A2(new_n283), .A3(new_n967), .A4(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT58), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G128), .A2(new_n784), .B1(new_n765), .B2(G125), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n779), .A2(G132), .B1(new_n791), .B2(new_n1149), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n860), .B2(new_n775), .C1(new_n963), .C2(new_n787), .ZN(new_n1197));
  XOR2_X1   g0997(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1198));
  XOR2_X1   g0998(.A(new_n1197), .B(new_n1198), .Z(new_n1199));
  AOI21_X1  g0999(.A(G41), .B1(new_n767), .B2(G124), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n864), .A2(G159), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1200), .A2(new_n266), .A3(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1184), .B(new_n1193), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1183), .B1(new_n1203), .B2(new_n759), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1181), .A2(new_n802), .B1(new_n1182), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1129), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1206));
  OAI211_X1 g1006(.A(KEYINPUT57), .B(new_n1181), .C1(new_n1206), .C2(new_n1097), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n707), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1181), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1205), .B1(new_n1208), .B2(new_n1210), .ZN(G375));
  NOR2_X1   g1011(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(new_n801), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n913), .A2(new_n805), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n779), .A2(new_n1149), .B1(new_n784), .B2(G137), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n867), .B2(new_n764), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT123), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1185), .B(new_n1217), .C1(G150), .C2(new_n776), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n791), .A2(G159), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n767), .A2(G128), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n283), .B1(new_n856), .B2(G50), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n764), .A2(new_n490), .B1(new_n432), .B2(new_n770), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G116), .B2(new_n779), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n283), .B1(new_n851), .B2(new_n612), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1037), .B(new_n1225), .C1(G97), .C2(new_n791), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n461), .B2(new_n775), .C1(new_n563), .C2(new_n783), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n760), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n804), .B(new_n1229), .C1(new_n255), .C2(new_n871), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1213), .B1(new_n1214), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1212), .A2(new_n1097), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n1024), .A3(new_n1129), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(G381));
  INV_X1    g1034(.A(new_n1025), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n1009), .A3(new_n1008), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1236), .A2(new_n980), .A3(new_n1092), .A4(new_n1095), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n826), .B(KEYINPUT101), .Z(new_n1238));
  NAND4_X1  g1038(.A1(new_n1238), .A2(new_n1059), .A3(new_n1057), .A4(new_n1061), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1237), .A2(G384), .A3(G381), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1205), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1174), .B1(new_n932), .B2(G330), .ZN(new_n1242));
  AND4_X1   g1042(.A1(G330), .A2(new_n935), .A3(new_n1174), .A4(new_n936), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n917), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1126), .B2(new_n1123), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n708), .B1(new_n1247), .B2(KEYINPUT57), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1209), .A2(new_n1181), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT57), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1241), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1133), .A2(new_n1155), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1132), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1240), .A2(new_n1252), .A3(new_n1255), .ZN(G407));
  NOR2_X1   g1056(.A1(new_n1240), .A2(new_n690), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1258));
  OAI21_X1  g1058(.A(G213), .B1(new_n1257), .B2(new_n1258), .ZN(G409));
  INV_X1    g1059(.A(G213), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(G343), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n708), .B1(new_n1232), .B2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n1129), .C1(new_n1263), .C2(new_n1232), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1231), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(G384), .A3(new_n1231), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G375), .B1(new_n1164), .B2(new_n1162), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1247), .A2(new_n1024), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1254), .B1(new_n1273), .B2(new_n1205), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1262), .B(new_n1271), .C1(new_n1272), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT62), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1261), .A2(G2897), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1268), .A2(new_n1269), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1278), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1270), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1274), .B1(G378), .B2(new_n1252), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1279), .B(new_n1281), .C1(new_n1282), .C2(new_n1261), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1164), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT120), .B1(new_n1133), .B2(new_n1155), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1158), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1163), .B1(new_n1287), .B2(new_n1132), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1252), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1274), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1262), .A4(new_n1271), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1276), .A2(new_n1277), .A3(new_n1283), .A4(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(G390), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1237), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G393), .A2(G396), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1239), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1239), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1239), .B2(new_n1297), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1237), .B(new_n1295), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1294), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1261), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1281), .A2(new_n1279), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1306), .B(new_n1307), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1261), .B(new_n1270), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT63), .B1(new_n1312), .B2(KEYINPUT124), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT124), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1275), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1311), .A2(new_n1313), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1305), .A2(new_n1317), .ZN(G405));
  NAND2_X1  g1118(.A1(G375), .A2(new_n1255), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1289), .A2(KEYINPUT127), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1271), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1304), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1306), .A2(new_n1320), .A3(new_n1271), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1289), .A2(new_n1319), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1322), .A2(new_n1326), .A3(new_n1325), .A4(new_n1323), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


