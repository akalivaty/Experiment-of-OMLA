//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT64), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT0), .B(G128), .Z(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  OAI211_X1 g005(.A(KEYINPUT0), .B(G128), .C1(new_n188), .C2(KEYINPUT64), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n198), .B(new_n188), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n194), .B1(G125), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G953), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G224), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n200), .B(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT3), .A3(G107), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT81), .A2(G104), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G107), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G107), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n206), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT84), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(new_n217), .A3(new_n214), .A4(G101), .ZN(new_n218));
  INV_X1    g032(.A(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT67), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n223), .B2(new_n224), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n216), .A2(new_n218), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n214), .B1(new_n213), .B2(G101), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n210), .A2(new_n233), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n232), .A2(KEYINPUT82), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n236));
  INV_X1    g050(.A(G107), .ZN(new_n237));
  INV_X1    g051(.A(new_n209), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT81), .A2(G104), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n205), .B1(new_n240), .B2(KEYINPUT3), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n238), .A2(new_n239), .ZN(new_n242));
  AOI21_X1  g056(.A(G101), .B1(new_n242), .B2(G107), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n230), .B(new_n231), .C1(new_n235), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT82), .B1(new_n232), .B2(new_n234), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n236), .A3(new_n243), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n231), .B1(new_n249), .B2(new_n230), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n229), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n224), .A2(KEYINPUT5), .ZN(new_n252));
  INV_X1    g066(.A(G116), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n253), .A2(KEYINPUT5), .A3(G119), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(new_n219), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n228), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT85), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n204), .A2(G107), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n233), .B1(new_n240), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n259), .B1(new_n249), .B2(new_n262), .ZN(new_n263));
  AOI211_X1 g077(.A(KEYINPUT85), .B(new_n261), .C1(new_n247), .C2(new_n248), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G122), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n251), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT87), .A2(KEYINPUT6), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n251), .A2(new_n265), .ZN(new_n271));
  INV_X1    g085(.A(new_n266), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n266), .B1(new_n251), .B2(new_n265), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n269), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n203), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n266), .B(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n249), .A2(new_n262), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT85), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n261), .B1(new_n247), .B2(new_n248), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n259), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n257), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n258), .A2(new_n281), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n202), .A2(KEYINPUT7), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n200), .B(new_n286), .Z(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n267), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n277), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n203), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n275), .B1(new_n269), .B2(new_n267), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n266), .B(new_n268), .C1(new_n251), .C2(new_n265), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n288), .A2(new_n289), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT88), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n291), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n274), .A2(new_n276), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n290), .B1(new_n301), .B2(new_n292), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT89), .B1(new_n302), .B2(new_n298), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n291), .A2(new_n297), .A3(KEYINPUT89), .A4(new_n299), .ZN(new_n306));
  XNOR2_X1  g120(.A(G113), .B(G122), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(new_n204), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT70), .B(G953), .ZN(new_n309));
  INV_X1    g123(.A(G237), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(G214), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT90), .ZN(new_n312));
  INV_X1    g126(.A(G143), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT90), .B(G143), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n309), .A2(new_n315), .A3(G214), .A4(new_n310), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT18), .ZN(new_n317));
  INV_X1    g131(.A(G131), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n314), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(new_n196), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n319), .B(new_n321), .C1(new_n323), .C2(new_n317), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT17), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n314), .A2(new_n318), .A3(new_n316), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n322), .A2(KEYINPUT17), .A3(G131), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n320), .A2(KEYINPUT16), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n330), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(G146), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(G146), .B1(new_n329), .B2(new_n331), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT91), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n334), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT91), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n332), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n328), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n308), .B(new_n324), .C1(new_n327), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n308), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n319), .A2(new_n321), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n317), .B(new_n318), .C1(new_n314), .C2(new_n316), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT19), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n320), .B(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n332), .B1(new_n346), .B2(G146), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n323), .B2(new_n326), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n341), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(G475), .A2(G902), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT20), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(G234), .A2(G237), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n357), .A2(G952), .A3(new_n201), .ZN(new_n358));
  INV_X1    g172(.A(new_n309), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(G902), .A3(new_n357), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n360), .B(KEYINPUT93), .Z(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT21), .B(G898), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n365), .A2(new_n366), .A3(G953), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n313), .A2(G128), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n195), .A2(G143), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G134), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G116), .B(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n237), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n253), .A2(KEYINPUT14), .A3(G122), .ZN(new_n376));
  INV_X1    g190(.A(new_n374), .ZN(new_n377));
  OAI211_X1 g191(.A(G107), .B(new_n376), .C1(new_n377), .C2(KEYINPUT14), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT92), .ZN(new_n380));
  INV_X1    g194(.A(new_n369), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n381), .A2(KEYINPUT13), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n370), .B1(new_n381), .B2(KEYINPUT13), .ZN(new_n383));
  OAI21_X1  g197(.A(G134), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n371), .A2(new_n372), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n374), .B(new_n237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n379), .A2(new_n380), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n380), .B1(new_n379), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n368), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n379), .A2(new_n387), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT92), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n367), .A3(new_n388), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n394), .A3(new_n289), .ZN(new_n395));
  INV_X1    g209(.A(G478), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(KEYINPUT15), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n395), .B(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n340), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n401), .A2(new_n328), .A3(new_n335), .A4(new_n338), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n308), .B1(new_n402), .B2(new_n324), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n289), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G475), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n356), .A2(new_n364), .A3(new_n399), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT94), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n353), .A2(new_n355), .B1(G475), .B2(new_n404), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT94), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n364), .A4(new_n399), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G110), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n195), .A2(G119), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT23), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n418));
  INV_X1    g232(.A(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G128), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n414), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n423), .B1(new_n422), .B2(new_n421), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n415), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT24), .B(G110), .ZN(new_n426));
  OAI221_X1 g240(.A(new_n424), .B1(new_n333), .B2(new_n334), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n320), .A2(new_n196), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n332), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n426), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT77), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n417), .A2(new_n418), .A3(new_n414), .A4(new_n420), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT77), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT78), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n432), .A2(KEYINPUT78), .A3(new_n433), .A4(new_n434), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n429), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT79), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI211_X1 g255(.A(KEYINPUT79), .B(new_n429), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n427), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G137), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n427), .B(new_n446), .C1(new_n441), .C2(new_n442), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n289), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n448), .A2(KEYINPUT25), .A3(new_n289), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n366), .B1(G234), .B2(new_n289), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(G902), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n449), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n460));
  INV_X1    g274(.A(G137), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT11), .A3(G134), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n372), .A2(G137), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT11), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n372), .B2(G137), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n464), .A2(KEYINPUT65), .A3(new_n318), .A4(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n466), .A2(new_n462), .A3(new_n318), .A4(new_n463), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n462), .A3(new_n463), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n467), .A2(new_n470), .B1(G131), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT68), .B1(new_n472), .B2(new_n193), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(G131), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n468), .A2(new_n469), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n468), .A2(new_n469), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n191), .A2(new_n192), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT68), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n461), .A2(G134), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n318), .B1(new_n481), .B2(new_n463), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n467), .B2(new_n470), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n199), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n473), .A2(new_n480), .A3(KEYINPUT30), .A4(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n472), .A2(new_n193), .ZN(new_n486));
  INV_X1    g300(.A(new_n199), .ZN(new_n487));
  INV_X1    g301(.A(new_n482), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n475), .B2(new_n476), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n483), .A2(KEYINPUT66), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n486), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n460), .B(new_n485), .C1(new_n493), .C2(KEYINPUT30), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n460), .B1(new_n483), .B2(new_n199), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n473), .A2(new_n480), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n473), .A2(new_n480), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n309), .A2(G210), .A3(new_n310), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT72), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(G101), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n503), .B(new_n506), .Z(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT73), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n501), .A2(new_n512), .A3(new_n508), .ZN(new_n513));
  INV_X1    g327(.A(new_n486), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT28), .B1(new_n514), .B2(new_n495), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n491), .A2(new_n492), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n514), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n499), .A2(new_n497), .B1(new_n518), .B2(new_n460), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n507), .B(new_n516), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n510), .A2(new_n511), .A3(new_n513), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n473), .A2(new_n480), .A3(new_n484), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n460), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(KEYINPUT74), .A3(new_n460), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n500), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n515), .B1(new_n528), .B2(KEYINPUT28), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n508), .A2(new_n511), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n522), .B1(new_n531), .B2(KEYINPUT75), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n533), .B(G902), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  OAI21_X1  g348(.A(G472), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT31), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n494), .A2(new_n500), .A3(new_n536), .A4(new_n507), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n494), .A2(new_n500), .A3(new_n507), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT31), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n518), .A2(new_n460), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n500), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n515), .B1(new_n541), .B2(KEYINPUT28), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n537), .B(new_n539), .C1(new_n542), .C2(new_n507), .ZN(new_n543));
  NOR2_X1   g357(.A1(G472), .A2(G902), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n543), .A2(KEYINPUT32), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT32), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n459), .B1(new_n535), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n193), .B1(new_n216), .B2(new_n218), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n246), .B2(new_n250), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n487), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n263), .B2(new_n264), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n281), .A2(new_n199), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n551), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n550), .A2(new_n553), .A3(new_n472), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n309), .A2(G227), .ZN(new_n557));
  XOR2_X1   g371(.A(G110), .B(G140), .Z(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n280), .A2(new_n282), .A3(new_n487), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n554), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(KEYINPUT86), .A3(new_n564), .A4(new_n477), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n564), .A2(KEYINPUT86), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(KEYINPUT86), .ZN(new_n567));
  INV_X1    g381(.A(new_n554), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n263), .A2(new_n264), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(new_n569), .B2(new_n487), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(new_n567), .C1(new_n570), .C2(new_n472), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n230), .B1(new_n235), .B2(new_n244), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT83), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n245), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n575), .A2(new_n549), .B1(new_n551), .B2(new_n554), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n472), .B1(new_n576), .B2(new_n553), .ZN(new_n577));
  INV_X1    g391(.A(new_n556), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n559), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G469), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n289), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n571), .A2(new_n556), .A3(new_n565), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n559), .ZN(new_n584));
  INV_X1    g398(.A(new_n577), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n561), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(G469), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n581), .A2(new_n289), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n582), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G221), .B1(new_n365), .B2(G902), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT80), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n413), .A2(new_n548), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n543), .B2(new_n289), .ZN(new_n599));
  INV_X1    g413(.A(new_n544), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n539), .A2(new_n537), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n508), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n459), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n590), .A3(new_n606), .A4(new_n593), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n305), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n298), .B1(new_n295), .B2(new_n296), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(KEYINPUT95), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n299), .B1(new_n277), .B2(new_n290), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n391), .A2(new_n394), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n391), .A2(new_n394), .A3(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n396), .A2(G902), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n620), .A2(new_n621), .B1(new_n396), .B2(new_n395), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n408), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g437(.A1(new_n364), .A2(new_n611), .A3(new_n615), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n608), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n356), .A2(KEYINPUT96), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT96), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n353), .A2(new_n629), .A3(new_n355), .ZN(new_n630));
  INV_X1    g444(.A(new_n399), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n628), .A2(new_n630), .A3(new_n405), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n363), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n633), .A2(new_n611), .A3(new_n615), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n608), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NOR2_X1   g451(.A1(new_n447), .A2(KEYINPUT36), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT97), .Z(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(new_n443), .Z(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n457), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n456), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n605), .A2(new_n590), .A3(new_n593), .A4(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n412), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  AOI22_X1  g460(.A1(new_n454), .A2(new_n455), .B1(new_n640), .B2(new_n457), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n535), .B2(new_n547), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n611), .A2(new_n615), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n358), .B1(new_n361), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n648), .A2(new_n595), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  NAND2_X1  g469(.A1(new_n304), .A2(new_n306), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT38), .Z(new_n657));
  XOR2_X1   g471(.A(new_n652), .B(KEYINPUT39), .Z(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n594), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT40), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n408), .A2(new_n399), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n647), .A2(new_n305), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT98), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n604), .A2(KEYINPUT32), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n543), .A2(new_n544), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT32), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n289), .B1(new_n528), .B2(new_n507), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n508), .B1(new_n494), .B2(new_n500), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n664), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n657), .A2(new_n661), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n408), .A2(new_n622), .A3(new_n652), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n677), .B1(new_n649), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n611), .A2(new_n615), .A3(KEYINPUT99), .A4(new_n678), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n680), .A2(new_n595), .A3(new_n648), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  AOI21_X1  g497(.A(G902), .B1(new_n572), .B2(new_n579), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n581), .ZN(new_n685));
  AOI211_X1 g499(.A(G469), .B(G902), .C1(new_n572), .C2(new_n579), .ZN(new_n686));
  INV_X1    g500(.A(new_n591), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n624), .A2(new_n548), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT41), .B(G113), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT100), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n689), .B(new_n691), .ZN(G15));
  NAND3_X1  g506(.A1(new_n634), .A2(new_n548), .A3(new_n688), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  INV_X1    g508(.A(new_n648), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n688), .A2(new_n411), .A3(new_n615), .A4(new_n611), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT101), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n580), .A2(new_n289), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n591), .A3(new_n582), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n407), .A2(new_n410), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n649), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n648), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n611), .A2(new_n615), .A3(new_n662), .ZN(new_n708));
  NOR4_X1   g522(.A1(new_n685), .A2(new_n686), .A3(new_n687), .A4(new_n363), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n539), .B1(new_n529), .B2(new_n507), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT102), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n713), .B(new_n539), .C1(new_n529), .C2(new_n507), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n537), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n544), .ZN(new_n716));
  INV_X1    g530(.A(new_n599), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n606), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n707), .B1(new_n710), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n611), .A2(new_n615), .A3(new_n662), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n699), .A2(new_n591), .A3(new_n582), .A4(new_n364), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n599), .B(new_n459), .C1(new_n715), .C2(new_n544), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(KEYINPUT103), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR2_X1   g540(.A1(new_n649), .A2(new_n700), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n599), .B(new_n647), .C1(new_n715), .C2(new_n544), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n678), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  XNOR2_X1  g544(.A(new_n588), .B(KEYINPUT104), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n684), .B2(new_n581), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n687), .B1(new_n733), .B2(new_n587), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n656), .A2(new_n305), .A3(new_n678), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n604), .B2(KEYINPUT32), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n546), .A2(KEYINPUT105), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n665), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n535), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n606), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT42), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n609), .B1(new_n304), .B2(new_n306), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n679), .A2(KEYINPUT42), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n548), .A3(new_n734), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n318), .ZN(G33));
  NAND4_X1  g561(.A1(new_n743), .A2(new_n548), .A3(new_n653), .A4(new_n734), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND2_X1  g563(.A1(new_n356), .A2(new_n405), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n750), .B2(new_n622), .ZN(new_n751));
  INV_X1    g565(.A(new_n622), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n408), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n647), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n605), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(KEYINPUT44), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n758), .A2(new_n762), .A3(KEYINPUT44), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT44), .B1(new_n758), .B2(new_n759), .ZN(new_n765));
  INV_X1    g579(.A(new_n743), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n583), .A2(new_n559), .B1(new_n585), .B2(new_n561), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT45), .ZN(new_n769));
  OAI21_X1  g583(.A(G469), .B1(new_n768), .B2(KEYINPUT45), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n731), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n686), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n687), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n775), .A2(new_n658), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n776), .B1(new_n775), .B2(new_n658), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n764), .B(new_n767), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  XNOR2_X1  g594(.A(new_n775), .B(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n535), .A2(new_n547), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n782), .A2(new_n606), .A3(new_n679), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n743), .A3(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT110), .B(G140), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G42));
  NOR3_X1   g600(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT101), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n703), .B1(new_n702), .B2(new_n648), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(new_n707), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT103), .B1(new_n722), .B2(new_n723), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n548), .B(new_n688), .C1(new_n624), .C2(new_n634), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n750), .A2(new_n622), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n408), .A2(new_n399), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n793), .A2(new_n364), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n304), .A2(new_n305), .A3(new_n795), .A4(new_n306), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(new_n607), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n596), .A2(new_n792), .A3(new_n644), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n582), .A2(new_n587), .A3(new_n731), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n591), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n720), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n642), .A2(new_n652), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n672), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT114), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n802), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n654), .A2(new_n729), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n811), .A3(new_n812), .A4(new_n682), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n802), .A2(new_n804), .A3(new_n807), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n807), .B1(new_n802), .B2(new_n804), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n682), .A2(new_n654), .A3(new_n729), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT52), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n743), .A2(new_n728), .A3(new_n678), .A4(new_n734), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n628), .A2(new_n405), .A3(new_n630), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n631), .A3(new_n652), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n743), .A2(new_n648), .A3(new_n595), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n748), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n746), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n799), .A2(new_n813), .A3(new_n818), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n782), .A2(new_n606), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n412), .A3(new_n594), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n412), .A2(new_n643), .B1(new_n796), .B2(new_n607), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n705), .A3(new_n725), .A4(new_n792), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n748), .A2(new_n822), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n742), .A3(new_n745), .A4(new_n819), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT53), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n835), .A2(new_n813), .A3(new_n818), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n827), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n827), .A2(new_n839), .A3(new_n841), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT115), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n836), .A2(new_n826), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n835), .A2(new_n813), .A3(new_n818), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n841), .B1(new_n827), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n842), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(new_n842), .C1(new_n844), .C2(new_n847), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n743), .A2(new_n688), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n606), .A2(new_n358), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n852), .A2(new_n672), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n408), .A3(new_n622), .ZN(new_n855));
  INV_X1    g669(.A(new_n852), .ZN(new_n856));
  INV_X1    g670(.A(new_n755), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n358), .A3(new_n728), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n688), .A2(new_n609), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT117), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n656), .B(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n358), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n718), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n859), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n685), .A2(new_n686), .A3(new_n593), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n743), .B(new_n864), .C1(new_n781), .C2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT51), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n852), .A2(new_n741), .A3(new_n863), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT48), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n854), .A2(new_n623), .ZN(new_n875));
  INV_X1    g689(.A(G952), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n876), .B(G953), .C1(new_n864), .C2(new_n727), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n871), .A3(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT118), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n869), .A2(new_n871), .A3(new_n881), .A4(KEYINPUT51), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n872), .B(new_n878), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n849), .A2(new_n851), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n876), .A2(new_n201), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n750), .A2(new_n622), .A3(new_n592), .A4(new_n609), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n606), .A2(new_n887), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT111), .Z(new_n889));
  INV_X1    g703(.A(KEYINPUT49), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n685), .A2(new_n686), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT112), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n672), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n862), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT113), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n896), .ZN(G75));
  NAND2_X1  g711(.A1(new_n827), .A2(new_n839), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n289), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n301), .A2(new_n292), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n277), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n309), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n900), .B2(G210), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n911), .B1(new_n912), .B2(new_n906), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n901), .A2(new_n902), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(KEYINPUT119), .A3(new_n905), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n913), .B2(new_n915), .ZN(G51));
  XNOR2_X1  g730(.A(new_n898), .B(new_n841), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n731), .B(KEYINPUT57), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n580), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n769), .A2(new_n770), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n900), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n919), .B2(new_n921), .ZN(G54));
  NAND3_X1  g736(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n923));
  INV_X1    g737(.A(new_n350), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n908), .ZN(G60));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n620), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n909), .B1(new_n917), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n851), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n827), .A2(new_n846), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT54), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(KEYINPUT115), .A3(new_n843), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n850), .B1(new_n936), .B2(new_n842), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n930), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n620), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n898), .A2(new_n640), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n448), .A2(new_n449), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n899), .B2(new_n942), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n898), .A2(new_n948), .A3(new_n640), .A4(new_n943), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n947), .A3(new_n909), .A4(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT61), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT61), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  INV_X1    g768(.A(new_n362), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n201), .B1(new_n955), .B2(G224), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n832), .B2(new_n309), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n274), .B(new_n276), .C1(G898), .C2(new_n309), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT122), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n957), .B(new_n959), .ZN(G69));
  NAND2_X1  g774(.A1(new_n779), .A2(new_n784), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n741), .A2(new_n720), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n777), .B2(new_n778), .ZN(new_n963));
  INV_X1    g777(.A(new_n748), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n746), .A2(new_n964), .A3(new_n817), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n961), .A2(new_n966), .A3(KEYINPUT125), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT125), .B1(new_n961), .B2(new_n966), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n309), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n485), .B1(new_n493), .B2(KEYINPUT30), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(new_n346), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n969), .B(new_n971), .C1(new_n651), .C2(new_n309), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n675), .A2(new_n682), .A3(new_n811), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n793), .A2(new_n794), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n660), .A2(new_n743), .A3(new_n548), .A4(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n779), .A2(new_n784), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT124), .B1(new_n973), .B2(KEYINPUT62), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n973), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n978), .B(new_n979), .C1(new_n980), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n309), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n971), .B(KEYINPUT123), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n972), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n309), .B1(G227), .B2(G900), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n988), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n972), .A2(new_n990), .A3(new_n986), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(G72));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n983), .B2(new_n832), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n670), .ZN(new_n997));
  INV_X1    g811(.A(new_n995), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n510), .A2(new_n513), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n999), .A2(KEYINPUT126), .ZN(new_n1000));
  INV_X1    g814(.A(new_n538), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n999), .B2(KEYINPUT126), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n998), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n908), .B1(new_n934), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n967), .A2(new_n799), .A3(new_n968), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n507), .B(new_n501), .C1(new_n1006), .C2(new_n995), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n993), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n995), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1009), .A2(new_n508), .A3(new_n500), .A4(new_n494), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1010), .A2(KEYINPUT127), .A3(new_n997), .A4(new_n1004), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n1011), .ZN(G57));
endmodule


