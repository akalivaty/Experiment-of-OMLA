

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(n322), .B(n321), .ZN(n324) );
  XNOR2_X1 U326 ( .A(n329), .B(n295), .ZN(n330) );
  XNOR2_X1 U327 ( .A(n366), .B(n413), .ZN(n353) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  AND2_X1 U329 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U330 ( .A(n384), .B(KEYINPUT64), .Z(n295) );
  XNOR2_X1 U331 ( .A(KEYINPUT104), .B(KEYINPUT47), .ZN(n456) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U333 ( .A(G197GAT), .ZN(n351) );
  XNOR2_X1 U334 ( .A(n460), .B(KEYINPUT48), .ZN(n517) );
  XNOR2_X1 U335 ( .A(n320), .B(n293), .ZN(n321) );
  XNOR2_X1 U336 ( .A(n352), .B(n351), .ZN(n366) );
  XNOR2_X1 U337 ( .A(n461), .B(KEYINPUT118), .ZN(n462) );
  XNOR2_X1 U338 ( .A(n355), .B(n294), .ZN(n356) );
  XNOR2_X1 U339 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U340 ( .A(n463), .B(n462), .ZN(n570) );
  NOR2_X1 U341 ( .A1(n584), .A2(n408), .ZN(n409) );
  XNOR2_X1 U342 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U343 ( .A(n443), .B(n442), .ZN(n576) );
  XNOR2_X1 U344 ( .A(n331), .B(n330), .ZN(n473) );
  XOR2_X1 U345 ( .A(KEYINPUT41), .B(n452), .Z(n561) );
  NOR2_X1 U346 ( .A1(n527), .A2(n526), .ZN(n536) );
  XNOR2_X1 U347 ( .A(n361), .B(n436), .ZN(n509) );
  XNOR2_X1 U348 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n447) );
  XNOR2_X1 U350 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  XNOR2_X1 U351 ( .A(n448), .B(n447), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n297) );
  XNOR2_X1 U353 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n315) );
  XOR2_X1 U355 ( .A(KEYINPUT65), .B(G190GAT), .Z(n299) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G15GAT), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n301) );
  XOR2_X1 U358 ( .A(G134GAT), .B(G99GAT), .Z(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n311) );
  XOR2_X1 U360 ( .A(G183GAT), .B(KEYINPUT19), .Z(n303) );
  XNOR2_X1 U361 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n359) );
  XOR2_X1 U363 ( .A(G127GAT), .B(KEYINPUT82), .Z(n305) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n393) );
  XNOR2_X1 U366 ( .A(n359), .B(n393), .ZN(n309) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G176GAT), .Z(n307) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(G71GAT), .ZN(n306) );
  XNOR2_X1 U369 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n313) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n523) );
  XOR2_X1 U375 ( .A(G99GAT), .B(G85GAT), .Z(n437) );
  XOR2_X1 U376 ( .A(G36GAT), .B(G190GAT), .Z(n355) );
  XOR2_X1 U377 ( .A(n437), .B(n355), .Z(n317) );
  XNOR2_X1 U378 ( .A(G162GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n322) );
  XOR2_X1 U380 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n319) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(G92GAT), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n320) );
  INV_X1 U383 ( .A(KEYINPUT10), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n331) );
  XOR2_X1 U385 ( .A(KEYINPUT7), .B(KEYINPUT71), .Z(n326) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(G43GAT), .ZN(n325) );
  XNOR2_X1 U387 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U388 ( .A(KEYINPUT8), .B(n327), .ZN(n424) );
  INV_X1 U389 ( .A(n424), .ZN(n329) );
  XNOR2_X1 U390 ( .A(G29GAT), .B(G134GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n328), .B(KEYINPUT77), .ZN(n384) );
  INV_X1 U392 ( .A(n473), .ZN(n551) );
  XOR2_X1 U393 ( .A(KEYINPUT36), .B(n551), .Z(n584) );
  XOR2_X1 U394 ( .A(G71GAT), .B(KEYINPUT13), .Z(n434) );
  XOR2_X1 U395 ( .A(G78GAT), .B(G211GAT), .Z(n333) );
  XNOR2_X1 U396 ( .A(G183GAT), .B(G155GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U398 ( .A(n434), .B(n334), .Z(n336) );
  NAND2_X1 U399 ( .A1(G231GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U401 ( .A(n337), .B(KEYINPUT79), .Z(n340) );
  XNOR2_X1 U402 ( .A(G22GAT), .B(G15GAT), .ZN(n338) );
  XNOR2_X1 U403 ( .A(n338), .B(G1GAT), .ZN(n416) );
  XNOR2_X1 U404 ( .A(n416), .B(KEYINPUT78), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n348) );
  XOR2_X1 U406 ( .A(G64GAT), .B(G57GAT), .Z(n342) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(G127GAT), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U409 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n344) );
  XNOR2_X1 U410 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U412 ( .A(n346), .B(n345), .Z(n347) );
  XOR2_X1 U413 ( .A(n348), .B(n347), .Z(n564) );
  INV_X1 U414 ( .A(n564), .ZN(n580) );
  XOR2_X1 U415 ( .A(KEYINPUT92), .B(G204GAT), .Z(n354) );
  XOR2_X1 U416 ( .A(KEYINPUT21), .B(G218GAT), .Z(n350) );
  XNOR2_X1 U417 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U418 ( .A(n350), .B(n349), .ZN(n352) );
  XOR2_X1 U419 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G92GAT), .ZN(n360) );
  XOR2_X1 U423 ( .A(n360), .B(G64GAT), .Z(n436) );
  XNOR2_X1 U424 ( .A(KEYINPUT27), .B(n509), .ZN(n516) );
  XNOR2_X1 U425 ( .A(G155GAT), .B(KEYINPUT87), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n362), .B(KEYINPUT2), .ZN(n363) );
  XOR2_X1 U427 ( .A(n363), .B(KEYINPUT3), .Z(n365) );
  XNOR2_X1 U428 ( .A(G141GAT), .B(G162GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n385) );
  XNOR2_X1 U430 ( .A(n385), .B(n366), .ZN(n378) );
  XOR2_X1 U431 ( .A(G148GAT), .B(KEYINPUT24), .Z(n368) );
  XNOR2_X1 U432 ( .A(G50GAT), .B(G22GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n371) );
  XOR2_X1 U434 ( .A(G78GAT), .B(G204GAT), .Z(n370) );
  XNOR2_X1 U435 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n430) );
  XOR2_X1 U437 ( .A(n371), .B(n430), .Z(n376) );
  XOR2_X1 U438 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n373) );
  NAND2_X1 U439 ( .A1(G228GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U441 ( .A(KEYINPUT23), .B(n374), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n464) );
  XOR2_X1 U444 ( .A(n464), .B(KEYINPUT66), .Z(n379) );
  XNOR2_X1 U445 ( .A(KEYINPUT28), .B(n379), .ZN(n527) );
  NOR2_X1 U446 ( .A1(n523), .A2(n527), .ZN(n396) );
  XOR2_X1 U447 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n381) );
  XNOR2_X1 U448 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U450 ( .A(G85GAT), .B(KEYINPUT89), .Z(n382) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n389) );
  XOR2_X1 U452 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n387) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n391) );
  NAND2_X1 U456 ( .A1(G225GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U459 ( .A(G120GAT), .B(G148GAT), .Z(n394) );
  XOR2_X1 U460 ( .A(G57GAT), .B(n394), .Z(n431) );
  XOR2_X1 U461 ( .A(n395), .B(n431), .Z(n404) );
  XNOR2_X1 U462 ( .A(KEYINPUT91), .B(n404), .ZN(n518) );
  NAND2_X1 U463 ( .A1(n396), .A2(n518), .ZN(n399) );
  NOR2_X1 U464 ( .A1(n523), .A2(n464), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n397), .B(KEYINPUT26), .ZN(n571) );
  NAND2_X1 U466 ( .A1(n571), .A2(n404), .ZN(n398) );
  NAND2_X1 U467 ( .A1(n399), .A2(n398), .ZN(n400) );
  NAND2_X1 U468 ( .A1(n516), .A2(n400), .ZN(n407) );
  NAND2_X1 U469 ( .A1(n523), .A2(n509), .ZN(n401) );
  XOR2_X1 U470 ( .A(KEYINPUT93), .B(n401), .Z(n402) );
  NAND2_X1 U471 ( .A1(n464), .A2(n402), .ZN(n403) );
  XNOR2_X1 U472 ( .A(KEYINPUT25), .B(n403), .ZN(n405) );
  NAND2_X1 U473 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U474 ( .A1(n407), .A2(n406), .ZN(n476) );
  NAND2_X1 U475 ( .A1(n580), .A2(n476), .ZN(n408) );
  XNOR2_X1 U476 ( .A(KEYINPUT37), .B(n409), .ZN(n507) );
  XOR2_X1 U477 ( .A(KEYINPUT69), .B(G113GAT), .Z(n411) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(G197GAT), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U480 ( .A(n412), .B(G36GAT), .Z(n415) );
  XNOR2_X1 U481 ( .A(n413), .B(G29GAT), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U483 ( .A(n416), .B(KEYINPUT29), .Z(n418) );
  NAND2_X1 U484 ( .A1(G229GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U485 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U486 ( .A(n420), .B(n419), .Z(n426) );
  XOR2_X1 U487 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n422) );
  XNOR2_X1 U488 ( .A(KEYINPUT68), .B(KEYINPUT70), .ZN(n421) );
  XNOR2_X1 U489 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U490 ( .A(n424), .B(n423), .Z(n425) );
  XOR2_X1 U491 ( .A(n426), .B(n425), .Z(n573) );
  INV_X1 U492 ( .A(n573), .ZN(n556) );
  XOR2_X1 U493 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n428) );
  NAND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U496 ( .A(n429), .B(KEYINPUT76), .Z(n433) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U499 ( .A(n435), .B(n434), .Z(n443) );
  XOR2_X1 U500 ( .A(n437), .B(n436), .Z(n441) );
  XOR2_X1 U501 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n439) );
  XNOR2_X1 U502 ( .A(KEYINPUT31), .B(KEYINPUT74), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U504 ( .A1(n556), .A2(n576), .ZN(n478) );
  NOR2_X1 U505 ( .A1(n507), .A2(n478), .ZN(n445) );
  XNOR2_X1 U506 ( .A(KEYINPUT98), .B(KEYINPUT38), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U508 ( .A(KEYINPUT97), .B(n446), .Z(n492) );
  NAND2_X1 U509 ( .A1(n523), .A2(n492), .ZN(n448) );
  INV_X1 U510 ( .A(n576), .ZN(n452) );
  NOR2_X1 U511 ( .A1(n584), .A2(n580), .ZN(n449) );
  XOR2_X1 U512 ( .A(KEYINPUT45), .B(n449), .Z(n450) );
  NOR2_X1 U513 ( .A1(n452), .A2(n450), .ZN(n451) );
  NAND2_X1 U514 ( .A1(n451), .A2(n573), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n556), .A2(n561), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n453), .B(KEYINPUT46), .ZN(n455) );
  NOR2_X1 U517 ( .A1(n551), .A2(n564), .ZN(n454) );
  AND2_X1 U518 ( .A1(n455), .A2(n454), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n509), .A2(n517), .ZN(n463) );
  INV_X1 U521 ( .A(KEYINPUT54), .ZN(n461) );
  INV_X1 U522 ( .A(n518), .ZN(n569) );
  AND2_X1 U523 ( .A1(n569), .A2(n464), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n570), .A2(n465), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(KEYINPUT55), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n467), .A2(n523), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT119), .ZN(n565) );
  NAND2_X1 U528 ( .A1(n565), .A2(n551), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n470) );
  XNOR2_X1 U530 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n564), .A2(n473), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT81), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(KEYINPUT16), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n494) );
  NOR2_X1 U535 ( .A1(n494), .A2(n478), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n479), .B(KEYINPUT94), .ZN(n487) );
  NAND2_X1 U537 ( .A1(n487), .A2(n518), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NAND2_X1 U540 ( .A1(n487), .A2(n509), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT35), .B(KEYINPUT96), .Z(n484) );
  NAND2_X1 U543 ( .A1(n487), .A2(n523), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n486) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT95), .Z(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n487), .A2(n527), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U549 ( .A1(n518), .A2(n492), .ZN(n490) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n509), .A2(n492), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n527), .A2(n492), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT42), .Z(n496) );
  NAND2_X1 U557 ( .A1(n561), .A2(n573), .ZN(n506) );
  NOR2_X1 U558 ( .A1(n494), .A2(n506), .ZN(n501) );
  NAND2_X1 U559 ( .A1(n501), .A2(n518), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n497), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n509), .A2(n501), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(KEYINPUT100), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(n499), .ZN(G1333GAT) );
  NAND2_X1 U565 ( .A1(n523), .A2(n501), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U568 ( .A1(n501), .A2(n527), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(n505) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT102), .Z(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n507), .A2(n506), .ZN(n513) );
  NAND2_X1 U573 ( .A1(n518), .A2(n513), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  XOR2_X1 U575 ( .A(G92GAT), .B(KEYINPUT103), .Z(n511) );
  NAND2_X1 U576 ( .A1(n513), .A2(n509), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n523), .A2(n513), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U580 ( .A1(n527), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT44), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n515), .ZN(G1339GAT) );
  XOR2_X1 U583 ( .A(G113GAT), .B(KEYINPUT107), .Z(n529) );
  INV_X1 U584 ( .A(KEYINPUT106), .ZN(n525) );
  INV_X1 U585 ( .A(KEYINPUT105), .ZN(n522) );
  INV_X1 U586 ( .A(n516), .ZN(n520) );
  NAND2_X1 U587 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U588 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n540) );
  AND2_X1 U590 ( .A1(n540), .A2(n523), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U592 ( .A1(n536), .A2(n556), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT109), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U595 ( .A1(n536), .A2(n561), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT108), .Z(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n564), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT110), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n551), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n540), .A2(n571), .ZN(n541) );
  XNOR2_X1 U607 ( .A(KEYINPUT111), .B(n541), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n556), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT113), .Z(n544) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U613 ( .A(KEYINPUT112), .B(n545), .Z(n547) );
  NAND2_X1 U614 ( .A1(n552), .A2(n561), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n549) );
  NAND2_X1 U617 ( .A1(n552), .A2(n564), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n554) );
  NAND2_X1 U621 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n565), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n559) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U629 ( .A(KEYINPUT56), .B(n560), .Z(n563) );
  NAND2_X1 U630 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n575) );
  AND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n583) );
  NOR2_X1 U639 ( .A1(n573), .A2(n583), .ZN(n574) );
  XOR2_X1 U640 ( .A(n575), .B(n574), .Z(G1352GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n583), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(G204GAT), .B(n579), .Z(G1353GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n583), .ZN(n581) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(n581), .Z(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

