

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785;

  BUF_X1 U383 ( .A(G128), .Z(n396) );
  AND2_X1 U384 ( .A1(n377), .A2(n378), .ZN(n389) );
  XOR2_X2 U385 ( .A(n733), .B(n734), .Z(n735) );
  XNOR2_X2 U386 ( .A(n701), .B(KEYINPUT59), .ZN(n702) );
  XNOR2_X2 U387 ( .A(G902), .B(KEYINPUT15), .ZN(n640) );
  NOR2_X1 U388 ( .A1(n548), .A2(n547), .ZN(n714) );
  AND2_X2 U389 ( .A1(n644), .A2(n382), .ZN(n383) );
  INV_X2 U390 ( .A(n380), .ZN(n414) );
  XNOR2_X2 U391 ( .A(n388), .B(n411), .ZN(n380) );
  AND2_X2 U392 ( .A1(n389), .A2(n393), .ZN(n374) );
  NAND2_X2 U393 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X2 U394 ( .A(n607), .B(KEYINPUT19), .ZN(n581) );
  AND2_X1 U395 ( .A1(n548), .A2(n547), .ZN(n718) );
  NOR2_X1 U396 ( .A1(n589), .A2(n674), .ZN(n591) );
  AND2_X1 U397 ( .A1(n366), .A2(n364), .ZN(n363) );
  AND2_X1 U398 ( .A1(n394), .A2(n392), .ZN(n391) );
  NOR2_X2 U399 ( .A1(n589), .A2(n604), .ZN(n577) );
  XNOR2_X1 U400 ( .A(n549), .B(KEYINPUT101), .ZN(n672) );
  NOR2_X1 U401 ( .A1(n714), .A2(n718), .ZN(n549) );
  XNOR2_X1 U402 ( .A(n429), .B(KEYINPUT89), .ZN(n431) );
  NAND2_X1 U403 ( .A1(n452), .A2(G224), .ZN(n429) );
  INV_X1 U404 ( .A(G953), .ZN(n452) );
  NAND2_X1 U405 ( .A1(n363), .A2(n360), .ZN(n368) );
  NAND2_X1 U406 ( .A1(n362), .A2(n361), .ZN(n360) );
  AND2_X1 U407 ( .A1(n555), .A2(n554), .ZN(n556) );
  OR2_X1 U408 ( .A1(n782), .A2(n561), .ZN(n555) );
  NAND2_X1 U409 ( .A1(n395), .A2(n391), .ZN(n390) );
  XNOR2_X1 U410 ( .A(n418), .B(KEYINPUT40), .ZN(n785) );
  NOR2_X1 U411 ( .A1(n587), .A2(n586), .ZN(n588) );
  AND2_X1 U412 ( .A1(n409), .A2(KEYINPUT103), .ZN(n392) );
  OR2_X1 U413 ( .A1(KEYINPUT103), .A2(n409), .ZN(n378) );
  OR2_X1 U414 ( .A1(n426), .A2(n508), .ZN(n410) );
  NOR2_X1 U415 ( .A1(n661), .A2(n573), .ZN(n574) );
  AND2_X1 U416 ( .A1(n365), .A2(n647), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n567), .B(n496), .ZN(n658) );
  INV_X1 U418 ( .A(n373), .ZN(n361) );
  OR2_X1 U419 ( .A1(n373), .A2(G472), .ZN(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT75), .B(n471), .Z(n499) );
  INV_X4 U421 ( .A(n385), .ZN(n691) );
  XOR2_X1 U422 ( .A(KEYINPUT91), .B(KEYINPUT17), .Z(n430) );
  XOR2_X1 U423 ( .A(G113), .B(G116), .Z(n498) );
  NOR2_X2 U424 ( .A1(G953), .A2(G237), .ZN(n471) );
  XNOR2_X2 U425 ( .A(n529), .B(n528), .ZN(n698) );
  INV_X1 U426 ( .A(n383), .ZN(n362) );
  NAND2_X1 U427 ( .A1(n383), .A2(n367), .ZN(n366) );
  AND2_X1 U428 ( .A1(n373), .A2(G472), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U430 ( .A(n770), .B(n399), .ZN(n504) );
  INV_X1 U431 ( .A(G146), .ZN(n399) );
  NOR2_X1 U432 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U433 ( .A1(n404), .A2(n597), .ZN(n402) );
  NAND2_X1 U434 ( .A1(n405), .A2(KEYINPUT34), .ZN(n404) );
  XNOR2_X1 U435 ( .A(n421), .B(n420), .ZN(n510) );
  INV_X1 U436 ( .A(KEYINPUT8), .ZN(n420) );
  NAND2_X1 U437 ( .A1(G237), .A2(G234), .ZN(n450) );
  INV_X1 U438 ( .A(KEYINPUT88), .ZN(n424) );
  INV_X1 U439 ( .A(KEYINPUT22), .ZN(n411) );
  INV_X1 U440 ( .A(G116), .ZN(n439) );
  XNOR2_X1 U441 ( .A(n535), .B(KEYINPUT33), .ZN(n687) );
  XNOR2_X1 U442 ( .A(n470), .B(n469), .ZN(n548) );
  XNOR2_X1 U443 ( .A(n493), .B(n504), .ZN(n741) );
  INV_X1 U444 ( .A(G237), .ZN(n443) );
  XNOR2_X1 U445 ( .A(G131), .B(G143), .ZN(n474) );
  XNOR2_X1 U446 ( .A(n488), .B(n487), .ZN(n770) );
  XOR2_X1 U447 ( .A(G134), .B(G131), .Z(n487) );
  AND2_X1 U448 ( .A1(n658), .A2(n589), .ZN(n426) );
  XNOR2_X1 U449 ( .A(n495), .B(n494), .ZN(n567) );
  XNOR2_X1 U450 ( .A(KEYINPUT3), .B(G119), .ZN(n501) );
  XNOR2_X1 U451 ( .A(n396), .B(G110), .ZN(n513) );
  NAND2_X1 U452 ( .A1(n691), .A2(G227), .ZN(n489) );
  XOR2_X1 U453 ( .A(G107), .B(G104), .Z(n490) );
  OR2_X2 U454 ( .A1(n613), .A2(n675), .ZN(n419) );
  AND2_X1 U455 ( .A1(n449), .A2(n424), .ZN(n422) );
  XNOR2_X1 U456 ( .A(n417), .B(KEYINPUT97), .ZN(n592) );
  AND2_X1 U457 ( .A1(n544), .A2(n567), .ZN(n417) );
  XNOR2_X1 U458 ( .A(n466), .B(n465), .ZN(n745) );
  XNOR2_X1 U459 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U460 ( .A(KEYINPUT80), .ZN(n653) );
  NAND2_X1 U461 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U462 ( .A1(n690), .A2(n427), .ZN(n692) );
  XNOR2_X1 U463 ( .A(n539), .B(n538), .ZN(n782) );
  XNOR2_X1 U464 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U465 ( .A(n741), .B(n740), .ZN(n742) );
  INV_X1 U466 ( .A(n412), .ZN(n551) );
  AND2_X1 U467 ( .A1(n526), .A2(n525), .ZN(n369) );
  AND2_X1 U468 ( .A1(n537), .A2(n406), .ZN(n370) );
  OR2_X1 U469 ( .A1(n449), .A2(n424), .ZN(n371) );
  INV_X1 U470 ( .A(KEYINPUT66), .ZN(n508) );
  INV_X1 U471 ( .A(KEYINPUT103), .ZN(n523) );
  AND2_X1 U472 ( .A1(KEYINPUT66), .A2(n523), .ZN(n372) );
  XOR2_X1 U473 ( .A(n645), .B(KEYINPUT62), .Z(n373) );
  INV_X1 U474 ( .A(KEYINPUT34), .ZN(n406) );
  XNOR2_X2 U475 ( .A(n388), .B(n411), .ZN(n413) );
  AND2_X1 U476 ( .A1(n410), .A2(n660), .ZN(n409) );
  NAND2_X1 U477 ( .A1(n691), .A2(G234), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n375), .B(n376), .ZN(n506) );
  XOR2_X1 U479 ( .A(n498), .B(n497), .Z(n375) );
  XNOR2_X1 U480 ( .A(n503), .B(n502), .ZN(n376) );
  NAND2_X1 U481 ( .A1(n413), .A2(n379), .ZN(n377) );
  AND2_X1 U482 ( .A1(n415), .A2(n523), .ZN(n379) );
  XNOR2_X1 U483 ( .A(n531), .B(n530), .ZN(n559) );
  NAND2_X1 U484 ( .A1(n414), .A2(KEYINPUT66), .ZN(n395) );
  NAND2_X1 U485 ( .A1(n414), .A2(n372), .ZN(n393) );
  NAND2_X2 U486 ( .A1(n536), .A2(n486), .ZN(n388) );
  NAND2_X1 U487 ( .A1(n374), .A2(n390), .ZN(n381) );
  NAND2_X1 U488 ( .A1(n374), .A2(n390), .ZN(n700) );
  NAND2_X1 U489 ( .A1(n763), .A2(n636), .ZN(n382) );
  NAND2_X1 U490 ( .A1(n763), .A2(n636), .ZN(n655) );
  AND2_X2 U491 ( .A1(n655), .A2(n644), .ZN(n749) );
  INV_X1 U492 ( .A(n423), .ZN(n384) );
  BUF_X2 U493 ( .A(G953), .Z(n385) );
  NAND2_X1 U494 ( .A1(n413), .A2(n415), .ZN(n394) );
  NOR2_X2 U495 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U496 ( .A1(n592), .A2(n593), .ZN(n416) );
  XNOR2_X1 U497 ( .A(n386), .B(n492), .ZN(n493) );
  XNOR2_X1 U498 ( .A(n771), .B(n387), .ZN(n386) );
  INV_X1 U499 ( .A(n491), .ZN(n387) );
  XNOR2_X2 U500 ( .A(G146), .B(G125), .ZN(n472) );
  NAND2_X1 U501 ( .A1(n639), .A2(n648), .ZN(n643) );
  XNOR2_X2 U502 ( .A(n566), .B(KEYINPUT45), .ZN(n648) );
  XNOR2_X2 U503 ( .A(n397), .B(n457), .ZN(n536) );
  NAND2_X1 U504 ( .A1(n581), .A2(n456), .ZN(n397) );
  XNOR2_X2 U505 ( .A(n461), .B(n398), .ZN(n488) );
  XNOR2_X2 U506 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n398) );
  XNOR2_X2 U507 ( .A(G143), .B(G128), .ZN(n461) );
  NAND2_X1 U508 ( .A1(n401), .A2(n400), .ZN(n539) );
  NAND2_X1 U509 ( .A1(n370), .A2(n687), .ZN(n400) );
  NOR2_X1 U510 ( .A1(n687), .A2(n406), .ZN(n403) );
  INV_X1 U511 ( .A(n537), .ZN(n405) );
  NAND2_X2 U512 ( .A1(n408), .A2(n407), .ZN(n607) );
  NAND2_X1 U513 ( .A1(n423), .A2(n422), .ZN(n407) );
  AND2_X2 U514 ( .A1(n425), .A2(n371), .ZN(n408) );
  OR2_X1 U515 ( .A1(n414), .A2(n626), .ZN(n412) );
  NAND2_X1 U516 ( .A1(n369), .A2(n380), .ZN(n529) );
  AND2_X1 U517 ( .A1(n426), .A2(n508), .ZN(n415) );
  NAND2_X1 U518 ( .A1(n594), .A2(n416), .ZN(n595) );
  NAND2_X1 U519 ( .A1(n623), .A2(n718), .ZN(n418) );
  XNOR2_X2 U520 ( .A(n419), .B(KEYINPUT39), .ZN(n623) );
  INV_X1 U521 ( .A(n596), .ZN(n423) );
  NAND2_X1 U522 ( .A1(n596), .A2(KEYINPUT88), .ZN(n425) );
  AND2_X1 U523 ( .A1(n382), .A2(n656), .ZN(n694) );
  OR2_X1 U524 ( .A1(n648), .A2(KEYINPUT2), .ZN(n652) );
  XNOR2_X2 U525 ( .A(n438), .B(G104), .ZN(n478) );
  XNOR2_X2 U526 ( .A(G122), .B(G113), .ZN(n438) );
  XOR2_X1 U527 ( .A(n689), .B(KEYINPUT118), .Z(n427) );
  NOR2_X1 U528 ( .A1(n694), .A2(n693), .ZN(n428) );
  XNOR2_X1 U529 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n618) );
  XNOR2_X1 U530 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n517), .B(n516), .ZN(n750) );
  INV_X1 U532 ( .A(n754), .ZN(n647) );
  INV_X1 U533 ( .A(KEYINPUT119), .ZN(n695) );
  XNOR2_X1 U534 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X2 U535 ( .A(KEYINPUT67), .B(G101), .ZN(n503) );
  XNOR2_X1 U536 ( .A(KEYINPUT70), .B(G110), .ZN(n432) );
  XNOR2_X1 U537 ( .A(n503), .B(n432), .ZN(n491) );
  XNOR2_X1 U538 ( .A(n433), .B(n491), .ZN(n437) );
  XNOR2_X1 U539 ( .A(KEYINPUT18), .B(KEYINPUT90), .ZN(n434) );
  XNOR2_X1 U540 ( .A(n472), .B(n434), .ZN(n435) );
  XNOR2_X1 U541 ( .A(n488), .B(n435), .ZN(n436) );
  XNOR2_X1 U542 ( .A(n437), .B(n436), .ZN(n442) );
  XNOR2_X1 U543 ( .A(n439), .B(G107), .ZN(n462) );
  XNOR2_X1 U544 ( .A(n478), .B(n462), .ZN(n441) );
  XNOR2_X1 U545 ( .A(n501), .B(KEYINPUT16), .ZN(n440) );
  XNOR2_X1 U546 ( .A(n441), .B(n440), .ZN(n757) );
  XNOR2_X1 U547 ( .A(n442), .B(n757), .ZN(n732) );
  NAND2_X1 U548 ( .A1(n732), .A2(n640), .ZN(n445) );
  INV_X1 U549 ( .A(G902), .ZN(n518) );
  NAND2_X1 U550 ( .A1(n518), .A2(n443), .ZN(n446) );
  NAND2_X1 U551 ( .A1(n446), .A2(G210), .ZN(n444) );
  XNOR2_X2 U552 ( .A(n445), .B(n444), .ZN(n596) );
  NAND2_X1 U553 ( .A1(n446), .A2(G214), .ZN(n448) );
  INV_X1 U554 ( .A(KEYINPUT92), .ZN(n447) );
  XNOR2_X1 U555 ( .A(n448), .B(n447), .ZN(n674) );
  INV_X1 U556 ( .A(n674), .ZN(n449) );
  XNOR2_X1 U557 ( .A(n450), .B(KEYINPUT14), .ZN(n451) );
  NAND2_X1 U558 ( .A1(n451), .A2(G952), .ZN(n686) );
  NOR2_X1 U559 ( .A1(n385), .A2(n686), .ZN(n571) );
  NAND2_X1 U560 ( .A1(n451), .A2(G902), .ZN(n568) );
  NOR2_X1 U561 ( .A1(G898), .A2(n691), .ZN(n453) );
  XNOR2_X1 U562 ( .A(KEYINPUT93), .B(n453), .ZN(n759) );
  NOR2_X1 U563 ( .A1(n568), .A2(n759), .ZN(n454) );
  OR2_X1 U564 ( .A1(n571), .A2(n454), .ZN(n455) );
  XNOR2_X1 U565 ( .A(n455), .B(KEYINPUT94), .ZN(n456) );
  INV_X1 U566 ( .A(KEYINPUT0), .ZN(n457) );
  NAND2_X1 U567 ( .A1(G217), .A2(n510), .ZN(n460) );
  XOR2_X1 U568 ( .A(G122), .B(KEYINPUT9), .Z(n458) );
  XNOR2_X1 U569 ( .A(n458), .B(G134), .ZN(n459) );
  XNOR2_X1 U570 ( .A(n460), .B(n459), .ZN(n466) );
  XNOR2_X1 U571 ( .A(n462), .B(n461), .ZN(n464) );
  XNOR2_X1 U572 ( .A(KEYINPUT7), .B(KEYINPUT98), .ZN(n463) );
  NOR2_X1 U573 ( .A1(G902), .A2(n745), .ZN(n470) );
  XNOR2_X1 U574 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n468) );
  INV_X1 U575 ( .A(G478), .ZN(n467) );
  NAND2_X1 U576 ( .A1(n499), .A2(G214), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n472), .B(KEYINPUT10), .ZN(n769) );
  XNOR2_X1 U578 ( .A(n473), .B(n769), .ZN(n480) );
  XNOR2_X1 U579 ( .A(G140), .B(KEYINPUT11), .ZN(n476) );
  XNOR2_X1 U580 ( .A(KEYINPUT12), .B(n474), .ZN(n475) );
  XNOR2_X1 U581 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U582 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U583 ( .A(n480), .B(n479), .ZN(n701) );
  NAND2_X1 U584 ( .A1(n701), .A2(n518), .ZN(n482) );
  XNOR2_X1 U585 ( .A(KEYINPUT13), .B(G475), .ZN(n481) );
  XNOR2_X1 U586 ( .A(n482), .B(n481), .ZN(n546) );
  AND2_X1 U587 ( .A1(n548), .A2(n546), .ZN(n677) );
  NAND2_X1 U588 ( .A1(G234), .A2(n640), .ZN(n483) );
  XNOR2_X1 U589 ( .A(KEYINPUT20), .B(n483), .ZN(n519) );
  NAND2_X1 U590 ( .A1(G221), .A2(n519), .ZN(n484) );
  XNOR2_X1 U591 ( .A(n484), .B(KEYINPUT21), .ZN(n661) );
  XNOR2_X1 U592 ( .A(n661), .B(KEYINPUT96), .ZN(n534) );
  INV_X1 U593 ( .A(n534), .ZN(n485) );
  AND2_X1 U594 ( .A1(n677), .A2(n485), .ZN(n486) );
  XNOR2_X1 U595 ( .A(KEYINPUT69), .B(G469), .ZN(n495) );
  XOR2_X2 U596 ( .A(G137), .B(G140), .Z(n509) );
  XNOR2_X1 U597 ( .A(n509), .B(KEYINPUT95), .ZN(n771) );
  XNOR2_X1 U598 ( .A(n490), .B(n489), .ZN(n492) );
  NOR2_X1 U599 ( .A1(G902), .A2(n741), .ZN(n494) );
  INV_X1 U600 ( .A(KEYINPUT1), .ZN(n496) );
  XNOR2_X1 U601 ( .A(G137), .B(KEYINPUT5), .ZN(n497) );
  NAND2_X1 U602 ( .A1(n499), .A2(G210), .ZN(n500) );
  XNOR2_X1 U603 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U604 ( .A(n504), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n506), .B(n505), .ZN(n645) );
  NOR2_X1 U606 ( .A1(n645), .A2(G902), .ZN(n507) );
  XNOR2_X2 U607 ( .A(n507), .B(G472), .ZN(n589) );
  XOR2_X1 U608 ( .A(G119), .B(n509), .Z(n512) );
  NAND2_X1 U609 ( .A1(G221), .A2(n510), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n512), .B(n511), .ZN(n517) );
  XOR2_X1 U611 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n514) );
  XNOR2_X1 U612 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U613 ( .A(n769), .B(n515), .ZN(n516) );
  NAND2_X1 U614 ( .A1(n750), .A2(n518), .ZN(n522) );
  NAND2_X1 U615 ( .A1(G217), .A2(n519), .ZN(n520) );
  XNOR2_X1 U616 ( .A(n520), .B(KEYINPUT25), .ZN(n521) );
  XNOR2_X2 U617 ( .A(n522), .B(n521), .ZN(n660) );
  INV_X1 U618 ( .A(n660), .ZN(n573) );
  NOR2_X1 U619 ( .A1(n658), .A2(n573), .ZN(n524) );
  XNOR2_X1 U620 ( .A(n524), .B(KEYINPUT102), .ZN(n526) );
  XNOR2_X1 U621 ( .A(n589), .B(KEYINPUT6), .ZN(n605) );
  INV_X1 U622 ( .A(n605), .ZN(n525) );
  INV_X1 U623 ( .A(KEYINPUT77), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n527), .B(KEYINPUT32), .ZN(n528) );
  NAND2_X1 U625 ( .A1(n700), .A2(n698), .ZN(n531) );
  INV_X1 U626 ( .A(KEYINPUT87), .ZN(n530) );
  NAND2_X1 U627 ( .A1(n559), .A2(KEYINPUT44), .ZN(n533) );
  INV_X1 U628 ( .A(KEYINPUT65), .ZN(n532) );
  XNOR2_X1 U629 ( .A(n533), .B(n532), .ZN(n557) );
  NOR2_X1 U630 ( .A1(n534), .A2(n660), .ZN(n544) );
  INV_X1 U631 ( .A(n544), .ZN(n657) );
  NOR2_X1 U632 ( .A1(n658), .A2(n657), .ZN(n540) );
  NAND2_X1 U633 ( .A1(n540), .A2(n605), .ZN(n535) );
  BUF_X1 U634 ( .A(n536), .Z(n537) );
  NOR2_X1 U635 ( .A1(n548), .A2(n546), .ZN(n597) );
  INV_X1 U636 ( .A(KEYINPUT35), .ZN(n538) );
  INV_X1 U637 ( .A(KEYINPUT44), .ZN(n561) );
  INV_X1 U638 ( .A(n589), .ZN(n664) );
  NAND2_X1 U639 ( .A1(n540), .A2(n664), .ZN(n667) );
  INV_X1 U640 ( .A(n667), .ZN(n541) );
  NAND2_X1 U641 ( .A1(n541), .A2(n537), .ZN(n543) );
  INV_X1 U642 ( .A(KEYINPUT31), .ZN(n542) );
  XNOR2_X1 U643 ( .A(n543), .B(n542), .ZN(n723) );
  NOR2_X1 U644 ( .A1(n592), .A2(n664), .ZN(n545) );
  NAND2_X1 U645 ( .A1(n537), .A2(n545), .ZN(n709) );
  NAND2_X1 U646 ( .A1(n723), .A2(n709), .ZN(n550) );
  INV_X1 U647 ( .A(n546), .ZN(n547) );
  NAND2_X1 U648 ( .A1(n550), .A2(n672), .ZN(n553) );
  NOR2_X1 U649 ( .A1(n605), .A2(n660), .ZN(n552) );
  NAND2_X1 U650 ( .A1(n551), .A2(n552), .ZN(n697) );
  AND2_X1 U651 ( .A1(n553), .A2(n697), .ZN(n554) );
  NAND2_X1 U652 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U653 ( .A(n558), .B(KEYINPUT85), .ZN(n565) );
  BUF_X1 U654 ( .A(n559), .Z(n560) );
  XNOR2_X1 U655 ( .A(n560), .B(KEYINPUT86), .ZN(n563) );
  NAND2_X1 U656 ( .A1(n782), .A2(n561), .ZN(n562) );
  OR2_X1 U657 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n565), .A2(n564), .ZN(n566) );
  BUF_X2 U659 ( .A(n648), .Z(n763) );
  INV_X1 U660 ( .A(n567), .ZN(n579) );
  OR2_X1 U661 ( .A1(n691), .A2(n568), .ZN(n569) );
  NOR2_X1 U662 ( .A1(G900), .A2(n569), .ZN(n570) );
  NOR2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U664 ( .A(KEYINPUT78), .B(n572), .ZN(n593) );
  INV_X1 U665 ( .A(n593), .ZN(n575) );
  NAND2_X1 U666 ( .A1(n575), .A2(n574), .ZN(n604) );
  XNOR2_X1 U667 ( .A(KEYINPUT28), .B(KEYINPUT107), .ZN(n576) );
  XNOR2_X1 U668 ( .A(n577), .B(n576), .ZN(n578) );
  NOR2_X1 U669 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U670 ( .A(n580), .B(KEYINPUT108), .ZN(n616) );
  BUF_X1 U671 ( .A(n581), .Z(n582) );
  NAND2_X1 U672 ( .A1(n616), .A2(n582), .ZN(n586) );
  INV_X1 U673 ( .A(n586), .ZN(n719) );
  NAND2_X1 U674 ( .A1(n719), .A2(n672), .ZN(n583) );
  NAND2_X1 U675 ( .A1(n583), .A2(KEYINPUT47), .ZN(n602) );
  INV_X1 U676 ( .A(n672), .ZN(n584) );
  NOR2_X1 U677 ( .A1(n584), .A2(KEYINPUT47), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n585), .B(KEYINPUT73), .ZN(n587) );
  XNOR2_X1 U679 ( .A(n588), .B(KEYINPUT72), .ZN(n600) );
  XNOR2_X1 U680 ( .A(KEYINPUT30), .B(KEYINPUT106), .ZN(n590) );
  XNOR2_X1 U681 ( .A(n591), .B(n590), .ZN(n594) );
  XNOR2_X1 U682 ( .A(KEYINPUT76), .B(n595), .ZN(n613) );
  INV_X1 U683 ( .A(n384), .ZN(n630) );
  NAND2_X1 U684 ( .A1(n597), .A2(n630), .ZN(n598) );
  NOR2_X1 U685 ( .A1(n613), .A2(n598), .ZN(n717) );
  XOR2_X1 U686 ( .A(KEYINPUT81), .B(n717), .Z(n599) );
  NOR2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U689 ( .A(n603), .B(KEYINPUT71), .ZN(n611) );
  INV_X1 U690 ( .A(n718), .ZN(n721) );
  NOR2_X1 U691 ( .A1(n721), .A2(n604), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n606), .A2(n605), .ZN(n625) );
  BUF_X1 U693 ( .A(n607), .Z(n608) );
  NOR2_X1 U694 ( .A1(n625), .A2(n608), .ZN(n609) );
  XNOR2_X1 U695 ( .A(n609), .B(KEYINPUT36), .ZN(n610) );
  INV_X1 U696 ( .A(n658), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n610), .A2(n626), .ZN(n729) );
  NAND2_X1 U698 ( .A1(n611), .A2(n729), .ZN(n621) );
  XOR2_X1 U699 ( .A(KEYINPUT38), .B(KEYINPUT74), .Z(n612) );
  XNOR2_X1 U700 ( .A(n384), .B(n612), .ZN(n675) );
  XOR2_X1 U701 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n615) );
  NOR2_X1 U702 ( .A1(n675), .A2(n674), .ZN(n673) );
  NAND2_X1 U703 ( .A1(n677), .A2(n673), .ZN(n614) );
  XNOR2_X1 U704 ( .A(n615), .B(n614), .ZN(n688) );
  NAND2_X1 U705 ( .A1(n616), .A2(n688), .ZN(n617) );
  XNOR2_X1 U706 ( .A(n617), .B(KEYINPUT42), .ZN(n783) );
  NAND2_X1 U707 ( .A1(n785), .A2(n783), .ZN(n619) );
  XNOR2_X1 U708 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U709 ( .A(n622), .B(KEYINPUT48), .ZN(n638) );
  INV_X1 U710 ( .A(n638), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n623), .A2(n714), .ZN(n731) );
  NAND2_X1 U712 ( .A1(n731), .A2(KEYINPUT2), .ZN(n624) );
  XNOR2_X1 U713 ( .A(n624), .B(KEYINPUT79), .ZN(n633) );
  OR2_X1 U714 ( .A1(n674), .A2(n625), .ZN(n627) );
  NOR2_X1 U715 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U716 ( .A(n628), .B(KEYINPUT104), .ZN(n629) );
  XNOR2_X1 U717 ( .A(KEYINPUT43), .B(n629), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U719 ( .A(n632), .B(KEYINPUT105), .ZN(n781) );
  NAND2_X1 U720 ( .A1(n633), .A2(n781), .ZN(n634) );
  NOR2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n636) );
  AND2_X1 U722 ( .A1(n781), .A2(n731), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n773) );
  NOR2_X1 U724 ( .A1(n773), .A2(n640), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n640), .B(KEYINPUT83), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n641), .A2(KEYINPUT2), .ZN(n642) );
  INV_X1 U727 ( .A(G952), .ZN(n646) );
  AND2_X1 U728 ( .A1(n646), .A2(n385), .ZN(n754) );
  INV_X1 U729 ( .A(KEYINPUT2), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n773), .A2(n649), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(KEYINPUT82), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n654), .B(n653), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(KEYINPUT50), .ZN(n666) );
  AND2_X1 U736 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U737 ( .A(KEYINPUT49), .B(n662), .Z(n663) );
  NOR2_X1 U738 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n670) );
  XOR2_X1 U741 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n669) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n671), .A2(n688), .ZN(n683) );
  NAND2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n679) );
  NAND2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U748 ( .A(KEYINPUT117), .B(n680), .Z(n681) );
  NAND2_X1 U749 ( .A1(n681), .A2(n687), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U751 ( .A(KEYINPUT52), .B(n684), .Z(n685) );
  NOR2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U754 ( .A(n695), .B(KEYINPUT53), .ZN(n696) );
  XNOR2_X1 U755 ( .A(n428), .B(n696), .ZN(G75) );
  XNOR2_X1 U756 ( .A(n697), .B(G101), .ZN(G3) );
  XOR2_X1 U757 ( .A(G119), .B(KEYINPUT126), .Z(n699) );
  XOR2_X1 U758 ( .A(n699), .B(n698), .Z(G21) );
  XNOR2_X1 U759 ( .A(n381), .B(G110), .ZN(G12) );
  NAND2_X1 U760 ( .A1(n749), .A2(G475), .ZN(n703) );
  XNOR2_X1 U761 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X2 U762 ( .A1(n704), .A2(n754), .ZN(n706) );
  XNOR2_X1 U763 ( .A(KEYINPUT120), .B(KEYINPUT60), .ZN(n705) );
  XNOR2_X1 U764 ( .A(n706), .B(n705), .ZN(G60) );
  NOR2_X1 U765 ( .A1(n721), .A2(n709), .ZN(n707) );
  XOR2_X1 U766 ( .A(KEYINPUT110), .B(n707), .Z(n708) );
  XNOR2_X1 U767 ( .A(G104), .B(n708), .ZN(G6) );
  INV_X1 U768 ( .A(n714), .ZN(n724) );
  NOR2_X1 U769 ( .A1(n709), .A2(n724), .ZN(n713) );
  XOR2_X1 U770 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n711) );
  XNOR2_X1 U771 ( .A(G107), .B(KEYINPUT111), .ZN(n710) );
  XNOR2_X1 U772 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U773 ( .A(n713), .B(n712), .ZN(G9) );
  XOR2_X1 U774 ( .A(n396), .B(KEYINPUT29), .Z(n716) );
  NAND2_X1 U775 ( .A1(n719), .A2(n714), .ZN(n715) );
  XNOR2_X1 U776 ( .A(n716), .B(n715), .ZN(G30) );
  XOR2_X1 U777 ( .A(G143), .B(n717), .Z(G45) );
  NAND2_X1 U778 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n720), .B(G146), .ZN(G48) );
  NOR2_X1 U780 ( .A1(n721), .A2(n723), .ZN(n722) );
  XOR2_X1 U781 ( .A(G113), .B(n722), .Z(G15) );
  NOR2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n726) );
  XNOR2_X1 U783 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n725) );
  XNOR2_X1 U784 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U785 ( .A(G116), .B(n727), .ZN(G18) );
  XOR2_X1 U786 ( .A(KEYINPUT37), .B(KEYINPUT114), .Z(n728) );
  XNOR2_X1 U787 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U788 ( .A(G125), .B(n730), .ZN(G27) );
  XNOR2_X1 U789 ( .A(G134), .B(n731), .ZN(G36) );
  NAND2_X1 U790 ( .A1(n749), .A2(G210), .ZN(n736) );
  BUF_X1 U791 ( .A(n732), .Z(n733) );
  XOR2_X1 U792 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n734) );
  XNOR2_X1 U793 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X2 U794 ( .A1(n737), .A2(n754), .ZN(n739) );
  XNOR2_X1 U795 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n738) );
  XNOR2_X1 U796 ( .A(n739), .B(n738), .ZN(G51) );
  NAND2_X1 U797 ( .A1(n383), .A2(G469), .ZN(n743) );
  XOR2_X1 U798 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n740) );
  NOR2_X1 U799 ( .A1(n754), .A2(n744), .ZN(G54) );
  NAND2_X1 U800 ( .A1(n383), .A2(G478), .ZN(n747) );
  XOR2_X1 U801 ( .A(n745), .B(KEYINPUT121), .Z(n746) );
  XNOR2_X1 U802 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U803 ( .A1(n754), .A2(n748), .ZN(G63) );
  NAND2_X1 U804 ( .A1(n383), .A2(G217), .ZN(n752) );
  XOR2_X1 U805 ( .A(KEYINPUT122), .B(n750), .Z(n751) );
  XNOR2_X1 U806 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U807 ( .A1(n754), .A2(n753), .ZN(G66) );
  XNOR2_X1 U808 ( .A(G101), .B(G110), .ZN(n755) );
  XOR2_X1 U809 ( .A(KEYINPUT125), .B(n755), .Z(n756) );
  XNOR2_X1 U810 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U811 ( .A1(n759), .A2(n758), .ZN(n768) );
  NAND2_X1 U812 ( .A1(n385), .A2(G224), .ZN(n760) );
  XNOR2_X1 U813 ( .A(KEYINPUT61), .B(n760), .ZN(n761) );
  NAND2_X1 U814 ( .A1(n761), .A2(G898), .ZN(n762) );
  XNOR2_X1 U815 ( .A(KEYINPUT123), .B(n762), .ZN(n766) );
  NAND2_X1 U816 ( .A1(n763), .A2(n691), .ZN(n764) );
  XOR2_X1 U817 ( .A(KEYINPUT124), .B(n764), .Z(n765) );
  NOR2_X1 U818 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(G69) );
  XNOR2_X1 U820 ( .A(n770), .B(n769), .ZN(n772) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(n775) );
  XNOR2_X1 U822 ( .A(n775), .B(n773), .ZN(n774) );
  NAND2_X1 U823 ( .A1(n774), .A2(n691), .ZN(n779) );
  XNOR2_X1 U824 ( .A(G227), .B(n775), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n776), .A2(G900), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n385), .A2(n777), .ZN(n778) );
  NAND2_X1 U827 ( .A1(n779), .A2(n778), .ZN(G72) );
  XOR2_X1 U828 ( .A(G140), .B(KEYINPUT115), .Z(n780) );
  XNOR2_X1 U829 ( .A(n781), .B(n780), .ZN(G42) );
  XNOR2_X1 U830 ( .A(G122), .B(n782), .ZN(G24) );
  XOR2_X1 U831 ( .A(G137), .B(n783), .Z(n784) );
  XNOR2_X1 U832 ( .A(KEYINPUT127), .B(n784), .ZN(G39) );
  XNOR2_X1 U833 ( .A(n785), .B(G131), .ZN(G33) );
endmodule

