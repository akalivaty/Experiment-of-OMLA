//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G68), .Z(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n247), .A2(new_n213), .A3(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT69), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n206), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G68), .ZN(new_n252));
  OR3_X1    g0052(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n249), .B2(new_n252), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n207), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n248), .A2(new_n213), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT11), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n247), .A2(G68), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT12), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n260), .A2(KEYINPUT11), .A3(new_n261), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n255), .A2(new_n264), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT70), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n267), .A2(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(new_n255), .A4(new_n264), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G97), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n284), .A2(new_n286), .A3(G226), .A4(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n278), .A2(KEYINPUT68), .A3(G226), .A4(new_n287), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n277), .B1(new_n282), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT64), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT64), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n296), .B(new_n206), .C1(G41), .C2(G45), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  INV_X1    g0099(.A(new_n213), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n276), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n277), .A2(new_n294), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G238), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT13), .B1(new_n293), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  INV_X1    g0107(.A(new_n305), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(new_n277), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT14), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(G169), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n310), .A3(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n311), .B2(G169), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n275), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n251), .A2(G50), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n249), .A2(new_n318), .B1(G50), .B2(new_n247), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n203), .A2(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n256), .A2(G150), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n320), .B(new_n321), .C1(new_n322), .C2(new_n259), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n323), .B2(new_n261), .ZN(new_n324));
  INV_X1    g0124(.A(new_n277), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n278), .A2(G1698), .ZN(new_n326));
  INV_X1    g0126(.A(G223), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(new_n258), .B2(new_n278), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n278), .A2(G222), .A3(new_n287), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n277), .A2(G274), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n295), .B2(new_n297), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(G226), .B2(new_n303), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(G179), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  AOI211_X1 g0136(.A(new_n324), .B(new_n335), .C1(new_n336), .C2(new_n334), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(G200), .B2(new_n334), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n324), .A2(KEYINPUT9), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT66), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n324), .A2(KEYINPUT9), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n343), .B(KEYINPUT67), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT10), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n340), .A2(new_n347), .A3(new_n342), .A4(new_n344), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n337), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n326), .A2(new_n219), .B1(new_n350), .B2(new_n278), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n284), .A2(new_n286), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n352), .A2(new_n225), .A3(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n325), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n332), .B1(G244), .B2(new_n303), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G200), .ZN(new_n357));
  INV_X1    g0157(.A(new_n261), .ZN(new_n358));
  INV_X1    g0158(.A(new_n322), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n361), .A2(new_n259), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n251), .A2(G77), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n249), .A2(new_n364), .B1(G77), .B2(new_n247), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n357), .B(new_n366), .C1(new_n338), .C2(new_n356), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n356), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(G169), .B1(new_n363), .B2(new_n365), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT65), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n370), .A2(KEYINPUT65), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n368), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n306), .A2(new_n310), .A3(G190), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n274), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n306), .B2(new_n310), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT71), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n382), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n274), .A4(new_n379), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  AND4_X1   g0187(.A1(new_n317), .A2(new_n349), .A3(new_n378), .A4(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n284), .A2(new_n286), .A3(G223), .A4(new_n287), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n283), .B2(new_n220), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n278), .A2(G226), .A3(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n325), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n277), .A2(G232), .A3(new_n294), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT73), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n277), .A2(new_n294), .A3(new_n396), .A4(G232), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n395), .A2(new_n397), .B1(new_n298), .B2(new_n301), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n397), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n400), .A2(KEYINPUT74), .A3(new_n302), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n399), .A2(new_n401), .A3(G179), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n399), .B2(new_n401), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n302), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(KEYINPUT75), .A3(new_n408), .A4(new_n393), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n402), .B1(new_n410), .B2(new_n336), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n359), .A2(new_n251), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n412), .A2(new_n249), .B1(new_n247), .B2(new_n359), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n224), .A2(new_n218), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n414), .B2(new_n201), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n256), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(KEYINPUT72), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT7), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n278), .B2(G20), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n352), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n218), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT72), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n415), .B2(new_n416), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n418), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n358), .B1(new_n425), .B2(KEYINPUT16), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n422), .B2(new_n417), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n413), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n411), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n411), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n389), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(KEYINPUT76), .A2(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(G200), .B1(new_n404), .B2(new_n409), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n399), .A2(new_n401), .A3(G190), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n429), .B(KEYINPUT17), .C1(new_n438), .C2(new_n439), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n388), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n221), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n277), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n206), .A2(G45), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n331), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n219), .A2(new_n287), .ZN(new_n454));
  INV_X1    g0254(.A(G244), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G1698), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n284), .A2(new_n454), .A3(new_n286), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n283), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n277), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(KEYINPUT80), .A3(new_n460), .ZN(new_n464));
  AOI211_X1 g0264(.A(G179), .B(new_n453), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n325), .A3(new_n464), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n301), .A2(new_n449), .B1(new_n450), .B2(new_n277), .ZN(new_n468));
  AOI21_X1  g0268(.A(G169), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n206), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n247), .A2(new_n471), .A3(new_n213), .A4(new_n248), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n361), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n284), .A2(new_n286), .A3(new_n207), .A4(G68), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n226), .A2(KEYINPUT77), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT77), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G97), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n259), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n476), .B1(new_n480), .B2(KEYINPUT19), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G87), .A2(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n207), .B1(new_n280), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n261), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n474), .A2(new_n247), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT81), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT77), .B(G97), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n484), .B1(new_n492), .B2(new_n259), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n483), .A2(new_n485), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(new_n476), .ZN(new_n495));
  AOI211_X1 g0295(.A(new_n491), .B(new_n488), .C1(new_n495), .C2(new_n261), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n475), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n470), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n487), .A2(new_n489), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n491), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n487), .A2(KEYINPUT81), .A3(new_n489), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n472), .A2(new_n220), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G238), .A2(G1698), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n455), .B2(G1698), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n459), .B1(new_n506), .B2(new_n278), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n325), .B1(new_n507), .B2(KEYINPUT80), .ZN(new_n508));
  INV_X1    g0308(.A(new_n464), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n338), .B(new_n468), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n453), .B1(new_n463), .B2(new_n464), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(G200), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n502), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n284), .A2(new_n286), .A3(new_n207), .A4(G87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n278), .A2(new_n516), .A3(new_n207), .A4(G87), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT23), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n207), .B2(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n350), .A2(KEYINPUT23), .A3(G20), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(new_n522), .B1(new_n459), .B2(new_n207), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n518), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n519), .B1(new_n518), .B2(new_n523), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n261), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n247), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(KEYINPUT25), .A3(new_n350), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n247), .B2(G107), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n473), .A2(G107), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n284), .A2(new_n286), .A3(G257), .A4(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n284), .A2(new_n286), .A3(G250), .A4(new_n287), .ZN(new_n533));
  INV_X1    g0333(.A(G294), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n283), .C2(new_n534), .ZN(new_n535));
  OR2_X1    g0335(.A1(KEYINPUT5), .A2(G41), .ZN(new_n536));
  NAND2_X1  g0336(.A1(KEYINPUT5), .A2(G41), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n452), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n325), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n535), .A2(new_n325), .B1(new_n539), .B2(G264), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n301), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(G190), .ZN(new_n543));
  AOI21_X1  g0343(.A(G200), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n526), .B(new_n531), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n498), .A2(new_n513), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n284), .A2(new_n286), .A3(G244), .A4(new_n287), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n287), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n549), .A2(new_n550), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n325), .ZN(new_n554));
  AND2_X1   g0354(.A1(KEYINPUT5), .A2(G41), .ZN(new_n555));
  NOR2_X1   g0355(.A1(KEYINPUT5), .A2(G41), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n449), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n277), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n541), .B1(new_n558), .B2(new_n227), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(KEYINPUT79), .A3(G200), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT79), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n559), .B1(new_n553), .B2(new_n325), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(new_n381), .ZN(new_n565));
  AND2_X1   g0365(.A1(G97), .A2(G107), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G97), .A2(G107), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n350), .A2(KEYINPUT6), .ZN(new_n569));
  OAI22_X1  g0369(.A1(new_n568), .A2(KEYINPUT6), .B1(new_n492), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n278), .A2(new_n419), .A3(G20), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT7), .B1(new_n352), .B2(new_n207), .ZN(new_n573));
  OAI21_X1  g0373(.A(G107), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n358), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n472), .A2(G97), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n247), .A2(new_n226), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n564), .A2(G190), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n562), .A2(new_n565), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n564), .A2(new_n372), .ZN(new_n585));
  OAI221_X1 g0385(.A(new_n585), .B1(G169), .B2(new_n564), .C1(new_n575), .C2(new_n581), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n546), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n247), .A2(G116), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n473), .B2(G116), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n207), .B(new_n551), .C1(new_n492), .C2(G33), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n248), .A2(new_n213), .B1(G20), .B2(new_n458), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT20), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(G33), .B1(new_n477), .B2(new_n479), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n551), .A2(new_n207), .ZN(new_n595));
  OAI211_X1 g0395(.A(KEYINPUT20), .B(new_n592), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n590), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n284), .A2(new_n286), .A3(G264), .A4(G1698), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n284), .A2(new_n286), .A3(G257), .A4(new_n287), .ZN(new_n600));
  XNOR2_X1  g0400(.A(KEYINPUT82), .B(G303), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n599), .B(new_n600), .C1(new_n278), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n325), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n539), .A2(G270), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n603), .A2(new_n541), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n598), .B1(new_n605), .B2(G190), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n381), .B2(new_n605), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n540), .A2(new_n372), .A3(new_n541), .ZN(new_n608));
  AOI21_X1  g0408(.A(G169), .B1(new_n540), .B2(new_n541), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n526), .A2(new_n531), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n605), .A2(new_n598), .A3(G179), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n603), .A2(new_n541), .A3(new_n604), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n598), .A2(new_n614), .A3(KEYINPUT21), .A4(G169), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n598), .A2(new_n614), .A3(G169), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n607), .A2(new_n612), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n447), .A2(new_n588), .A3(new_n620), .ZN(G372));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n588), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n612), .A2(new_n616), .A3(new_n619), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT83), .B1(new_n546), .B2(new_n587), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n498), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n498), .A2(new_n513), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n586), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n503), .B1(new_n500), .B2(new_n501), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n512), .B1(new_n470), .B2(new_n497), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n575), .A2(new_n581), .B1(new_n564), .B2(G169), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n561), .A2(G179), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(KEYINPUT26), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n627), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n626), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n447), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n434), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n433), .B1(new_n411), .B2(new_n430), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n317), .ZN(new_n643));
  INV_X1    g0443(.A(new_n380), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n384), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n374), .A2(new_n376), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n442), .A2(new_n443), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n642), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n346), .A2(new_n348), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n337), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n639), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT84), .Z(G369));
  INV_X1    g0454(.A(G13), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n655), .A2(G1), .A3(G20), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n598), .A2(new_n616), .A3(new_n619), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n598), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n616), .A2(new_n607), .A3(new_n619), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n545), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n611), .A2(new_n662), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n612), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n662), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n610), .A3(new_n611), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n662), .B1(new_n616), .B2(new_n619), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n670), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT86), .Z(G399));
  INV_X1    g0479(.A(new_n210), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n483), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n216), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n511), .A2(new_n540), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n614), .A2(new_n372), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n564), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n687), .A2(KEYINPUT30), .A3(new_n564), .A4(new_n688), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n605), .A2(new_n511), .A3(G179), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n561), .A3(new_n542), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(new_n662), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n588), .A2(new_n620), .A3(new_n671), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(KEYINPUT31), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(G330), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n662), .B1(new_n626), .B2(new_n637), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n498), .A2(new_n513), .A3(new_n545), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n584), .A2(new_n586), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(new_n624), .ZN(new_n707));
  AOI211_X1 g0507(.A(KEYINPUT87), .B(new_n662), .C1(new_n637), .C2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT87), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT26), .B1(new_n632), .B2(new_n635), .ZN(new_n710));
  AND4_X1   g0510(.A1(KEYINPUT26), .A2(new_n498), .A3(new_n513), .A4(new_n635), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n707), .B(new_n498), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n709), .B1(new_n712), .B2(new_n671), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT29), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n702), .B1(new_n704), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n686), .B1(new_n715), .B2(G1), .ZN(G364));
  NOR2_X1   g0516(.A1(new_n666), .A2(G330), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT88), .Z(new_n718));
  NOR2_X1   g0518(.A1(new_n655), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n206), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n681), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n667), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n381), .A2(G179), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(G20), .A3(G190), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n207), .A2(new_n372), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G190), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n278), .B1(new_n220), .B2(new_n726), .C1(new_n730), .C2(new_n218), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n728), .A2(new_n338), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(G50), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n338), .A2(G20), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n725), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G107), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n372), .A2(new_n381), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT92), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n735), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G159), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT32), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n727), .A2(KEYINPUT90), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(G190), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G58), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n733), .A2(new_n738), .A3(new_n744), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n740), .A2(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G97), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n746), .A2(new_n338), .A3(new_n747), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n754), .B1(new_n258), .B2(new_n755), .C1(new_n743), .C2(KEYINPUT32), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G329), .A2(new_n742), .B1(new_n737), .B2(G283), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n352), .B1(new_n726), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n759), .B1(G326), .B2(new_n732), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  OAI211_X1 g0561(.A(new_n757), .B(new_n760), .C1(new_n730), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n755), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G311), .A2(new_n763), .B1(new_n749), .B2(G322), .ZN(new_n764));
  INV_X1    g0564(.A(new_n753), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n534), .B2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n751), .A2(new_n756), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n213), .B1(G20), .B2(new_n336), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n210), .A2(G355), .A3(new_n278), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n680), .A2(new_n278), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G45), .B2(new_n216), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n245), .A2(new_n448), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n770), .B1(G116), .B2(new_n210), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n207), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT89), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n768), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n723), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n769), .B(new_n780), .C1(new_n666), .C2(new_n777), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n724), .A2(new_n781), .ZN(G396));
  NAND3_X1  g0582(.A1(new_n377), .A2(new_n373), .A3(new_n371), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n783), .B(new_n367), .C1(new_n366), .C2(new_n671), .ZN(new_n784));
  INV_X1    g0584(.A(new_n366), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n646), .A2(new_n785), .A3(new_n662), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n703), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n703), .A2(new_n787), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n702), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT95), .Z(new_n792));
  OAI211_X1 g0592(.A(new_n792), .B(new_n723), .C1(new_n702), .C2(new_n790), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n768), .A2(new_n775), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n722), .B1(G77), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n732), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n352), .B1(new_n350), .B2(new_n726), .C1(new_n797), .C2(new_n758), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n737), .A2(G87), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(G311), .C2(new_n742), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n755), .A2(new_n458), .B1(new_n802), .B2(new_n730), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT93), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n749), .A2(G294), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n801), .A2(new_n804), .A3(new_n754), .A4(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n729), .A2(G150), .B1(new_n732), .B2(G137), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n755), .B2(new_n808), .C1(new_n809), .C2(new_n748), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n278), .B1(new_n741), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT94), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n753), .A2(G58), .ZN(new_n817));
  INV_X1    g0617(.A(new_n726), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n737), .A2(G68), .B1(G50), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n806), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n796), .B1(new_n821), .B2(new_n768), .ZN(new_n822));
  INV_X1    g0622(.A(new_n775), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n787), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n793), .A2(new_n824), .ZN(G384));
  AOI211_X1 g0625(.A(new_n458), .B(new_n215), .C1(new_n570), .C2(KEYINPUT35), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(KEYINPUT35), .B2(new_n570), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT36), .Z(new_n828));
  NOR3_X1   g0628(.A1(new_n414), .A2(new_n216), .A3(new_n258), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT96), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n829), .A2(new_n830), .B1(new_n202), .B2(G68), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n206), .B(G13), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n426), .B1(KEYINPUT16), .B2(new_n425), .ZN(new_n835));
  INV_X1    g0635(.A(new_n413), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n660), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n435), .B2(new_n444), .ZN(new_n838));
  AOI21_X1  g0638(.A(G169), .B1(new_n404), .B2(new_n409), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n660), .B1(new_n839), .B2(new_n402), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n835), .A2(new_n836), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n440), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n844));
  INV_X1    g0644(.A(new_n440), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n840), .A2(new_n430), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n838), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n317), .A2(KEYINPUT97), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT97), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n275), .C1(new_n315), .C2(new_n316), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n274), .A2(new_n671), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n644), .B2(new_n384), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n315), .A2(new_n316), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n387), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n858), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n783), .A2(new_n662), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n789), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n854), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n642), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n660), .ZN(new_n870));
  INV_X1    g0670(.A(new_n848), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n440), .A2(KEYINPUT98), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT98), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n429), .B(new_n873), .C1(new_n438), .C2(new_n439), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n847), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(KEYINPUT99), .A3(KEYINPUT37), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n429), .B(new_n660), .C1(new_n642), .C2(new_n648), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n851), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n853), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n882), .A2(new_n884), .B1(new_n854), .B2(KEYINPUT39), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n855), .A2(new_n857), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n671), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n868), .B(new_n870), .C1(new_n885), .C2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n704), .A2(new_n714), .A3(new_n447), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n652), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n888), .B(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(G330), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n699), .A2(KEYINPUT100), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT100), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n695), .A2(new_n894), .A3(KEYINPUT31), .A4(new_n662), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n787), .B1(new_n698), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n864), .ZN(new_n898));
  INV_X1    g0698(.A(new_n853), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n838), .B2(new_n849), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n897), .A2(new_n864), .A3(new_n902), .ZN(new_n904));
  INV_X1    g0704(.A(new_n879), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT99), .B1(new_n875), .B2(KEYINPUT37), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n848), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n429), .A2(new_n660), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n649), .B2(new_n869), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n904), .B1(new_n910), .B2(new_n899), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n388), .B(new_n445), .C1(new_n698), .C2(new_n896), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n892), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n891), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n206), .B2(new_n719), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n891), .A2(new_n915), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n834), .B1(new_n917), .B2(new_n918), .ZN(G367));
  NOR2_X1   g0719(.A1(new_n671), .A2(new_n631), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n627), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n629), .B2(new_n920), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n706), .B1(new_n582), .B2(new_n671), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n635), .A2(new_n662), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT42), .B1(new_n926), .B2(new_n676), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n586), .B1(new_n924), .B2(new_n612), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n671), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n926), .A2(KEYINPUT42), .A3(new_n676), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT101), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n674), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n926), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n933), .A2(new_n935), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n940), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n942), .A2(new_n936), .B1(new_n938), .B2(new_n926), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n681), .B(KEYINPUT41), .Z(new_n944));
  XNOR2_X1  g0744(.A(new_n673), .B(new_n675), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n667), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n715), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n926), .A2(new_n677), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT44), .Z(new_n949));
  NOR2_X1   g0749(.A1(new_n926), .A2(new_n677), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT45), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n949), .A2(new_n938), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n938), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  OR3_X1    g0753(.A1(new_n947), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n944), .B1(new_n954), .B2(new_n715), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n941), .B(new_n943), .C1(new_n955), .C2(new_n721), .ZN(new_n956));
  INV_X1    g0756(.A(new_n771), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n238), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n779), .B1(new_n210), .B2(new_n361), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT46), .B1(new_n818), .B2(G116), .ZN(new_n960));
  INV_X1    g0760(.A(G311), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n730), .A2(new_n534), .B1(new_n797), .B2(new_n961), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(G283), .C2(new_n763), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n818), .A2(KEYINPUT46), .A3(G116), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n352), .B(new_n964), .C1(new_n736), .C2(new_n492), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G317), .B2(new_n742), .ZN(new_n966));
  INV_X1    g0766(.A(new_n601), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n967), .A2(new_n749), .B1(new_n753), .B2(G107), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n963), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n749), .A2(G150), .B1(G143), .B2(new_n732), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n218), .B2(new_n765), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT102), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G137), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n741), .A2(new_n974), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n278), .B1(new_n224), .B2(new_n726), .C1(new_n730), .C2(new_n808), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(G77), .C2(new_n737), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n973), .B(new_n977), .C1(new_n202), .C2(new_n755), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n971), .A2(new_n972), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n969), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  INV_X1    g0781(.A(new_n768), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n722), .B1(new_n958), .B2(new_n959), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT103), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(new_n777), .C2(new_n922), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n956), .A2(new_n987), .ZN(G387));
  NOR2_X1   g0788(.A1(new_n235), .A2(new_n448), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n322), .A2(G50), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT50), .ZN(new_n991));
  INV_X1    g0791(.A(new_n683), .ZN(new_n992));
  AOI211_X1 g0792(.A(G45), .B(new_n992), .C1(G68), .C2(G77), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n957), .B(new_n989), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(new_n210), .A3(new_n278), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(G107), .B2(new_n210), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT104), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n779), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n753), .A2(new_n474), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n202), .B2(new_n748), .C1(new_n218), .C2(new_n755), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n352), .B1(new_n818), .B2(G77), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n797), .B2(new_n808), .C1(new_n322), .C2(new_n730), .ZN(new_n1002));
  INV_X1    g0802(.A(G150), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n741), .A2(new_n1003), .B1(new_n736), .B2(new_n226), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT105), .B(G322), .Z(new_n1006));
  AOI22_X1  g0806(.A1(G311), .A2(new_n729), .B1(new_n732), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(new_n755), .B2(new_n601), .C1(new_n1008), .C2(new_n748), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT48), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n753), .A2(G283), .B1(G294), .B2(new_n818), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT49), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n736), .A2(new_n458), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n742), .A2(G326), .ZN(new_n1018));
  NOR4_X1   g0818(.A1(new_n1016), .A2(new_n278), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1005), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n722), .B(new_n998), .C1(new_n1021), .C2(new_n982), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n673), .B2(new_n778), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n946), .B2(new_n721), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n947), .A2(new_n681), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n715), .A2(new_n946), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT106), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(G393));
  AND2_X1   g0831(.A1(new_n954), .A2(new_n681), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n952), .A2(new_n953), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n947), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n720), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n957), .A2(new_n242), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n779), .B1(new_n210), .B2(new_n492), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n755), .A2(new_n322), .B1(new_n202), .B2(new_n730), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n352), .B1(new_n818), .B2(G68), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n799), .B(new_n1040), .C1(new_n809), .C2(new_n741), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT107), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(G77), .C2(new_n753), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n748), .A2(new_n808), .B1(new_n1003), .B2(new_n797), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT51), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n748), .A2(new_n961), .B1(new_n1008), .B2(new_n797), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n278), .B1(new_n818), .B2(G283), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n738), .B(new_n1048), .C1(new_n601), .C2(new_n730), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n765), .A2(new_n458), .B1(new_n534), .B2(new_n755), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n742), .C2(new_n1006), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1043), .A2(new_n1045), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n722), .B1(new_n1037), .B2(new_n1038), .C1(new_n1052), .C2(new_n982), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT108), .Z(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n778), .B2(new_n926), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1036), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1035), .A2(new_n1056), .ZN(G390));
  INV_X1    g0857(.A(KEYINPUT109), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n787), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n498), .B1(new_n710), .B2(new_n711), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n705), .A2(new_n706), .A3(new_n624), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n671), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT87), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n712), .A2(new_n709), .A3(new_n671), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1059), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1058), .B1(new_n1065), .B2(new_n865), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n787), .B1(new_n708), .B2(new_n713), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(KEYINPUT109), .A3(new_n866), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n864), .B(KEYINPUT110), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n887), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n882), .B2(new_n853), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n882), .A2(new_n884), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n1071), .C2(new_n867), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n787), .B(G330), .C1(new_n698), .C2(new_n700), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n860), .A2(new_n863), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1073), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n698), .A2(new_n896), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1082), .A2(G330), .A3(new_n787), .A4(new_n1079), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n721), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n722), .B1(new_n359), .B2(new_n795), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT114), .Z(new_n1088));
  OAI22_X1  g0888(.A1(new_n741), .A2(new_n534), .B1(new_n736), .B2(new_n218), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n352), .B1(new_n220), .B2(new_n726), .C1(new_n730), .C2(new_n350), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G283), .C2(new_n732), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G116), .A2(new_n749), .B1(new_n753), .B2(G77), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n492), .C2(new_n755), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n726), .B2(new_n1003), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n818), .A2(new_n1094), .A3(G150), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n730), .C2(new_n974), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G132), .B2(new_n749), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n737), .A2(G50), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT54), .B(G143), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n763), .A2(new_n1102), .B1(new_n753), .B2(G159), .ZN(new_n1103));
  INV_X1    g0903(.A(G128), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n278), .B1(new_n797), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G125), .B2(new_n742), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .A4(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1093), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1088), .B1(new_n982), .B2(new_n1108), .C1(new_n1109), .C2(new_n823), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1086), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT113), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1077), .A2(new_n864), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1083), .A2(new_n1114), .B1(new_n789), .B2(new_n866), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1079), .B(KEYINPUT110), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1082), .A2(G330), .A3(new_n787), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1117), .A2(new_n1118), .B1(new_n1079), .B2(new_n1078), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1115), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n447), .A2(KEYINPUT111), .A3(new_n1082), .A4(G330), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT111), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n913), .B2(new_n892), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1124), .A2(new_n652), .A3(new_n889), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT112), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n682), .B1(new_n1085), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1115), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1125), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(KEYINPUT112), .B(new_n1132), .C1(new_n1081), .C2(new_n1084), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1113), .B1(new_n1127), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1073), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n867), .A2(new_n1071), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n885), .A2(new_n1136), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1126), .B(new_n1135), .C1(new_n1137), .C2(new_n1083), .ZN(new_n1138));
  AND4_X1   g0938(.A1(new_n1113), .A2(new_n1133), .A3(new_n681), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1112), .B1(new_n1134), .B2(new_n1139), .ZN(G378));
  OAI211_X1 g0940(.A(new_n1135), .B(new_n1130), .C1(new_n1137), .C2(new_n1083), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1131), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n660), .A2(new_n324), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT117), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n349), .B(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1147));
  XOR2_X1   g0947(.A(new_n1146), .B(new_n1147), .Z(new_n1148));
  NAND2_X1  g0948(.A1(new_n882), .A2(new_n853), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1149), .A2(new_n904), .B1(new_n901), .B2(new_n902), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1148), .B1(new_n1150), .B2(G330), .ZN(new_n1151));
  AND4_X1   g0951(.A1(G330), .A2(new_n903), .A3(new_n911), .A4(new_n1148), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n888), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1148), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n912), .B2(new_n892), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(G330), .A3(new_n1148), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n868), .A2(new_n870), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1071), .B2(new_n1109), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1143), .B1(new_n1153), .B2(new_n1159), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1159), .A2(new_n1143), .ZN(new_n1161));
  OAI211_X1 g0961(.A(KEYINPUT57), .B(new_n1142), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1142), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1166), .A3(new_n681), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n721), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n732), .A2(G125), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n729), .A2(G132), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n818), .A2(new_n1102), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n765), .A2(new_n1003), .B1(new_n1104), .B2(new_n748), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G137), .C2(new_n763), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n737), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n742), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n736), .A2(new_n224), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n278), .A2(G41), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(new_n258), .B2(new_n726), .C1(new_n730), .C2(new_n226), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(G283), .C2(new_n742), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n350), .B2(new_n748), .C1(new_n361), .C2(new_n755), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n753), .A2(G68), .B1(G116), .B2(new_n732), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT116), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1179), .A2(new_n1180), .B1(KEYINPUT58), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1182), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n768), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n723), .B1(new_n202), .B2(new_n794), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n1148), .C2(new_n823), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1168), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1167), .A2(new_n1196), .ZN(G375));
  INV_X1    g0997(.A(new_n944), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1132), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n999), .B1(new_n802), .B2(new_n748), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT119), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n741), .A2(new_n758), .B1(new_n736), .B2(new_n258), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n278), .B1(new_n818), .B2(G97), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n797), .B2(new_n534), .C1(new_n458), .C2(new_n730), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G107), .C2(new_n763), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n352), .B1(new_n818), .B2(G159), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n797), .B2(new_n812), .C1(new_n730), .C2(new_n1101), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1181), .B(new_n1208), .C1(G128), .C2(new_n742), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n974), .A2(new_n748), .B1(new_n755), .B2(new_n1003), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G50), .B2(new_n753), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1202), .A2(new_n1206), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n722), .B1(G68), .B2(new_n795), .C1(new_n1212), .C2(new_n982), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1117), .B2(new_n775), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1130), .B2(new_n721), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1200), .A2(new_n1215), .ZN(G381));
  XOR2_X1   g1016(.A(G375), .B(KEYINPUT120), .Z(new_n1217));
  AOI21_X1  g1017(.A(new_n1111), .B1(new_n1133), .B2(new_n1127), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G393), .A2(G396), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1220), .A2(new_n1215), .A3(new_n1200), .A4(new_n1221), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1217), .A2(new_n1219), .A3(new_n1222), .ZN(G407));
  NAND2_X1  g1023(.A1(new_n661), .A2(G213), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1218), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(new_n1217), .C2(new_n1226), .ZN(G409));
  NAND3_X1  g1027(.A1(G390), .A2(new_n956), .A3(new_n987), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT124), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G387), .A2(new_n1035), .A3(new_n1056), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(G390), .A2(KEYINPUT124), .A3(new_n956), .A4(new_n987), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT123), .B1(new_n1234), .B2(new_n1221), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1234), .A2(new_n1221), .A3(KEYINPUT123), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1231), .B(new_n1228), .C1(new_n1221), .C2(new_n1234), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(G378), .A2(new_n1167), .A3(new_n1196), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1142), .A2(new_n1198), .A3(new_n1163), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT121), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n721), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1142), .A2(new_n1163), .A3(KEYINPUT121), .A4(new_n1198), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1245), .A2(new_n1195), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1218), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1225), .B1(new_n1242), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1132), .A2(KEYINPUT60), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1199), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1125), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n681), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1215), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n793), .A3(new_n824), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(G384), .A3(new_n1215), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1258), .A2(KEYINPUT63), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1241), .B1(new_n1250), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1242), .A2(new_n1249), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT122), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1242), .A2(new_n1249), .A3(KEYINPUT122), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1224), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1225), .A2(G2897), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1256), .A2(new_n1257), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1265), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1263), .A2(new_n1224), .A3(new_n1258), .A4(new_n1264), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1260), .A2(new_n1270), .A3(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1240), .B1(new_n1275), .B2(new_n1250), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1271), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1250), .A2(KEYINPUT62), .A3(new_n1258), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1276), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1280), .B2(new_n1239), .ZN(G405));
  NAND2_X1  g1081(.A1(G375), .A2(new_n1218), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1242), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(KEYINPUT126), .A3(new_n1258), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1258), .A2(KEYINPUT126), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1242), .A3(new_n1282), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  XOR2_X1   g1087(.A(new_n1287), .B(new_n1239), .Z(G402));
endmodule


