

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U326 ( .A(n553), .B(KEYINPUT55), .ZN(n554) );
  XOR2_X1 U327 ( .A(n312), .B(n311), .Z(n556) );
  XNOR2_X1 U328 ( .A(n363), .B(n362), .ZN(n364) );
  NOR2_X1 U329 ( .A1(n546), .A2(n388), .ZN(n385) );
  INV_X1 U330 ( .A(G183GAT), .ZN(n305) );
  XNOR2_X1 U331 ( .A(n306), .B(n305), .ZN(n307) );
  INV_X1 U332 ( .A(KEYINPUT97), .ZN(n360) );
  XNOR2_X1 U333 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U334 ( .A(n308), .B(n307), .ZN(n354) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(n578) );
  XNOR2_X1 U336 ( .A(n555), .B(n554), .ZN(n557) );
  NOR2_X1 U337 ( .A1(n489), .A2(n461), .ZN(n454) );
  XNOR2_X1 U338 ( .A(n454), .B(KEYINPUT38), .ZN(n474) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U340 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n294) );
  XNOR2_X1 U342 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U344 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n296) );
  XOR2_X1 U345 ( .A(G43GAT), .B(G134GAT), .Z(n319) );
  XOR2_X1 U346 ( .A(G15GAT), .B(G127GAT), .Z(n397) );
  XNOR2_X1 U347 ( .A(n319), .B(n397), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U349 ( .A(n298), .B(n297), .Z(n300) );
  NAND2_X1 U350 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U352 ( .A(G99GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n301), .B(G120GAT), .ZN(n437) );
  XOR2_X1 U354 ( .A(n302), .B(n437), .Z(n312) );
  XOR2_X1 U355 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n304) );
  XNOR2_X1 U356 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n308) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G176GAT), .ZN(n306) );
  XOR2_X1 U359 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n310) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n345) );
  XNOR2_X1 U362 ( .A(n354), .B(n345), .ZN(n311) );
  XNOR2_X1 U363 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n417) );
  XOR2_X1 U364 ( .A(KEYINPUT77), .B(KEYINPUT65), .Z(n314) );
  XNOR2_X1 U365 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n313) );
  XOR2_X1 U366 ( .A(n314), .B(n313), .Z(n330) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G92GAT), .Z(n445) );
  XOR2_X1 U368 ( .A(G36GAT), .B(KEYINPUT78), .Z(n355) );
  XOR2_X1 U369 ( .A(n445), .B(n355), .Z(n316) );
  XNOR2_X1 U370 ( .A(G190GAT), .B(G218GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n323) );
  XOR2_X1 U372 ( .A(G29GAT), .B(KEYINPUT7), .Z(n318) );
  XNOR2_X1 U373 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n431) );
  XOR2_X1 U375 ( .A(n319), .B(n431), .Z(n321) );
  NAND2_X1 U376 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U378 ( .A(n323), .B(n322), .Z(n328) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G162GAT), .Z(n371) );
  XOR2_X1 U380 ( .A(KEYINPUT9), .B(KEYINPUT79), .Z(n325) );
  XNOR2_X1 U381 ( .A(G99GAT), .B(G106GAT), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n371), .B(n326), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n568) );
  XOR2_X1 U386 ( .A(KEYINPUT36), .B(n568), .Z(n586) );
  XOR2_X1 U387 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n332) );
  XNOR2_X1 U388 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n338) );
  XOR2_X1 U390 ( .A(KEYINPUT91), .B(KEYINPUT3), .Z(n334) );
  XNOR2_X1 U391 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n369) );
  XOR2_X1 U393 ( .A(n369), .B(KEYINPUT4), .Z(n336) );
  NAND2_X1 U394 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n352) );
  XOR2_X1 U397 ( .A(G148GAT), .B(G155GAT), .Z(n340) );
  XNOR2_X1 U398 ( .A(G120GAT), .B(G127GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U400 ( .A(G57GAT), .B(KEYINPUT6), .Z(n342) );
  XNOR2_X1 U401 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U403 ( .A(n344), .B(n343), .Z(n350) );
  XOR2_X1 U404 ( .A(G85GAT), .B(G162GAT), .Z(n347) );
  XNOR2_X1 U405 ( .A(n345), .B(G134GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(n348), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U409 ( .A(n352), .B(n351), .Z(n384) );
  XNOR2_X1 U410 ( .A(G92GAT), .B(KEYINPUT96), .ZN(n353) );
  XOR2_X1 U411 ( .A(G204GAT), .B(G64GAT), .Z(n446) );
  XOR2_X1 U412 ( .A(n353), .B(n446), .Z(n365) );
  XOR2_X1 U413 ( .A(n355), .B(n354), .Z(n357) );
  NAND2_X1 U414 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n363) );
  XOR2_X1 U416 ( .A(G211GAT), .B(KEYINPUT21), .Z(n359) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(G218GAT), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n368) );
  XNOR2_X1 U419 ( .A(G8GAT), .B(n368), .ZN(n361) );
  XOR2_X1 U420 ( .A(n365), .B(n364), .Z(n491) );
  XOR2_X1 U421 ( .A(n491), .B(KEYINPUT27), .Z(n390) );
  NOR2_X1 U422 ( .A1(n384), .A2(n390), .ZN(n531) );
  XOR2_X1 U423 ( .A(G204GAT), .B(KEYINPUT22), .Z(n367) );
  XNOR2_X1 U424 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n366) );
  XNOR2_X1 U425 ( .A(n367), .B(n366), .ZN(n380) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n378) );
  XNOR2_X1 U427 ( .A(G106GAT), .B(G78GAT), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n370), .B(G148GAT), .ZN(n436) );
  XOR2_X1 U429 ( .A(n436), .B(n371), .Z(n373) );
  NAND2_X1 U430 ( .A1(G228GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n374), .B(KEYINPUT23), .Z(n376) );
  XOR2_X1 U433 ( .A(G22GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U434 ( .A(n398), .B(KEYINPUT92), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n552) );
  XOR2_X1 U438 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n381) );
  XOR2_X1 U439 ( .A(n552), .B(n381), .Z(n495) );
  INV_X1 U440 ( .A(n495), .ZN(n382) );
  NAND2_X1 U441 ( .A1(n531), .A2(n382), .ZN(n512) );
  XOR2_X1 U442 ( .A(KEYINPUT89), .B(n556), .Z(n383) );
  NOR2_X1 U443 ( .A1(n512), .A2(n383), .ZN(n396) );
  INV_X1 U444 ( .A(n384), .ZN(n549) );
  INV_X1 U445 ( .A(n491), .ZN(n546) );
  INV_X1 U446 ( .A(n556), .ZN(n388) );
  NOR2_X1 U447 ( .A1(n385), .A2(n552), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n386), .B(KEYINPUT25), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n387), .B(KEYINPUT99), .ZN(n393) );
  NAND2_X1 U450 ( .A1(n552), .A2(n388), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n389), .B(KEYINPUT26), .ZN(n571) );
  NOR2_X1 U452 ( .A1(n571), .A2(n390), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n391), .B(KEYINPUT98), .ZN(n392) );
  NOR2_X1 U454 ( .A1(n393), .A2(n392), .ZN(n394) );
  NOR2_X1 U455 ( .A1(n549), .A2(n394), .ZN(n395) );
  NOR2_X1 U456 ( .A1(n396), .A2(n395), .ZN(n459) );
  NOR2_X1 U457 ( .A1(n586), .A2(n459), .ZN(n415) );
  XOR2_X1 U458 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U459 ( .A1(G231GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n402) );
  XNOR2_X1 U462 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U464 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U465 ( .A(G1GAT), .B(G8GAT), .Z(n426) );
  XOR2_X1 U466 ( .A(G78GAT), .B(G211GAT), .Z(n406) );
  XNOR2_X1 U467 ( .A(G183GAT), .B(G71GAT), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n426), .B(n407), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U471 ( .A(n410), .B(KEYINPUT80), .Z(n414) );
  XOR2_X1 U472 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n412) );
  XNOR2_X1 U473 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n443) );
  XNOR2_X1 U475 ( .A(n443), .B(KEYINPUT15), .ZN(n413) );
  XOR2_X1 U476 ( .A(n414), .B(n413), .Z(n564) );
  NAND2_X1 U477 ( .A1(n415), .A2(n564), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n489) );
  XOR2_X1 U479 ( .A(G113GAT), .B(G22GAT), .Z(n419) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G197GAT), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U482 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n421) );
  XNOR2_X1 U483 ( .A(G15GAT), .B(KEYINPUT30), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n435) );
  XOR2_X1 U486 ( .A(G141GAT), .B(G50GAT), .Z(n425) );
  XNOR2_X1 U487 ( .A(G43GAT), .B(G36GAT), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n429) );
  AND2_X1 U490 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U492 ( .A(KEYINPUT68), .B(n430), .Z(n433) );
  XNOR2_X1 U493 ( .A(n431), .B(KEYINPUT29), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n532) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n442) );
  XNOR2_X1 U497 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n439) );
  AND2_X1 U498 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n440), .B(KEYINPUT32), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U504 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n448) );
  XNOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  NOR2_X1 U507 ( .A1(n532), .A2(n578), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT76), .B(n453), .Z(n461) );
  NAND2_X1 U509 ( .A1(n556), .A2(n474), .ZN(n456) );
  XNOR2_X1 U510 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n463) );
  NOR2_X1 U511 ( .A1(n568), .A2(n564), .ZN(n457) );
  XOR2_X1 U512 ( .A(KEYINPUT16), .B(n457), .Z(n458) );
  NOR2_X1 U513 ( .A1(n459), .A2(n458), .ZN(n460) );
  XOR2_X1 U514 ( .A(KEYINPUT100), .B(n460), .Z(n476) );
  NOR2_X1 U515 ( .A1(n461), .A2(n476), .ZN(n468) );
  NAND2_X1 U516 ( .A1(n549), .A2(n468), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n463), .B(n462), .ZN(G1324GAT) );
  XOR2_X1 U518 ( .A(G8GAT), .B(KEYINPUT101), .Z(n465) );
  NAND2_X1 U519 ( .A1(n468), .A2(n491), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n465), .B(n464), .ZN(G1325GAT) );
  XOR2_X1 U521 ( .A(G15GAT), .B(KEYINPUT35), .Z(n467) );
  NAND2_X1 U522 ( .A1(n468), .A2(n556), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n467), .B(n466), .ZN(G1326GAT) );
  NAND2_X1 U524 ( .A1(n495), .A2(n468), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT102), .ZN(n470) );
  XNOR2_X1 U526 ( .A(G22GAT), .B(n470), .ZN(G1327GAT) );
  NAND2_X1 U527 ( .A1(n549), .A2(n474), .ZN(n472) );
  XOR2_X1 U528 ( .A(G29GAT), .B(KEYINPUT39), .Z(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(G1328GAT) );
  NAND2_X1 U530 ( .A1(n474), .A2(n491), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U532 ( .A1(n474), .A2(n495), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U534 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n480) );
  XOR2_X1 U535 ( .A(G57GAT), .B(KEYINPUT105), .Z(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT41), .B(n578), .Z(n559) );
  NAND2_X1 U537 ( .A1(n532), .A2(n559), .ZN(n488) );
  NOR2_X1 U538 ( .A1(n476), .A2(n488), .ZN(n485) );
  NAND2_X1 U539 ( .A1(n485), .A2(n549), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1332GAT) );
  NAND2_X1 U542 ( .A1(n491), .A2(n485), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n481), .B(KEYINPUT106), .ZN(n482) );
  XNOR2_X1 U544 ( .A(G64GAT), .B(n482), .ZN(G1333GAT) );
  XOR2_X1 U545 ( .A(G71GAT), .B(KEYINPUT107), .Z(n484) );
  NAND2_X1 U546 ( .A1(n485), .A2(n556), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(G1334GAT) );
  XOR2_X1 U548 ( .A(G78GAT), .B(KEYINPUT43), .Z(n487) );
  NAND2_X1 U549 ( .A1(n485), .A2(n495), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1335GAT) );
  NOR2_X1 U551 ( .A1(n489), .A2(n488), .ZN(n496) );
  NAND2_X1 U552 ( .A1(n549), .A2(n496), .ZN(n490) );
  XNOR2_X1 U553 ( .A(G85GAT), .B(n490), .ZN(G1336GAT) );
  NAND2_X1 U554 ( .A1(n491), .A2(n496), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n492), .B(KEYINPUT108), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G92GAT), .B(n493), .ZN(G1337GAT) );
  NAND2_X1 U557 ( .A1(n556), .A2(n496), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n498) );
  NAND2_X1 U560 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G106GAT), .B(n499), .ZN(G1339GAT) );
  INV_X1 U563 ( .A(n532), .ZN(n573) );
  NAND2_X1 U564 ( .A1(n559), .A2(n573), .ZN(n501) );
  INV_X1 U565 ( .A(KEYINPUT46), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U567 ( .A(n568), .ZN(n542) );
  NOR2_X1 U568 ( .A1(n502), .A2(n568), .ZN(n503) );
  NAND2_X1 U569 ( .A1(n503), .A2(n564), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT47), .ZN(n510) );
  NOR2_X1 U571 ( .A1(n586), .A2(n564), .ZN(n505) );
  XOR2_X1 U572 ( .A(n505), .B(KEYINPUT45), .Z(n508) );
  INV_X1 U573 ( .A(n578), .ZN(n506) );
  NAND2_X1 U574 ( .A1(n532), .A2(n506), .ZN(n507) );
  NOR2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n509) );
  NOR2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(KEYINPUT48), .ZN(n545) );
  NOR2_X1 U578 ( .A1(n545), .A2(n512), .ZN(n513) );
  NAND2_X1 U579 ( .A1(n513), .A2(n556), .ZN(n526) );
  NOR2_X1 U580 ( .A1(n532), .A2(n526), .ZN(n514) );
  XOR2_X1 U581 ( .A(KEYINPUT110), .B(n514), .Z(n515) );
  XNOR2_X1 U582 ( .A(G113GAT), .B(n515), .ZN(G1340GAT) );
  INV_X1 U583 ( .A(n559), .ZN(n535) );
  NOR2_X1 U584 ( .A1(n526), .A2(n535), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n517) );
  XNOR2_X1 U586 ( .A(G120GAT), .B(KEYINPUT112), .ZN(n516) );
  XNOR2_X1 U587 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(G1341GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n521) );
  XNOR2_X1 U590 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n521), .B(n520), .ZN(n523) );
  NOR2_X1 U592 ( .A1(n564), .A2(n526), .ZN(n522) );
  XOR2_X1 U593 ( .A(n523), .B(n522), .Z(G1342GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n525) );
  XNOR2_X1 U595 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n524) );
  XNOR2_X1 U596 ( .A(n525), .B(n524), .ZN(n528) );
  NOR2_X1 U597 ( .A1(n542), .A2(n526), .ZN(n527) );
  XOR2_X1 U598 ( .A(n528), .B(n527), .Z(n529) );
  XNOR2_X1 U599 ( .A(KEYINPUT115), .B(n529), .ZN(G1343GAT) );
  NOR2_X1 U600 ( .A1(n571), .A2(n545), .ZN(n530) );
  NAND2_X1 U601 ( .A1(n531), .A2(n530), .ZN(n541) );
  NOR2_X1 U602 ( .A1(n532), .A2(n541), .ZN(n533) );
  XOR2_X1 U603 ( .A(KEYINPUT118), .B(n533), .Z(n534) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(n534), .ZN(G1344GAT) );
  NOR2_X1 U605 ( .A1(n541), .A2(n535), .ZN(n539) );
  XOR2_X1 U606 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n537) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n536) );
  XNOR2_X1 U608 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U609 ( .A(n539), .B(n538), .ZN(G1345GAT) );
  NOR2_X1 U610 ( .A1(n564), .A2(n541), .ZN(n540) );
  XOR2_X1 U611 ( .A(G155GAT), .B(n540), .Z(G1346GAT) );
  NOR2_X1 U612 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U613 ( .A(KEYINPUT120), .B(n543), .Z(n544) );
  XNOR2_X1 U614 ( .A(G162GAT), .B(n544), .ZN(G1347GAT) );
  NOR2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n548) );
  INV_X1 U616 ( .A(KEYINPUT54), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n548), .B(n547), .ZN(n550) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT64), .B(n551), .Z(n572) );
  NOR2_X1 U620 ( .A1(n572), .A2(n552), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n553) );
  AND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n567), .A2(n573), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT57), .Z(n561) );
  NAND2_X1 U626 ( .A1(n567), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  INV_X1 U630 ( .A(n564), .ZN(n582) );
  NAND2_X1 U631 ( .A1(n567), .A2(n582), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT124), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G183GAT), .B(n566), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT125), .Z(n575) );
  NOR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U639 ( .A1(n584), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n584), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

