//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT68), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n465), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n479), .B2(G2105), .ZN(G160));
  NOR2_X1   g055(.A1(new_n473), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n473), .A2(new_n466), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(KEYINPUT70), .A2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT70), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2105), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n483), .A2(G126), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n466), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .A4(new_n466), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n498), .A2(new_n499), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n502), .A2(new_n503), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n506), .A2(new_n507), .A3(new_n499), .A4(new_n498), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT74), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(new_n519), .A3(G88), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G50), .A3(G543), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT73), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT73), .B1(new_n520), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT75), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n526), .B(new_n518), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n514), .A2(new_n519), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n519), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n531), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n533), .A2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n511), .A2(new_n513), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n540), .B(new_n545), .C1(new_n546), .C2(new_n529), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n529), .A2(new_n552), .B1(new_n532), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n533), .A2(KEYINPUT76), .A3(G53), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n532), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(KEYINPUT9), .A3(new_n565), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n542), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n530), .A2(G91), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n566), .A2(new_n567), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND2_X1  g148(.A1(new_n530), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n533), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT77), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n542), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n519), .A2(G48), .A3(G543), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n529), .ZN(G305));
  AOI22_X1  g160(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n550), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT78), .B(G85), .Z(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n529), .A2(new_n588), .B1(new_n532), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n550), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n529), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n533), .A2(G54), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n529), .B2(new_n596), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n595), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G321));
  XNOR2_X1  g178(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  XNOR2_X1  g182(.A(G297), .B(KEYINPUT81), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NOR2_X1   g185(.A1(new_n601), .A2(G559), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n611), .A2(KEYINPUT82), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT82), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(G868), .C2(new_n555), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n465), .A2(new_n463), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n483), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n481), .A2(G135), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n466), .A2(G111), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n622), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT15), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2435), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2435), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT86), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT87), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT18), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n649), .A2(new_n651), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n654), .B2(KEYINPUT17), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n649), .B2(new_n651), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(KEYINPUT17), .A3(new_n650), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n662), .A2(new_n663), .ZN(new_n669));
  AOI22_X1  g244(.A1(new_n667), .A2(new_n668), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OR3_X1    g245(.A1(new_n664), .A2(new_n669), .A3(new_n666), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n670), .B(new_n671), .C1(new_n668), .C2(new_n667), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT89), .B(G1981), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(G229));
  XOR2_X1   g254(.A(KEYINPUT31), .B(G11), .Z(new_n680));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT30), .B(G28), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(KEYINPUT96), .B1(G5), .B2(G16), .ZN(new_n684));
  OR3_X1    g259(.A1(KEYINPUT96), .A2(G5), .A3(G16), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n684), .B(new_n685), .C1(G301), .C2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(G1961), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(G1961), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n683), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n627), .A2(new_n681), .ZN(new_n691));
  INV_X1    g266(.A(G34), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n692), .A2(KEYINPUT24), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(KEYINPUT24), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n681), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G160), .B2(new_n681), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2084), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n690), .A2(new_n691), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G27), .A2(G29), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G164), .B2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G2078), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n681), .A2(G33), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n463), .A2(G103), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT92), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT25), .ZN(new_n706));
  NAND2_X1  g281(.A1(G115), .A2(G2104), .ZN(new_n707));
  INV_X1    g282(.A(G127), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n473), .B2(new_n708), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n709), .A2(G2105), .B1(new_n481), .B2(G139), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n703), .B1(new_n711), .B2(G29), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT93), .B(G2072), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n698), .A2(new_n702), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(G29), .A2(G32), .ZN(new_n716));
  AOI22_X1  g291(.A1(G129), .A2(new_n483), .B1(new_n481), .B2(G141), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n463), .A2(G105), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT26), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(new_n681), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT94), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n722), .B(new_n724), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G21), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G168), .B2(G16), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT95), .B(G1966), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n715), .A2(KEYINPUT97), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT97), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n698), .A2(new_n730), .A3(new_n714), .A4(new_n702), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(new_n725), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT91), .B1(G4), .B2(G16), .ZN(new_n735));
  OR3_X1    g310(.A1(KEYINPUT91), .A2(G4), .A3(G16), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n735), .B(new_n736), .C1(new_n601), .C2(new_n686), .ZN(new_n737));
  INV_X1    g312(.A(G1348), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n686), .A2(G19), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n555), .B2(new_n686), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1341), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n731), .A2(new_n734), .A3(new_n743), .ZN(new_n744));
  MUX2_X1   g319(.A(G6), .B(G305), .S(G16), .Z(new_n745));
  XOR2_X1   g320(.A(KEYINPUT32), .B(G1981), .Z(new_n746));
  XOR2_X1   g321(.A(new_n745), .B(new_n746), .Z(new_n747));
  AOI21_X1  g322(.A(new_n686), .B1(new_n525), .B2(new_n527), .ZN(new_n748));
  NOR2_X1   g323(.A1(G16), .A2(G22), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n748), .A2(G1971), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(G1971), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n686), .A2(G23), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n577), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT33), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n757), .A2(G1976), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(G1976), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n752), .A2(new_n753), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n753), .B1(new_n752), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT36), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n686), .A2(G24), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n591), .B2(new_n686), .ZN(new_n767));
  INV_X1    g342(.A(G1986), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G25), .A2(G29), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n483), .A2(G119), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n481), .A2(G131), .ZN(new_n772));
  OAI21_X1  g347(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n466), .A2(G107), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n771), .B(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT90), .Z(new_n776));
  AOI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT35), .B(G1991), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n764), .A2(new_n765), .A3(new_n769), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n750), .A2(new_n751), .ZN(new_n781));
  INV_X1    g356(.A(new_n747), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n761), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(KEYINPUT34), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n752), .A2(new_n753), .A3(new_n761), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n784), .A2(new_n769), .A3(new_n785), .A4(new_n779), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT36), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n744), .B1(new_n780), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G35), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G162), .B2(G29), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2090), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n681), .A2(G26), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n483), .A2(G128), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n481), .A2(G140), .ZN(new_n797));
  OR2_X1    g372(.A1(G104), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(new_n681), .ZN(new_n802));
  MUX2_X1   g377(.A(new_n795), .B(new_n802), .S(KEYINPUT28), .Z(new_n803));
  INV_X1    g378(.A(G2067), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n686), .A2(KEYINPUT23), .A3(G20), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n807));
  INV_X1    g382(.A(G20), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G16), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n806), .B(new_n809), .C1(new_n606), .C2(new_n686), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT99), .B(G1956), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT100), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n788), .A2(new_n794), .A3(new_n805), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(G311));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT101), .ZN(new_n816));
  INV_X1    g391(.A(new_n813), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n817), .B(new_n744), .C1(new_n780), .C2(new_n787), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n818), .A2(new_n819), .A3(new_n794), .A4(new_n805), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(G150));
  AOI22_X1  g396(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n550), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n529), .A2(new_n824), .B1(new_n532), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n555), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n551), .B2(new_n554), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT39), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n602), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT102), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n828), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  NAND2_X1  g415(.A1(new_n483), .A2(G130), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n481), .A2(G142), .ZN(new_n842));
  OR2_X1    g417(.A1(G106), .A2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n800), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n619), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n504), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n506), .A2(KEYINPUT103), .A3(new_n499), .A4(new_n498), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n847), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G160), .B(new_n627), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n488), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n706), .A2(KEYINPUT104), .A3(new_n710), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n721), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n775), .B(KEYINPUT105), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n859), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g439(.A1(G166), .A2(G290), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n525), .A2(new_n527), .A3(new_n591), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n577), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(G305), .B(KEYINPUT107), .Z(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n577), .A3(new_n866), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT42), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n869), .ZN(new_n875));
  INV_X1    g450(.A(new_n870), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n867), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT42), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n871), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n831), .B(new_n611), .Z(new_n881));
  NOR2_X1   g456(.A1(G299), .A2(new_n601), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(G299), .A2(new_n601), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n885), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n881), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n880), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n890), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n874), .A2(new_n894), .A3(new_n879), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G868), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n827), .A2(G868), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(G295));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n901), .A3(new_n899), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n612), .B1(new_n893), .B2(new_n895), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT108), .B1(new_n903), .B2(new_n898), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(G331));
  NAND2_X1  g480(.A1(G168), .A2(G301), .ZN(new_n906));
  NAND2_X1  g481(.A1(G171), .A2(G286), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n831), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n907), .A2(new_n906), .B1(new_n829), .B2(new_n830), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n909), .A2(new_n885), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n887), .A2(new_n889), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n909), .A2(new_n910), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n871), .B2(new_n877), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT109), .B1(new_n915), .B2(G37), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n872), .A2(new_n873), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n917), .B(new_n861), .C1(new_n918), .C2(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n914), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n891), .A2(new_n886), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n913), .B(new_n924), .C1(KEYINPUT41), .C2(new_n891), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT110), .B1(new_n913), .B2(new_n885), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n911), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n872), .B2(new_n873), .ZN(new_n930));
  AND4_X1   g505(.A1(KEYINPUT43), .A2(new_n930), .A3(new_n861), .A4(new_n920), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n923), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n930), .A2(new_n920), .A3(new_n922), .A4(new_n861), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n937), .ZN(G397));
  OAI21_X1  g513(.A(new_n583), .B1(new_n529), .B2(new_n584), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT116), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT116), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n583), .B(new_n941), .C1(new_n529), .C2(new_n584), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n582), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT117), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(G1981), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n943), .A2(G1981), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT117), .B1(G305), .B2(G1981), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT49), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n951));
  AOI211_X1 g526(.A(G1976), .B(G288), .C1(new_n949), .C2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(G305), .A2(G1981), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  NAND4_X1  g530(.A1(G160), .A2(new_n504), .A3(G40), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G8), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(KEYINPUT114), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n956), .B2(G8), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n952), .A2(new_n954), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n949), .B(new_n951), .C1(new_n958), .C2(new_n960), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT115), .B(G1976), .Z(new_n963));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(G288), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1976), .ZN(new_n965));
  OAI221_X1 g540(.A(new_n964), .B1(new_n965), .B2(new_n577), .C1(new_n958), .C2(new_n960), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n958), .A2(new_n960), .B1(new_n965), .B2(new_n577), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT52), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n962), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(G166), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(KEYINPUT55), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(KEYINPUT55), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n851), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n849), .B2(new_n850), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n979), .A2(KEYINPUT113), .A3(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n479), .A2(G2105), .ZN(new_n982));
  INV_X1    g557(.A(new_n469), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(G40), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n505), .A2(new_n955), .A3(new_n508), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G1971), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n984), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n504), .A2(new_n955), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G2090), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n975), .B(G8), .C1(new_n988), .C2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n961), .B1(new_n970), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT63), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n973), .A2(new_n974), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n984), .B1(KEYINPUT50), .B2(new_n990), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(KEYINPUT50), .B2(new_n985), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2090), .ZN(new_n1000));
  INV_X1    g575(.A(new_n980), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT113), .B1(new_n979), .B2(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n987), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1971), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n997), .B1(new_n1005), .B2(new_n971), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(new_n969), .A3(new_n994), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n984), .B1(new_n986), .B2(new_n990), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n955), .A4(new_n508), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1966), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT118), .ZN(new_n1013));
  INV_X1    g588(.A(G2084), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n989), .A2(new_n1014), .A3(new_n991), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(new_n1016), .A3(new_n1011), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G8), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G286), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n996), .B1(new_n1007), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n988), .B2(new_n993), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n996), .B1(new_n1023), .B2(new_n997), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(new_n994), .A3(new_n969), .A4(new_n1020), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n995), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G286), .A2(G8), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT123), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n989), .A2(new_n1014), .A3(new_n991), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1016), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1031));
  AOI211_X1 g606(.A(KEYINPUT118), .B(G1966), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1027), .B(new_n1029), .C1(new_n1033), .C2(new_n971), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT51), .B1(new_n1033), .B2(new_n1029), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1029), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n1018), .B2(G8), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1034), .B(KEYINPUT62), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1003), .B2(G2078), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT120), .B1(new_n989), .B2(new_n991), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1961), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n989), .A2(KEYINPUT120), .A3(new_n991), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1010), .B2(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1008), .A2(new_n1009), .A3(KEYINPUT124), .A4(new_n701), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT53), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1042), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G171), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1007), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1019), .A2(new_n1029), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1027), .B1(new_n1018), .B2(new_n1036), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1034), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1040), .A2(new_n1054), .A3(new_n1058), .A4(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(G299), .B(KEYINPUT57), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n981), .A2(new_n987), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1956), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n999), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1064), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1064), .A3(new_n1068), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n989), .A2(KEYINPUT120), .A3(new_n991), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1072), .A2(new_n1043), .A3(G1348), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n956), .A2(G2067), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT119), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1070), .B1(new_n1077), .B2(new_n601), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT60), .B(new_n602), .C1(new_n1073), .C2(new_n1076), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1044), .A2(new_n738), .A3(new_n1046), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1075), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1071), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT61), .B1(new_n1085), .B2(new_n1069), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT61), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1070), .A2(new_n1087), .A3(new_n1071), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1084), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1996), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n987), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT121), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n981), .A2(new_n1093), .A3(new_n1090), .A4(new_n987), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n956), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1098));
  AND3_X1   g673(.A1(new_n1097), .A2(new_n555), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1097), .B2(new_n555), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1078), .B1(new_n1089), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G2078), .B1(new_n978), .B2(new_n980), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n979), .A2(KEYINPUT45), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n984), .B(KEYINPUT125), .Z(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(KEYINPUT53), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1042), .A2(new_n1047), .A3(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G301), .B(KEYINPUT54), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1007), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1052), .A2(new_n1109), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1057), .A3(new_n1034), .A4(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1026), .B(new_n1062), .C1(new_n1102), .C2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1105), .A2(new_n984), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n800), .B(new_n804), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n721), .B(G1996), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n775), .B(new_n778), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1115), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n591), .A2(new_n768), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT111), .Z(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(G1986), .B2(G290), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1122), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT112), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1114), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1119), .A2(new_n778), .A3(new_n776), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n801), .A2(new_n804), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1123), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT46), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1123), .B2(G1996), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1115), .B1(new_n721), .B2(new_n1117), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1115), .A2(KEYINPUT46), .A3(new_n1090), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT47), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1115), .A2(new_n1125), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT48), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1132), .B(new_n1138), .C1(new_n1122), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1129), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g717(.A1(G227), .A2(new_n460), .ZN(new_n1144));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n1145));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g720(.A1(new_n863), .A2(new_n646), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1148));
  NOR2_X1   g722(.A1(new_n1148), .A2(G229), .ZN(new_n1149));
  AND3_X1   g723(.A1(new_n1147), .A2(new_n935), .A3(new_n1149), .ZN(G308));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n935), .A3(new_n1149), .ZN(G225));
endmodule


