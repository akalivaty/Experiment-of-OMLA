//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT92), .B1(new_n187), .B2(G143), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT92), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n187), .A2(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT93), .ZN(new_n196));
  XNOR2_X1  g010(.A(G116), .B(G122), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT93), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n192), .A2(new_n200), .A3(new_n193), .A4(new_n194), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT13), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n192), .A2(new_n203), .B1(new_n187), .B2(G143), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n188), .A2(new_n191), .A3(KEYINPUT13), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n193), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G122), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G116), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n198), .B1(new_n209), .B2(KEYINPUT14), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n210), .B(new_n197), .ZN(new_n211));
  INV_X1    g025(.A(new_n195), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n193), .B1(new_n192), .B2(new_n194), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT9), .B(G234), .ZN(new_n215));
  INV_X1    g029(.A(G217), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n215), .A2(new_n216), .A3(G953), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n207), .A2(KEYINPUT94), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(new_n217), .C1(new_n206), .C2(new_n202), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT94), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n214), .B1(new_n202), .B2(new_n206), .ZN(new_n222));
  INV_X1    g036(.A(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n218), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G478), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n228), .A2(KEYINPUT15), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n227), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G140), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G125), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT16), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT74), .A2(G125), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(new_n232), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n237), .B2(new_n234), .ZN(new_n238));
  INV_X1    g052(.A(G146), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(G237), .A2(G953), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(G143), .A3(G214), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(G143), .B1(new_n241), .B2(G214), .ZN(new_n244));
  OAI21_X1  g058(.A(G131), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n242), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT91), .B1(new_n249), .B2(KEYINPUT17), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n245), .A2(new_n248), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n245), .A2(new_n252), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n240), .A2(new_n250), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G113), .B(G122), .ZN(new_n256));
  INV_X1    g070(.A(G104), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n243), .A2(new_n244), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(KEYINPUT18), .A2(G131), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G140), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n233), .A2(new_n264), .A3(KEYINPUT76), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT76), .B1(new_n233), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n239), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n239), .B2(new_n237), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n261), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n262), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n255), .A2(new_n258), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n258), .B1(new_n255), .B2(new_n270), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n226), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G475), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n276));
  INV_X1    g090(.A(new_n258), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n238), .A2(G146), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n249), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n265), .B2(new_n266), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n236), .B(G140), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT19), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT90), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n239), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n283), .A3(new_n239), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT90), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n279), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n270), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n277), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n271), .ZN(new_n292));
  NOR2_X1   g106(.A1(G475), .A2(G902), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n276), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n293), .ZN(new_n295));
  AOI211_X1 g109(.A(KEYINPUT20), .B(new_n295), .C1(new_n291), .C2(new_n271), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n275), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n231), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(G234), .A2(G237), .ZN(new_n299));
  INV_X1    g113(.A(G953), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n299), .A2(G952), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n299), .A2(G902), .A3(G953), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT21), .B(G898), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G210), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n239), .A2(G143), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n190), .B2(G146), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n239), .A2(KEYINPUT64), .A3(G143), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n309), .B(new_n310), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n190), .A2(G146), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(G143), .B2(new_n239), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(new_n187), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n190), .A2(G146), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT64), .B1(new_n239), .B2(G143), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n311), .A2(new_n190), .A3(G146), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(KEYINPUT0), .A2(G128), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT0), .A2(G128), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n324), .A2(new_n325), .B1(new_n327), .B2(new_n316), .ZN(new_n328));
  MUX2_X1   g142(.A(new_n320), .B(new_n328), .S(G125), .Z(new_n329));
  INV_X1    g143(.A(G224), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G953), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT80), .B1(new_n198), .B2(G104), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(new_n257), .A3(G107), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n198), .A2(KEYINPUT3), .A3(G104), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT3), .B1(new_n198), .B2(G104), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n333), .B(new_n335), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G101), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n257), .B2(G107), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n198), .A2(KEYINPUT3), .A3(G104), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G101), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n333), .A4(new_n335), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G119), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G116), .ZN(new_n348));
  INV_X1    g162(.A(G116), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G119), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT2), .B(G113), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT66), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT66), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n352), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n338), .A2(new_n358), .A3(G101), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n346), .A2(new_n353), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n351), .A2(new_n352), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n348), .A2(KEYINPUT5), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(G113), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n350), .A3(KEYINPUT5), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n257), .A2(G107), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n198), .A2(G104), .ZN(new_n368));
  OAI21_X1  g182(.A(G101), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n345), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n366), .B1(new_n345), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n365), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT85), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n360), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G122), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n360), .A2(new_n372), .A3(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT6), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n377), .B1(new_n373), .B2(KEYINPUT85), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n332), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n365), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n345), .A2(new_n369), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n386), .B(new_n387), .C1(KEYINPUT81), .C2(KEYINPUT86), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n377), .B(KEYINPUT8), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n370), .A2(new_n371), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n388), .B(new_n389), .C1(new_n392), .C2(new_n386), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT7), .B1(new_n330), .B2(G953), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n329), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n380), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n226), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n308), .B1(new_n385), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n332), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n383), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n383), .A2(new_n376), .B1(KEYINPUT6), .B2(new_n380), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n397), .ZN(new_n404));
  AOI21_X1  g218(.A(G902), .B1(new_n404), .B2(new_n393), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n307), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  OAI211_X1 g223(.A(KEYINPUT87), .B(new_n308), .C1(new_n385), .C2(new_n398), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT88), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n408), .A2(new_n413), .A3(new_n409), .A4(new_n410), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n306), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n216), .B1(G234), .B2(new_n226), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n187), .A2(G119), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(KEYINPUT73), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n347), .A2(G128), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT73), .B(KEYINPUT23), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n420), .B(new_n421), .C1(new_n422), .C2(new_n418), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G110), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n421), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT24), .B(G110), .ZN(new_n426));
  INV_X1    g240(.A(new_n278), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n238), .A2(G146), .ZN(new_n428));
  OAI221_X1 g242(.A(new_n424), .B1(new_n425), .B2(new_n426), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n426), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(KEYINPUT75), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n423), .A2(G110), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n278), .B(new_n267), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G137), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n300), .A2(G221), .A3(G234), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n429), .A2(new_n433), .A3(new_n437), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n226), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT25), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n439), .A2(KEYINPUT25), .A3(new_n226), .A4(new_n440), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n417), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n440), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT77), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n416), .A2(G902), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n357), .A2(new_n353), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n320), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n193), .B2(G137), .ZN(new_n455));
  INV_X1    g269(.A(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT11), .A3(G134), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n193), .A2(G137), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n455), .A2(new_n457), .A3(new_n247), .A4(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n193), .A2(G137), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n456), .A2(G134), .ZN(new_n461));
  OAI21_X1  g275(.A(G131), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n314), .A2(KEYINPUT67), .A3(new_n319), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n453), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G131), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n459), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n328), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(KEYINPUT30), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n320), .A2(new_n463), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT65), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n475));
  AOI211_X1 g289(.A(new_n475), .B(KEYINPUT30), .C1(new_n469), .C2(new_n471), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n451), .B(new_n470), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n465), .A2(new_n469), .A3(new_n450), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n479));
  NAND2_X1  g293(.A1(new_n241), .A2(G210), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G101), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n481), .B(new_n482), .Z(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT31), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n477), .A2(KEYINPUT31), .A3(new_n478), .A4(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n483), .B(KEYINPUT69), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n451), .A2(new_n472), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n478), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT28), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n478), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n492), .B2(KEYINPUT71), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n489), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G472), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n488), .A2(KEYINPUT72), .A3(new_n498), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n226), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(G902), .B1(new_n499), .B2(new_n500), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n507), .A2(KEYINPUT32), .A3(new_n502), .A4(new_n503), .ZN(new_n508));
  INV_X1    g322(.A(new_n496), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n465), .A2(new_n469), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n451), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n511), .B2(KEYINPUT28), .ZN(new_n512));
  INV_X1    g326(.A(new_n483), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n478), .A2(new_n491), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(new_n490), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n493), .A3(new_n496), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n489), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n477), .A2(new_n478), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n513), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n514), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n516), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G472), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n506), .A2(new_n508), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G469), .ZN(new_n528));
  XNOR2_X1  g342(.A(G110), .B(G140), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT79), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n300), .A2(G227), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n530), .B(new_n531), .Z(new_n532));
  NOR2_X1   g346(.A1(new_n318), .A2(new_n187), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n314), .B1(new_n533), .B2(new_n324), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n387), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n346), .A2(new_n328), .A3(new_n359), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n453), .A2(KEYINPUT10), .A3(new_n464), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n537), .B(new_n538), .C1(new_n390), .C2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n532), .B1(new_n540), .B2(new_n468), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT84), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n390), .A2(new_n539), .ZN(new_n543));
  INV_X1    g357(.A(new_n468), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n537), .A4(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT84), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n532), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n345), .A2(new_n369), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT81), .ZN(new_n550));
  INV_X1    g364(.A(new_n320), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n345), .A2(new_n366), .A3(new_n369), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT82), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT82), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n550), .A2(new_n555), .A3(new_n551), .A4(new_n552), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n535), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT12), .B1(new_n557), .B2(new_n468), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n553), .A2(KEYINPUT82), .B1(new_n387), .B2(new_n534), .ZN(new_n560));
  AOI211_X1 g374(.A(new_n559), .B(new_n544), .C1(new_n560), .C2(new_n556), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n561), .B2(KEYINPUT83), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(KEYINPUT12), .A3(new_n468), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n548), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n540), .A2(new_n468), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n532), .B1(new_n545), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n528), .B(new_n226), .C1(new_n566), .C2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n545), .A2(new_n567), .A3(new_n532), .ZN(new_n570));
  INV_X1    g384(.A(new_n545), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n562), .B2(new_n565), .ZN(new_n572));
  OAI211_X1 g386(.A(G469), .B(new_n570), .C1(new_n572), .C2(new_n532), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n528), .A2(new_n226), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G221), .B1(new_n215), .B2(G902), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT78), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n415), .A2(new_n449), .A3(new_n527), .A4(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  NOR2_X1   g396(.A1(new_n502), .A2(KEYINPUT95), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n486), .A2(new_n487), .B1(new_n520), .B2(new_n489), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n226), .B1(new_n584), .B2(KEYINPUT72), .ZN(new_n585));
  INV_X1    g399(.A(new_n503), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n583), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n507), .A2(new_n503), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n587), .A2(new_n449), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n409), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n307), .B1(new_n403), .B2(new_n405), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(KEYINPUT96), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n399), .A2(new_n406), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n228), .A2(G902), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n214), .B(KEYINPUT98), .C1(new_n206), .C2(new_n202), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n217), .A2(KEYINPUT97), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n599), .A2(new_n219), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND4_X1   g418(.A1(new_n598), .A2(new_n218), .A3(new_n221), .A4(new_n224), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n597), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n227), .A2(new_n228), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n297), .A2(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n596), .A2(new_n609), .A3(new_n304), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n590), .A2(new_n580), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  INV_X1    g427(.A(new_n297), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n231), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n596), .A2(new_n304), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n590), .A2(new_n580), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  NAND2_X1  g433(.A1(new_n443), .A2(new_n444), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n416), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT99), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n434), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n448), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT100), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n625), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n445), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n587), .A2(new_n630), .A3(new_n589), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n415), .A2(new_n580), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT37), .B(G110), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT101), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n632), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n301), .B1(new_n302), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n615), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n576), .A2(new_n638), .A3(new_n579), .ZN(new_n639));
  INV_X1    g453(.A(new_n596), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n527), .A2(new_n639), .A3(new_n640), .A4(new_n630), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  XOR2_X1   g456(.A(new_n637), .B(KEYINPUT39), .Z(new_n643));
  NAND2_X1  g457(.A1(new_n580), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT40), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n408), .A2(new_n410), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT38), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n621), .A2(new_n625), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n614), .A2(new_n230), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR4_X1   g464(.A1(new_n647), .A2(new_n591), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n644), .A2(KEYINPUT40), .ZN(new_n652));
  INV_X1    g466(.A(new_n522), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n483), .B1(new_n489), .B2(new_n511), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n654), .B2(G902), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n506), .A2(new_n508), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n645), .A2(new_n651), .A3(new_n652), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  INV_X1    g472(.A(new_n637), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n297), .A2(new_n608), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n576), .A2(new_n579), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n527), .A2(new_n662), .A3(new_n640), .A4(new_n630), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT102), .B(G146), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G48));
  INV_X1    g479(.A(new_n548), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n544), .B1(new_n560), .B2(new_n556), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(KEYINPUT83), .A3(KEYINPUT12), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n565), .B(new_n668), .C1(KEYINPUT12), .C2(new_n667), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n568), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(G469), .B1(new_n670), .B2(G902), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n569), .A3(new_n579), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n527), .A2(new_n610), .A3(new_n449), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT41), .B(G113), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NAND4_X1  g490(.A1(new_n527), .A2(new_n449), .A3(new_n616), .A4(new_n673), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  NOR2_X1   g492(.A1(new_n672), .A2(new_n596), .ZN(new_n679));
  INV_X1    g493(.A(new_n306), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n527), .A2(new_n679), .A3(new_n680), .A4(new_n630), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT103), .B(G119), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G21));
  OAI21_X1  g497(.A(G472), .B1(new_n585), .B2(new_n586), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n501), .A2(new_n226), .A3(new_n503), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(KEYINPUT104), .A3(G472), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n649), .A2(new_n593), .A3(new_n305), .A4(new_n595), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n672), .ZN(new_n691));
  INV_X1    g505(.A(new_n489), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n512), .A2(new_n692), .ZN(new_n693));
  AOI211_X1 g507(.A(G472), .B(G902), .C1(new_n693), .C2(new_n488), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n689), .A2(new_n449), .A3(new_n691), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  NAND2_X1  g511(.A1(new_n660), .A2(KEYINPUT106), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n297), .A2(new_n608), .A3(new_n699), .A4(new_n659), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n679), .A2(new_n701), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n685), .B(new_n502), .C1(new_n507), .C2(new_n503), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT104), .B1(new_n687), .B2(G472), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n648), .B(new_n695), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n689), .A2(KEYINPUT105), .A3(new_n648), .A4(new_n695), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n263), .ZN(G27));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n570), .B(KEYINPUT107), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n712), .B(G469), .C1(new_n572), .C2(new_n532), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n569), .A2(new_n713), .A3(new_n575), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n714), .A2(new_n579), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n591), .B1(new_n408), .B2(new_n410), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n701), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n527), .A2(new_n449), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n711), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n579), .A2(new_n701), .A3(new_n716), .A4(new_n714), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(KEYINPUT42), .A3(new_n449), .A4(new_n527), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT108), .B(G131), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G33));
  NAND3_X1  g538(.A1(new_n715), .A2(new_n638), .A3(new_n716), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n718), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n193), .ZN(G36));
  NAND2_X1  g541(.A1(new_n614), .A2(new_n608), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT110), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT43), .Z(new_n730));
  INV_X1    g544(.A(new_n648), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n587), .A2(new_n589), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n732), .A2(KEYINPUT44), .A3(new_n733), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n716), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  OAI211_X1 g553(.A(KEYINPUT45), .B(new_n712), .C1(new_n572), .C2(new_n532), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(G469), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n532), .B1(new_n669), .B2(new_n545), .ZN(new_n744));
  INV_X1    g558(.A(new_n570), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n741), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(G469), .A3(new_n740), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT109), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n739), .B1(new_n750), .B2(new_n574), .ZN(new_n751));
  INV_X1    g565(.A(new_n569), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n747), .A2(new_n749), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n574), .A2(new_n739), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n578), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n643), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n738), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n456), .ZN(G39));
  XNOR2_X1  g573(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n753), .A2(new_n754), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n569), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n574), .B1(new_n747), .B2(new_n749), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(KEYINPUT46), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n579), .B(new_n761), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n716), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n527), .A2(new_n449), .A3(new_n660), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n766), .B(new_n768), .C1(new_n756), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  NOR2_X1   g586(.A1(G952), .A2(G953), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT118), .Z(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n301), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n730), .A2(new_n776), .A3(new_n672), .A4(new_n767), .ZN(new_n777));
  INV_X1    g591(.A(new_n718), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT48), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n673), .A2(new_n449), .A3(new_n301), .A4(new_n716), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n656), .A3(new_n609), .ZN(new_n782));
  INV_X1    g596(.A(G952), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n783), .A3(G953), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n694), .B1(new_n686), .B2(new_n688), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n449), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n776), .A3(new_n730), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n679), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n780), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n716), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n766), .B1(new_n756), .B2(new_n770), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n671), .A2(new_n569), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n579), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n707), .A2(new_n708), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n781), .A2(new_n656), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n297), .A2(new_n608), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n777), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n647), .A2(new_n591), .A3(new_n673), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT117), .Z(new_n805));
  AND3_X1   g619(.A1(new_n805), .A2(KEYINPUT50), .A3(new_n787), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT50), .B1(new_n805), .B2(new_n787), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT51), .B(new_n803), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n790), .B1(new_n799), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n641), .A2(new_n663), .ZN(new_n812));
  INV_X1    g626(.A(new_n702), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n812), .B1(new_n800), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n596), .A2(new_n650), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n715), .A2(new_n731), .A3(new_n659), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n656), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n811), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n412), .A2(new_n414), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n615), .A2(new_n609), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n304), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n590), .A2(new_n821), .A3(new_n580), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n581), .A2(new_n824), .A3(new_n674), .A4(new_n677), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n696), .A2(new_n632), .A3(new_n681), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n630), .A2(new_n298), .A3(new_n659), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n527), .A2(new_n828), .A3(new_n580), .A4(new_n716), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n800), .B2(new_n720), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n726), .B1(new_n719), .B2(new_n721), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n820), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n814), .A2(new_n811), .A3(new_n819), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n709), .A2(new_n812), .A3(KEYINPUT52), .A4(new_n818), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n820), .A2(new_n832), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n810), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n827), .A2(new_n830), .A3(new_n831), .ZN(new_n840));
  INV_X1    g654(.A(new_n708), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT105), .B1(new_n785), .B2(new_n648), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n813), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n812), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n819), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n846), .A3(new_n834), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n837), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n840), .A2(new_n846), .A3(KEYINPUT53), .A4(new_n834), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n809), .B1(new_n839), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n791), .B(KEYINPUT114), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n796), .B1(new_n794), .B2(KEYINPUT115), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n766), .B(new_n857), .C1(new_n756), .C2(new_n770), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n855), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n854), .B1(new_n859), .B2(KEYINPUT116), .ZN(new_n860));
  INV_X1    g674(.A(new_n766), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n755), .B1(KEYINPUT46), .B2(new_n764), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n770), .B1(new_n862), .B2(new_n579), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT115), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n858), .A3(new_n797), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n865), .A2(KEYINPUT116), .A3(new_n793), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n852), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n775), .B1(new_n851), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n449), .A2(new_n579), .A3(new_n409), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT112), .Z(new_n870));
  AOI211_X1 g684(.A(new_n728), .B(new_n870), .C1(KEYINPUT49), .C2(new_n795), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT113), .Z(new_n872));
  OR2_X1    g686(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n647), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n817), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT119), .B1(new_n868), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n808), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n793), .A2(new_n798), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n789), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT54), .B1(new_n848), .B2(new_n849), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n865), .A2(new_n793), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n853), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n859), .A2(KEYINPUT116), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT51), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n774), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n875), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n877), .A2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n300), .A2(G952), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT120), .Z(new_n894));
  OAI211_X1 g708(.A(G210), .B(G902), .C1(new_n835), .C2(new_n838), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n401), .A2(new_n402), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n332), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n403), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n895), .B2(new_n896), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT121), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n894), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(G51));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n574), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n839), .A2(new_n850), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n911));
  INV_X1    g725(.A(new_n670), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n226), .B1(new_n848), .B2(new_n849), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n750), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(new_n912), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT123), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n893), .B1(new_n916), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n292), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n893), .ZN(G60));
  INV_X1    g738(.A(new_n894), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n881), .A2(new_n882), .ZN(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n604), .B2(new_n605), .ZN(new_n931));
  INV_X1    g745(.A(new_n604), .ZN(new_n932));
  INV_X1    g746(.A(new_n605), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n926), .A2(new_n932), .A3(new_n933), .A4(new_n929), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n925), .B1(new_n931), .B2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(new_n848), .A2(new_n849), .ZN(new_n936));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n447), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n624), .A3(new_n938), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n894), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G66));
  OAI21_X1  g759(.A(G953), .B1(new_n303), .B2(new_n330), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n827), .B2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n897), .B1(G898), .B2(new_n300), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  INV_X1    g764(.A(new_n758), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n951), .A2(new_n814), .A3(new_n831), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n756), .A2(new_n778), .A3(new_n643), .A4(new_n815), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n300), .A3(new_n771), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n470), .B1(new_n474), .B2(new_n476), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(new_n284), .Z(new_n956));
  NAND2_X1  g770(.A1(G900), .A2(G953), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n950), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n814), .A2(new_n657), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n822), .B(KEYINPUT124), .ZN(new_n963));
  OR4_X1    g777(.A1(new_n718), .A2(new_n963), .A3(new_n644), .A4(new_n767), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n962), .A2(new_n771), .A3(new_n951), .A4(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n951), .A2(new_n964), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(KEYINPUT125), .A3(new_n771), .A4(new_n962), .ZN(new_n969));
  AOI21_X1  g783(.A(G953), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n959), .B1(new_n970), .B2(new_n956), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n300), .B1(G227), .B2(G900), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n959), .B(new_n974), .C1(new_n970), .C2(new_n956), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(G72));
  NAND3_X1  g790(.A1(new_n967), .A2(new_n969), .A3(new_n827), .ZN(new_n977));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  AOI211_X1 g793(.A(new_n513), .B(new_n653), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n771), .A2(new_n952), .A3(new_n827), .A4(new_n953), .ZN(new_n981));
  INV_X1    g795(.A(new_n979), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n513), .B(new_n653), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n523), .B2(new_n484), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT127), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n893), .B1(new_n936), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n980), .A2(new_n987), .ZN(G57));
endmodule


