//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n471), .B1(G2104), .B2(new_n460), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n473), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(G101), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XOR2_X1   g050(.A(KEYINPUT67), .B(G2105), .Z(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(G137), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(new_n463), .A2(new_n477), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G124), .B1(new_n482), .B2(G136), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n476), .C2(G112), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n460), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n461), .B(new_n462), .C1(new_n489), .C2(new_n490), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n476), .A2(new_n496), .A3(G138), .A4(new_n477), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT70), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n502), .B(G651), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n501), .A2(G543), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G50), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT71), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n500), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(new_n502), .B1(KEYINPUT6), .B2(new_n500), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT72), .B1(new_n521), .B2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(new_n519), .A3(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n518), .A2(G88), .A3(new_n501), .A4(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(G62), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT73), .Z(new_n529));
  OAI21_X1  g104(.A(G651), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n512), .A2(new_n514), .A3(new_n526), .A4(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n525), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n509), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n501), .A2(new_n507), .A3(new_n525), .A4(new_n508), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT74), .B1(new_n539), .B2(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G168));
  NAND2_X1  g122(.A1(new_n510), .A2(G52), .ZN(new_n548));
  AND4_X1   g123(.A1(new_n501), .A2(new_n508), .A3(new_n507), .A4(new_n525), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G90), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n525), .A2(G64), .ZN(new_n551));
  AND2_X1   g126(.A1(G77), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n548), .A2(new_n550), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AND3_X1   g130(.A1(new_n501), .A2(new_n508), .A3(new_n507), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n556), .A2(G43), .A3(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n549), .A2(G81), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n525), .A2(G56), .ZN(new_n559));
  AND2_X1   g134(.A1(G68), .A2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT75), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(KEYINPUT76), .A2(G53), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n556), .A2(new_n569), .A3(G543), .A4(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n509), .B2(new_n570), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n540), .A2(new_n575), .B1(new_n576), .B2(new_n500), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  NAND2_X1  g155(.A1(new_n510), .A2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n549), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND4_X1  g159(.A1(new_n518), .A2(G86), .A3(new_n501), .A4(new_n525), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n518), .A2(G48), .A3(G543), .A4(new_n501), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI211_X1 g162(.A(new_n587), .B(new_n520), .C1(new_n522), .C2(new_n524), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(G305));
  AND2_X1   g167(.A1(new_n525), .A2(G60), .ZN(new_n593));
  AND2_X1   g168(.A1(G72), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT77), .B(G85), .Z(new_n597));
  OAI221_X1 g172(.A(new_n595), .B1(new_n596), .B2(new_n509), .C1(new_n540), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G54), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT78), .B(G66), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n525), .A2(new_n601), .B1(G79), .B2(G543), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n509), .A2(new_n600), .B1(new_n602), .B2(new_n500), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  NOR3_X1   g180(.A1(new_n540), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(new_n540), .B2(new_n605), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n599), .B1(new_n609), .B2(G868), .ZN(G321));
  NOR2_X1   g186(.A1(G299), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g188(.A(new_n612), .B1(G868), .B2(G168), .ZN(G280));
  XNOR2_X1  g189(.A(KEYINPUT79), .B(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(G860), .B2(new_n615), .ZN(G148));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g195(.A1(new_n481), .A2(G123), .B1(new_n482), .B2(G135), .ZN(new_n621));
  OAI221_X1 g196(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n476), .C2(G111), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  OR2_X1    g199(.A1(new_n472), .A2(new_n474), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n477), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  OAI21_X1  g203(.A(new_n624), .B1(new_n628), .B2(G2100), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G2100), .B2(new_n628), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT80), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n651), .B2(new_n648), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n651), .A3(new_n648), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n655), .A2(new_n651), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n667), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n667), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1981), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(G229));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT33), .ZN(new_n689));
  INV_X1    g264(.A(G1976), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n685), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n685), .ZN(new_n693));
  INV_X1    g268(.A(G1971), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G6), .A2(G16), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n585), .A2(new_n586), .A3(new_n591), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n689), .B2(new_n690), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n696), .A2(KEYINPUT34), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(KEYINPUT34), .B1(new_n696), .B2(new_n702), .ZN(new_n704));
  MUX2_X1   g279(.A(G24), .B(G290), .S(G16), .Z(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(G1986), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(G1986), .ZN(new_n707));
  OAI221_X1 g282(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n476), .C2(G107), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n481), .A2(G119), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n482), .A2(G131), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n711), .S(G29), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT86), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT87), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n712), .B(new_n715), .ZN(new_n716));
  NOR4_X1   g291(.A1(new_n706), .A2(new_n707), .A3(KEYINPUT88), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n703), .A2(new_n704), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G32), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT26), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n482), .A2(G141), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n725), .B(new_n727), .C1(G129), .C2(new_n481), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n625), .A2(G105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT96), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n723), .B1(new_n732), .B2(new_n722), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  NOR2_X1   g311(.A1(G27), .A2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G164), .B2(G29), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n735), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n722), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n722), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n748));
  OR2_X1    g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n623), .B2(new_n722), .ZN(new_n752));
  INV_X1    g327(.A(G2084), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT24), .B(G34), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(new_n722), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT94), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n479), .B2(new_n722), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n752), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G2078), .B2(new_n738), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n740), .A2(new_n745), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n685), .A2(G19), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT89), .Z(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n562), .B2(new_n685), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1341), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n722), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT28), .Z(new_n766));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n463), .A2(new_n477), .ZN(new_n768));
  INV_X1    g343(.A(G128), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n463), .A2(new_n477), .A3(KEYINPUT90), .A4(G128), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(G116), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n463), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G140), .B2(new_n482), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n772), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n773), .B1(new_n772), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n766), .B1(new_n781), .B2(G29), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT92), .B(G2067), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n760), .A2(new_n764), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n609), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G4), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1348), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n685), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n577), .B1(new_n572), .B2(new_n573), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n685), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT98), .B(G1956), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n789), .A2(new_n790), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n722), .A2(G33), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(new_n476), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT93), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n476), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT25), .ZN(new_n806));
  NAND2_X1  g381(.A1(G103), .A2(G2104), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n463), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n805), .A2(new_n808), .B1(G139), .B2(new_n482), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n803), .A2(new_n804), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n800), .B1(new_n811), .B2(new_n722), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G2072), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n685), .A2(G5), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G171), .B2(new_n685), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G1961), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n757), .A2(new_n753), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT95), .Z(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n743), .B2(new_n744), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(G1961), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n813), .A2(new_n816), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n685), .A2(G21), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G168), .B2(new_n685), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1966), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n785), .A2(new_n799), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n720), .A2(new_n721), .A3(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  AND2_X1   g402(.A1(new_n525), .A2(G67), .ZN(new_n828));
  AND2_X1   g403(.A1(G80), .A2(G543), .ZN(new_n829));
  OAI21_X1  g404(.A(G651), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n518), .A2(G93), .A3(new_n501), .A4(new_n525), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n518), .A2(G55), .A3(G543), .A4(new_n501), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n836));
  INV_X1    g411(.A(new_n833), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n562), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n836), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n609), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT100), .Z(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n846), .B2(new_n847), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n835), .B1(new_n849), .B2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n623), .B(new_n479), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n485), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n495), .A2(new_n497), .ZN(new_n855));
  INV_X1    g430(.A(new_n492), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n778), .B2(new_n779), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n772), .A2(new_n777), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT91), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n772), .A2(new_n773), .A3(new_n777), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(G164), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n858), .A2(new_n862), .A3(new_n810), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n810), .B1(new_n858), .B2(new_n862), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n863), .A2(new_n864), .A3(new_n731), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n778), .A2(new_n779), .A3(new_n857), .ZN(new_n866));
  AOI21_X1  g441(.A(G164), .B1(new_n860), .B2(new_n861), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n811), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n858), .A2(new_n862), .A3(new_n810), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n732), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n711), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT101), .A4(new_n710), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n627), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI221_X1 g452(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n476), .C2(G118), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n481), .A2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n482), .A2(G142), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n627), .A2(new_n873), .A3(new_n874), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n877), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n877), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n854), .B1(new_n871), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n865), .B2(new_n870), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n888), .A2(new_n865), .A3(new_n870), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(KEYINPUT102), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n888), .B(new_n893), .C1(new_n865), .C2(new_n870), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n854), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n890), .B(KEYINPUT103), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(G395));
  XNOR2_X1  g478(.A(new_n843), .B(new_n617), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n510), .A2(G54), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n602), .A2(new_n500), .ZN(new_n907));
  INV_X1    g482(.A(new_n608), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n906), .B(new_n907), .C1(new_n908), .C2(new_n606), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(G299), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n609), .A2(new_n794), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(G299), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n609), .A2(new_n794), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n904), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT105), .Z(new_n918));
  NOR2_X1   g493(.A1(new_n910), .A2(new_n911), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n904), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(new_n920), .B(KEYINPUT104), .Z(new_n921));
  XNOR2_X1  g496(.A(new_n687), .B(G290), .ZN(new_n922));
  XNOR2_X1  g497(.A(G303), .B(new_n698), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT42), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n918), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n918), .B2(new_n921), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n837), .A2(G868), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(G295));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n929), .ZN(G331));
  AND3_X1   g506(.A1(new_n838), .A2(G168), .A3(new_n842), .ZN(new_n932));
  AOI21_X1  g507(.A(G168), .B1(new_n838), .B2(new_n842), .ZN(new_n933));
  OAI21_X1  g508(.A(G301), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n843), .A2(G286), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n838), .A2(G168), .A3(new_n842), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(G171), .A3(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n934), .A2(new_n937), .A3(new_n919), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n916), .B1(new_n934), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n940), .B2(new_n924), .ZN(new_n941));
  INV_X1    g516(.A(new_n924), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n937), .A3(new_n919), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  AOI211_X1 g520(.A(KEYINPUT106), .B(new_n916), .C1(new_n934), .C2(new_n937), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n941), .A2(new_n947), .A3(KEYINPUT43), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n942), .B1(new_n938), .B2(new_n939), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT43), .B1(new_n941), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n941), .A2(new_n947), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n939), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n924), .A3(new_n943), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n949), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n951), .A2(new_n961), .ZN(G397));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n470), .A2(new_n478), .A3(G40), .A4(new_n475), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G164), .B2(G1384), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1966), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT116), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n857), .A2(new_n973), .A3(new_n963), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n753), .A4(new_n966), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n969), .A2(KEYINPUT116), .A3(new_n970), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(G8), .A3(G286), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n976), .ZN(new_n981));
  OAI211_X1 g556(.A(KEYINPUT123), .B(G8), .C1(new_n981), .C2(new_n971), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n545), .A2(G8), .A3(new_n546), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT124), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(KEYINPUT123), .A2(KEYINPUT51), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n983), .B2(KEYINPUT51), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n978), .B2(G8), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n979), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT62), .B(new_n979), .C1(new_n985), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n969), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n964), .A2(new_n968), .A3(KEYINPUT110), .A4(new_n966), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n694), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n974), .A2(new_n966), .A3(new_n975), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n744), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(KEYINPUT111), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n514), .A2(new_n526), .A3(new_n530), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n509), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1004), .A2(KEYINPUT111), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1009), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G303), .A2(new_n1005), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1002), .A2(KEYINPUT115), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1003), .B1(new_n997), .B2(new_n1000), .ZN(new_n1016));
  AND3_X1   g591(.A1(G303), .A2(new_n1005), .A3(new_n1011), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1011), .B1(G303), .B2(new_n1005), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1016), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n525), .A2(G61), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n500), .B1(new_n1027), .B2(new_n589), .ZN(new_n1028));
  OAI21_X1  g603(.A(G1981), .B1(new_n1028), .B2(KEYINPUT114), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n698), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n591), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G305), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1026), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G164), .A2(G1384), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1003), .B1(new_n1036), .B2(new_n966), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n698), .A2(new_n1029), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G305), .A2(new_n1033), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n581), .A2(new_n582), .A3(G1976), .A4(new_n583), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  INV_X1    g618(.A(G87), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n583), .B1(new_n540), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G49), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n509), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n690), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1037), .A2(new_n1042), .A3(new_n1043), .A4(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1043), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n690), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1053), .A2(KEYINPUT113), .A3(new_n1037), .A4(new_n1042), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1041), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1014), .A2(new_n1020), .A3(new_n1025), .A4(new_n1056), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n999), .A2(G1961), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n736), .A2(KEYINPUT53), .ZN(new_n1059));
  AOI21_X1  g634(.A(G2078), .B1(new_n995), .B2(new_n996), .ZN(new_n1060));
  OAI221_X1 g635(.A(new_n1058), .B1(new_n969), .B2(new_n1059), .C1(new_n1060), .C2(KEYINPUT53), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1057), .A2(G301), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n993), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n966), .A2(new_n964), .A3(new_n968), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1066), .A2(new_n1067), .B1(new_n1068), .B2(new_n998), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1071));
  NAND3_X1  g646(.A1(G299), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n794), .B2(KEYINPUT118), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n964), .A2(new_n968), .A3(new_n966), .A4(new_n1065), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT120), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1069), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n998), .A2(new_n788), .ZN(new_n1080));
  NOR4_X1   g655(.A1(G164), .A2(new_n965), .A3(G1384), .A4(G2067), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g658(.A(KEYINPUT121), .B(new_n1081), .C1(new_n998), .C2(new_n788), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n909), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1075), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1078), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1083), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1080), .A2(new_n1079), .A3(new_n1082), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n609), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1036), .A2(new_n966), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT122), .ZN(new_n1097));
  INV_X1    g672(.A(G1996), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n964), .A2(new_n968), .A3(new_n1098), .A4(new_n966), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(new_n1100), .A3(new_n1095), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1102), .A2(KEYINPUT59), .A3(new_n562), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT59), .B1(new_n1102), .B2(new_n562), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(KEYINPUT60), .B(new_n909), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1093), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n964), .A2(new_n968), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1109), .A2(new_n1067), .A3(new_n966), .A4(new_n1065), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n998), .A2(new_n1068), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1077), .A3(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1108), .B1(new_n1114), .B2(new_n1086), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1078), .A3(KEYINPUT61), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1087), .B1(new_n1107), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(G301), .B(KEYINPUT54), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1061), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n478), .A2(new_n475), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT125), .ZN(new_n1123));
  INV_X1    g698(.A(G40), .ZN(new_n1124));
  INV_X1    g699(.A(new_n470), .ZN(new_n1125));
  NOR4_X1   g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1059), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1120), .B1(new_n1109), .B2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1058), .C1(KEYINPUT53), .C2(new_n1060), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1121), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1057), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(new_n989), .A3(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1017), .A2(new_n1018), .A3(KEYINPUT112), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(new_n1023), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1055), .B1(new_n1133), .B2(new_n1016), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n978), .A2(G8), .A3(G168), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1134), .A2(new_n1020), .A3(new_n1014), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1134), .A2(new_n1140), .A3(new_n1136), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT117), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1134), .A2(new_n1140), .A3(new_n1143), .A4(new_n1136), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1139), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1025), .A2(new_n1055), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1041), .A2(new_n690), .A3(new_n687), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(G1981), .B2(G305), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1037), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1064), .A2(new_n1131), .A3(new_n1145), .A4(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n780), .B(G2067), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT108), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n857), .A2(new_n963), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1153), .A2(new_n967), .A3(new_n966), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n732), .A2(new_n1154), .A3(new_n1098), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1157), .A2(KEYINPUT107), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(KEYINPUT107), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1154), .A2(G1996), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1158), .A2(new_n1159), .B1(new_n732), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n711), .A2(new_n714), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n711), .A2(new_n714), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1155), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(G290), .B(G1986), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1155), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1156), .A2(new_n1161), .A3(new_n1164), .A4(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT109), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1150), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1156), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(G2067), .B2(new_n781), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1156), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1154), .A2(G290), .A3(G1986), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT48), .Z(new_n1174));
  AOI22_X1  g749(.A1(new_n1171), .A2(new_n1155), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1155), .B1(new_n1152), .B2(new_n731), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT46), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1160), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g755(.A(KEYINPUT126), .B(KEYINPUT46), .C1(new_n1154), .C2(G1996), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1180), .A2(new_n1181), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1177), .A2(KEYINPUT47), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT47), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1176), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1185), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1187), .A2(KEYINPUT127), .A3(new_n1183), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1175), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1169), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g765(.A1(new_n899), .A2(new_n900), .ZN(new_n1192));
  NOR4_X1   g766(.A1(G229), .A2(new_n457), .A3(G401), .A4(G227), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n1192), .A2(new_n959), .A3(new_n1193), .ZN(G308));
  NAND3_X1  g768(.A1(new_n1192), .A2(new_n959), .A3(new_n1193), .ZN(G225));
endmodule


