//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT75), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n194), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(KEYINPUT11), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G137), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n202), .A2(new_n208), .A3(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n199), .A2(G134), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n200), .B2(new_n198), .ZN(new_n212));
  OAI22_X1  g026(.A1(KEYINPUT65), .A2(new_n206), .B1(new_n203), .B2(G137), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(G143), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n219), .A2(G143), .ZN(new_n224));
  OAI22_X1  g038(.A1(new_n220), .A2(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(G146), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n218), .A4(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(KEYINPUT76), .ZN(new_n232));
  INV_X1    g046(.A(G107), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT77), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G107), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT76), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT3), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n232), .A2(new_n234), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n231), .B2(G107), .ZN(new_n240));
  AOI21_X1  g054(.A(G101), .B1(new_n231), .B2(G107), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(G104), .B1(new_n234), .B2(new_n236), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n231), .A2(G107), .ZN(new_n244));
  OAI21_X1  g058(.A(G101), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n229), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n229), .B1(new_n242), .B2(new_n245), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n217), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT12), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n242), .A2(new_n245), .ZN(new_n252));
  INV_X1    g066(.A(new_n229), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n246), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT12), .A3(new_n217), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n246), .A2(KEYINPUT10), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n229), .A2(new_n242), .A3(new_n245), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n231), .A2(G107), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n239), .A2(new_n240), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G101), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n265));
  INV_X1    g079(.A(G101), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT4), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n226), .A2(new_n227), .A3(new_n268), .ZN(new_n269));
  OR2_X1    g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n268), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n223), .B2(new_n224), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n263), .A2(new_n267), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n261), .A2(new_n275), .A3(new_n216), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n196), .B1(new_n257), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n196), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n216), .B1(new_n261), .B2(new_n275), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n250), .B(new_n216), .C1(new_n246), .C2(new_n254), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT12), .B1(new_n255), .B2(new_n217), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n196), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n258), .A2(new_n260), .B1(new_n265), .B2(new_n274), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n288), .B2(new_n216), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n261), .A2(new_n275), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n217), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT78), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n190), .B1(new_n282), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G469), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT79), .B(G469), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n283), .A2(new_n284), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(new_n278), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n196), .B1(new_n291), .B2(new_n276), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n190), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n191), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G217), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n188), .A2(new_n302), .A3(G953), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(KEYINPUT67), .A2(G116), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT67), .A2(G116), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(G122), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n308), .A2(G122), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT14), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT14), .ZN(new_n312));
  OAI21_X1  g126(.A(G107), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n234), .A2(new_n236), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n307), .A3(new_n309), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT90), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n221), .B2(G143), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n222), .A2(KEYINPUT90), .A3(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n221), .A2(G143), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n320), .A2(new_n203), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n203), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n316), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n203), .A3(new_n321), .ZN(new_n326));
  INV_X1    g140(.A(new_n316), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n315), .B1(new_n307), .B2(new_n309), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n318), .A2(KEYINPUT13), .A3(new_n319), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT13), .B1(new_n318), .B2(new_n319), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n321), .B(new_n330), .C1(new_n331), .C2(KEYINPUT91), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT91), .ZN(new_n333));
  AOI211_X1 g147(.A(new_n333), .B(KEYINPUT13), .C1(new_n318), .C2(new_n319), .ZN(new_n334));
  OAI21_X1  g148(.A(G134), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n329), .B1(new_n335), .B2(KEYINPUT92), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(G134), .C1(new_n332), .C2(new_n334), .ZN(new_n338));
  AOI211_X1 g152(.A(new_n304), .B(new_n325), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(KEYINPUT92), .ZN(new_n340));
  INV_X1    g154(.A(new_n329), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n325), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n303), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n190), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT15), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G478), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G237), .A2(G953), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n349), .A2(G143), .A3(G214), .ZN(new_n350));
  AOI21_X1  g164(.A(G143), .B1(new_n349), .B2(G214), .ZN(new_n351));
  OAI21_X1  g165(.A(G131), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT17), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n192), .A3(G214), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n222), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n349), .A2(G143), .A3(G214), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n210), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G125), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT69), .B1(new_n361), .B2(KEYINPUT16), .ZN(new_n362));
  INV_X1    g176(.A(G125), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G140), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n364), .A3(KEYINPUT16), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT69), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT16), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n360), .A4(G125), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n362), .A2(new_n365), .A3(G146), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(new_n365), .A3(new_n368), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n219), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT17), .B(G131), .C1(new_n350), .C2(new_n351), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n359), .A2(new_n369), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(KEYINPUT18), .A2(G131), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n356), .A2(new_n357), .A3(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT18), .B(G131), .C1(new_n350), .C2(new_n351), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n363), .A2(G140), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n360), .A2(G125), .ZN(new_n378));
  OAI21_X1  g192(.A(G146), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n361), .A2(new_n364), .A3(new_n219), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n379), .A2(KEYINPUT85), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT85), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n375), .B(new_n376), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G113), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n231), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n373), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT87), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n373), .A2(new_n383), .A3(new_n388), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n385), .B1(new_n373), .B2(new_n383), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT89), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n392), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n190), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n377), .A2(new_n378), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT19), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT19), .B1(new_n397), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n219), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n352), .A2(new_n358), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n369), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n385), .B1(new_n403), .B2(new_n383), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n390), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT20), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT88), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n404), .B1(new_n387), .B2(new_n389), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n412), .B2(new_n409), .ZN(new_n413));
  AOI22_X1  g227(.A1(G475), .A2(new_n396), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G952), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  INV_X1    g230(.A(G234), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n354), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n190), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(G898), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n348), .A2(new_n414), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT2), .B(G113), .ZN(new_n426));
  INV_X1    g240(.A(new_n306), .ZN(new_n427));
  NOR2_X1   g241(.A1(KEYINPUT67), .A2(G116), .ZN(new_n428));
  INV_X1    g242(.A(G119), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n308), .A2(G119), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n426), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n305), .A2(G119), .A3(new_n306), .ZN(new_n434));
  INV_X1    g248(.A(new_n431), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n432), .A2(new_n436), .B1(new_n263), .B2(new_n267), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n265), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n252), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n430), .A2(new_n431), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(KEYINPUT5), .A3(new_n435), .ZN(new_n441));
  INV_X1    g255(.A(G113), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n440), .A2(new_n433), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT80), .ZN(new_n448));
  XOR2_X1   g262(.A(G110), .B(G122), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n265), .A2(new_n437), .B1(new_n439), .B2(new_n445), .ZN(new_n453));
  INV_X1    g267(.A(new_n451), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT80), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n453), .B2(new_n450), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n447), .A2(new_n449), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n229), .A2(new_n363), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n273), .A2(new_n270), .A3(new_n269), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G224), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G953), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT81), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n464), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n456), .A2(new_n460), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(KEYINPUT7), .B1(new_n465), .B2(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n461), .A2(new_n463), .A3(new_n470), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n453), .B2(new_n450), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n449), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT83), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n242), .A2(new_n245), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n445), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n445), .B2(new_n479), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n483), .B(KEYINPUT84), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n469), .B2(new_n482), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n425), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n424), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n301), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n302), .B1(G234), .B2(new_n190), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT22), .B(G137), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n371), .A2(new_n369), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n429), .B2(G128), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n429), .A2(G128), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G110), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT24), .B(G110), .Z(new_n506));
  XNOR2_X1  g320(.A(G119), .B(G128), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n504), .A2(G110), .B1(new_n506), .B2(new_n507), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n369), .A3(new_n380), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(KEYINPUT72), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n509), .B1(new_n369), .B2(new_n371), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n512), .A2(new_n369), .A3(new_n380), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n498), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n511), .A2(new_n513), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n497), .B1(new_n520), .B2(new_n515), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT25), .B1(new_n522), .B2(new_n190), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n524));
  NOR4_X1   g338(.A1(new_n519), .A2(new_n521), .A3(new_n524), .A4(G902), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n492), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n514), .A2(new_n518), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n497), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n518), .A2(new_n498), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n190), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n524), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT73), .A3(new_n492), .ZN(new_n536));
  INV_X1    g350(.A(new_n492), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n190), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT74), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n522), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n528), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n432), .A2(new_n436), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n462), .B1(new_n209), .B2(new_n215), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n212), .A2(new_n214), .A3(new_n210), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT66), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n200), .B1(new_n204), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n549));
  OAI21_X1  g363(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n229), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n544), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n544), .A3(new_n551), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n553), .A2(KEYINPUT28), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(KEYINPUT28), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n349), .A2(G210), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT27), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G101), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT29), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n553), .B(KEYINPUT28), .ZN(new_n565));
  OAI21_X1  g379(.A(G131), .B1(new_n202), .B2(new_n208), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT64), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n566), .A2(new_n546), .B1(new_n462), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n271), .A2(KEYINPUT64), .A3(new_n273), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n202), .A2(new_n208), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n570), .A2(new_n210), .B1(new_n228), .B2(new_n225), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n568), .A2(new_n569), .B1(new_n571), .B2(new_n550), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n572), .A2(new_n544), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n562), .B1(new_n574), .B2(new_n561), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n545), .A2(KEYINPUT30), .A3(new_n551), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n543), .B(new_n576), .C1(new_n572), .C2(KEYINPUT30), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n553), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n560), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n564), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n574), .A2(new_n561), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT68), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n553), .A2(new_n584), .A3(new_n560), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n553), .B2(new_n560), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT31), .B1(new_n587), .B2(new_n577), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n553), .A2(new_n560), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT68), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n553), .A2(new_n584), .A3(new_n560), .ZN(new_n591));
  AND4_X1   g405(.A1(KEYINPUT31), .A2(new_n577), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n583), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G472), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n593), .A2(KEYINPUT32), .A3(new_n594), .A4(new_n190), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT32), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n560), .B1(new_n565), .B2(new_n573), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n577), .A2(new_n590), .A3(new_n591), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT31), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n587), .A2(KEYINPUT31), .A3(new_n577), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n594), .A2(new_n190), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n596), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n582), .A2(new_n595), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n542), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n491), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n266), .ZN(G3));
  NAND2_X1  g422(.A1(new_n484), .A2(KEYINPUT94), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n469), .A2(new_n482), .ZN(new_n610));
  INV_X1    g424(.A(new_n483), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n469), .A2(new_n613), .A3(new_n482), .A4(new_n483), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n609), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n425), .A3(new_n423), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n407), .B1(new_n406), .B2(new_n410), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n412), .A2(KEYINPUT20), .A3(new_n409), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n391), .B(KEYINPUT89), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n619), .B2(new_n390), .ZN(new_n620));
  INV_X1    g434(.A(G475), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n617), .A2(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n190), .A2(G478), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n339), .B2(new_n344), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n342), .A2(new_n343), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n304), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n342), .A2(new_n343), .A3(new_n303), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT95), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(KEYINPUT33), .B(new_n625), .C1(new_n629), .C2(new_n624), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n339), .B2(new_n344), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(KEYINPUT96), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n623), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n345), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(G478), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n622), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n616), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n528), .A2(new_n536), .A3(new_n541), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n594), .A2(KEYINPUT93), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n602), .B2(G902), .ZN(new_n643));
  INV_X1    g457(.A(new_n642), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n593), .A2(new_n190), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n301), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NOR2_X1   g465(.A1(new_n348), .A2(new_n622), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n425), .A2(new_n652), .A3(new_n615), .A4(new_n423), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n648), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT35), .B(G107), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(new_n646), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n301), .A2(new_n490), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n520), .B(KEYINPUT97), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n540), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n528), .A2(new_n536), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n528), .A2(new_n536), .A3(KEYINPUT98), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n659), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT37), .B(G110), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  AND2_X1   g485(.A1(new_n615), .A2(new_n425), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n345), .A2(new_n346), .A3(G478), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n627), .A2(new_n628), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n190), .A3(new_n347), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n414), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n419), .B1(new_n420), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n672), .A2(KEYINPUT99), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n301), .A2(new_n666), .A3(new_n605), .A4(new_n667), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XOR2_X1   g503(.A(new_n679), .B(KEYINPUT39), .Z(new_n690));
  AND2_X1   g504(.A1(new_n301), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  INV_X1    g508(.A(new_n553), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n561), .B1(new_n695), .B2(new_n552), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n598), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n697), .B2(G902), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n595), .A2(new_n604), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n595), .A2(new_n604), .A3(KEYINPUT100), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n485), .A2(new_n488), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT38), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n396), .A2(G475), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n411), .A2(new_n413), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n706), .A2(new_n707), .B1(new_n673), .B2(new_n675), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n425), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n705), .A2(new_n664), .A3(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n693), .A2(new_n694), .A3(new_n703), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND2_X1  g526(.A1(new_n615), .A2(new_n425), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n686), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n624), .B1(new_n674), .B2(new_n631), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n625), .A2(KEYINPUT33), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n634), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n623), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n637), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  INV_X1    g536(.A(new_n679), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n722), .A3(new_n622), .A4(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n622), .B(new_n723), .C1(new_n635), .C2(new_n637), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT101), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n714), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  AND2_X1   g544(.A1(new_n542), .A2(new_n605), .ZN(new_n731));
  INV_X1    g545(.A(new_n191), .ZN(new_n732));
  INV_X1    g546(.A(G469), .ZN(new_n733));
  INV_X1    g547(.A(new_n276), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n286), .B1(new_n734), .B2(new_n279), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n257), .A2(new_n289), .ZN(new_n736));
  AOI21_X1  g550(.A(G902), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n300), .B(new_n732), .C1(new_n733), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT102), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n298), .A2(new_n299), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n732), .A4(new_n300), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n640), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT41), .B(G113), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n654), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n308), .ZN(G18));
  NAND2_X1  g564(.A1(new_n739), .A2(new_n743), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n713), .A3(new_n424), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n605), .A3(new_n666), .A4(new_n667), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  NAND3_X1  g568(.A1(new_n739), .A2(new_n743), .A3(new_n423), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n602), .A2(G902), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n600), .A2(new_n601), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n556), .A2(new_n560), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g573(.A1(new_n756), .A2(new_n594), .B1(new_n759), .B2(new_n603), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n755), .A2(new_n641), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n453), .A2(new_n450), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n472), .A2(new_n473), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n481), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n190), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n452), .A2(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n766), .B2(new_n468), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n614), .B1(new_n767), .B2(new_n483), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n613), .B1(new_n767), .B2(new_n483), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n708), .B(new_n425), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT103), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n615), .A2(KEYINPUT103), .A3(new_n425), .A4(new_n708), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n761), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n761), .A2(new_n774), .A3(KEYINPUT104), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G122), .ZN(G24));
  AOI21_X1  g594(.A(new_n603), .B1(new_n757), .B2(new_n758), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n593), .A2(new_n190), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(G472), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n744), .A2(new_n672), .A3(new_n664), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT105), .B1(new_n727), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n664), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n751), .A3(new_n713), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT105), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n724), .A4(new_n726), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G125), .ZN(G27));
  AOI22_X1  g605(.A1(new_n251), .A2(new_n256), .B1(new_n288), .B2(new_n216), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n292), .B1(new_n792), .B2(new_n196), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n190), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(G469), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n191), .B1(new_n795), .B2(new_n300), .ZN(new_n796));
  INV_X1    g610(.A(new_n425), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n485), .A2(new_n488), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n799), .A2(new_n542), .A3(new_n605), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(KEYINPUT42), .A3(new_n724), .A4(new_n726), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT42), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n542), .A3(new_n605), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n802), .B1(new_n727), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  NAND4_X1  g620(.A1(new_n799), .A2(new_n542), .A3(new_n605), .A4(new_n680), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT106), .B(G134), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G36));
  INV_X1    g623(.A(new_n798), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n721), .A2(new_n414), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT43), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(KEYINPUT43), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n664), .A2(new_n646), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n810), .B1(new_n816), .B2(KEYINPUT44), .ZN(new_n817));
  NAND2_X1  g631(.A1(G469), .A2(G902), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n282), .A2(new_n293), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT45), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n821));
  OAI21_X1  g635(.A(G469), .B1(new_n793), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT46), .B(new_n818), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(KEYINPUT107), .A3(new_n300), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n820), .A2(new_n822), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(G469), .B2(G902), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n826), .B2(KEYINPUT46), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT107), .B1(new_n823), .B2(new_n300), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n732), .B(new_n690), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n815), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT44), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n817), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(KEYINPUT108), .B(G137), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(G39));
  OAI21_X1  g650(.A(new_n732), .B1(new_n827), .B2(new_n828), .ZN(new_n837));
  NAND2_X1  g651(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n542), .A2(new_n605), .A3(new_n810), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n728), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n837), .B1(new_n845), .B2(new_n839), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  AND3_X1   g662(.A1(new_n812), .A2(new_n419), .A3(new_n813), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n751), .A2(new_n810), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n703), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n542), .A3(new_n419), .A4(new_n850), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n719), .A2(new_n414), .A3(new_n720), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n851), .A2(new_n786), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n760), .A2(new_n641), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n705), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n744), .A2(new_n797), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n858), .A2(KEYINPUT50), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  INV_X1    g679(.A(new_n863), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n857), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n855), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n741), .A2(new_n300), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n840), .A2(new_n846), .B1(new_n191), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n858), .A2(new_n798), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n868), .B(KEYINPUT51), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n851), .A2(KEYINPUT118), .A3(new_n606), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT118), .B1(new_n851), .B2(new_n606), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(KEYINPUT48), .A3(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n849), .A2(new_n672), .A3(new_n744), .A4(new_n856), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n853), .A2(new_n638), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n416), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT117), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT48), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n874), .A2(new_n875), .A3(new_n878), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n425), .B(new_n423), .C1(new_n485), .C2(new_n488), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n677), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n647), .A2(new_n301), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n659), .B2(new_n668), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT111), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n648), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n638), .A2(new_n887), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n301), .A2(new_n490), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n893), .A2(new_n894), .B1(new_n895), .B2(new_n731), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n889), .B(KEYINPUT111), .C1(new_n659), .C2(new_n668), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n783), .A2(new_n664), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n724), .A2(new_n726), .A3(new_n899), .A4(new_n799), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n622), .A2(new_n676), .A3(new_n679), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT112), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n798), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n901), .B2(new_n798), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n900), .B(new_n807), .C1(new_n686), .C2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n886), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n638), .A2(new_n887), .ZN(new_n908));
  OAI22_X1  g722(.A1(new_n908), .A2(new_n648), .B1(new_n491), .B2(new_n606), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n891), .B2(new_n890), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n807), .B1(new_n905), .B2(new_n686), .ZN(new_n911));
  INV_X1    g725(.A(new_n900), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n910), .A2(new_n913), .A3(KEYINPUT114), .A4(new_n897), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n731), .B(new_n744), .C1(new_n639), .C2(new_n653), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n761), .A2(new_n774), .A3(KEYINPUT104), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT104), .B1(new_n761), .B2(new_n774), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n753), .B(new_n916), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT115), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n753), .A2(new_n916), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT115), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n779), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n801), .B2(new_n804), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n920), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT52), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT73), .B1(new_n535), .B2(new_n492), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n527), .B(new_n537), .C1(new_n533), .C2(new_n534), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(new_n663), .A3(new_n796), .A4(new_n723), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n701), .B2(new_n702), .ZN(new_n932));
  AOI22_X1  g746(.A1(new_n714), .A2(new_n728), .B1(new_n774), .B2(new_n932), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n927), .A2(new_n933), .A3(new_n790), .A4(new_n688), .ZN(new_n934));
  XOR2_X1   g748(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n935));
  AOI22_X1  g749(.A1(new_n785), .A2(new_n789), .B1(new_n685), .B2(new_n687), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n933), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n915), .A2(new_n926), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n933), .A2(new_n790), .A3(new_n688), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT52), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n927), .A3(new_n933), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n919), .A2(new_n898), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n906), .B1(new_n804), .B2(new_n801), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n941), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n924), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n939), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(KEYINPUT53), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n913), .A2(new_n805), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n919), .A3(new_n898), .ZN(new_n951));
  INV_X1    g765(.A(new_n935), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n940), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n951), .A2(new_n924), .A3(new_n942), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n949), .A2(KEYINPUT54), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n948), .A2(new_n955), .ZN(new_n956));
  OAI22_X1  g770(.A1(new_n885), .A2(new_n956), .B1(G952), .B2(G953), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n869), .B(KEYINPUT49), .Z(new_n958));
  NAND3_X1  g772(.A1(new_n542), .A2(new_n732), .A3(new_n425), .ZN(new_n959));
  OR4_X1    g773(.A1(new_n859), .A2(new_n958), .A3(new_n811), .A4(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n957), .B1(new_n703), .B2(new_n960), .ZN(G75));
  NAND2_X1  g775(.A1(new_n415), .A2(G953), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT119), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n939), .A2(new_n946), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(G902), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(new_n487), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n766), .B(new_n468), .Z(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT55), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT56), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n963), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n964), .A2(G210), .A3(G902), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n968), .B1(new_n972), .B2(new_n969), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n973), .ZN(G51));
  INV_X1    g788(.A(new_n963), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n818), .B(KEYINPUT57), .Z(new_n976));
  INV_X1    g790(.A(new_n948), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n947), .B1(new_n939), .B2(new_n946), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n740), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n964), .A2(G902), .A3(new_n825), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(G54));
  NAND2_X1  g797(.A1(KEYINPUT58), .A2(G475), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n965), .A2(new_n406), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n406), .B1(new_n965), .B2(new_n984), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n975), .B1(new_n985), .B2(new_n986), .ZN(G60));
  NAND2_X1  g801(.A1(G478), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT59), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n956), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT120), .ZN(new_n992));
  INV_X1    g806(.A(new_n717), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n892), .A2(new_n897), .A3(new_n896), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n753), .A2(new_n916), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n777), .B2(new_n778), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n944), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n927), .B1(new_n936), .B2(new_n933), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(KEYINPUT53), .B1(new_n1000), .B2(new_n942), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n953), .A2(new_n942), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n907), .A2(new_n914), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n920), .A2(new_n925), .A3(new_n923), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(KEYINPUT54), .B1(new_n1001), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n948), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n993), .A2(new_n989), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n975), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n989), .B1(new_n948), .B2(new_n955), .ZN(new_n1010));
  OAI21_X1  g824(.A(KEYINPUT120), .B1(new_n1010), .B2(new_n717), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n994), .A2(new_n1009), .A3(new_n1011), .ZN(G63));
  INV_X1    g826(.A(KEYINPUT61), .ZN(new_n1013));
  XNOR2_X1  g827(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n302), .A2(new_n190), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n939), .B2(new_n946), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n662), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n963), .B1(new_n1018), .B2(new_n522), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1013), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n1018), .A2(new_n522), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1023), .A2(KEYINPUT61), .A3(new_n963), .A4(new_n1019), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1024), .ZN(G66));
  NOR3_X1   g839(.A1(new_n421), .A2(new_n465), .A3(new_n192), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n943), .B2(new_n192), .ZN(new_n1027));
  INV_X1    g841(.A(G898), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n766), .B1(new_n1028), .B2(G953), .ZN(new_n1029));
  XNOR2_X1  g843(.A(KEYINPUT122), .B(KEYINPUT123), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1027), .B(new_n1031), .ZN(G69));
  OAI21_X1  g846(.A(new_n576), .B1(new_n572), .B2(KEYINPUT30), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n399), .A2(new_n400), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1034), .B(KEYINPUT124), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1033), .B(new_n1035), .Z(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n638), .A2(new_n677), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n691), .A2(new_n731), .A3(new_n798), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n834), .A2(new_n192), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n936), .A2(new_n711), .A3(new_n729), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(KEYINPUT62), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n847), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n1042), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1042), .A2(KEYINPUT62), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT125), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1041), .B(new_n1045), .C1(new_n1046), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(G227), .ZN(new_n1051));
  NOR3_X1   g865(.A1(new_n1051), .A2(new_n678), .A3(new_n192), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1037), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n830), .A2(new_n731), .A3(new_n774), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n834), .A2(new_n805), .A3(new_n807), .A4(new_n1055), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n847), .A2(new_n729), .A3(new_n936), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n192), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1051), .A2(G900), .A3(G953), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n1036), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g874(.A(KEYINPUT126), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1062), .A2(new_n1037), .ZN(new_n1063));
  INV_X1    g877(.A(KEYINPUT126), .ZN(new_n1064));
  NOR2_X1   g878(.A1(new_n1049), .A2(new_n1046), .ZN(new_n1065));
  NOR2_X1   g879(.A1(new_n1065), .A2(new_n1044), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1052), .B1(new_n1066), .B2(new_n1041), .ZN(new_n1067));
  OAI211_X1 g881(.A(new_n1063), .B(new_n1064), .C1(new_n1067), .C2(new_n1037), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1061), .A2(new_n1068), .ZN(G72));
  NAND2_X1  g883(.A1(new_n578), .A2(new_n560), .ZN(new_n1070));
  NAND4_X1  g884(.A1(new_n1066), .A2(new_n834), .A3(new_n943), .A4(new_n1039), .ZN(new_n1071));
  NAND2_X1  g885(.A1(G472), .A2(G902), .ZN(new_n1072));
  XOR2_X1   g886(.A(new_n1072), .B(KEYINPUT63), .Z(new_n1073));
  AOI21_X1  g887(.A(new_n1070), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g888(.A(new_n1073), .ZN(new_n1075));
  INV_X1    g889(.A(new_n580), .ZN(new_n1076));
  AOI21_X1  g890(.A(new_n1075), .B1(new_n1076), .B2(new_n598), .ZN(new_n1077));
  NAND3_X1  g891(.A1(new_n949), .A2(new_n954), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n1075), .B1(new_n1079), .B2(new_n943), .ZN(new_n1080));
  NAND2_X1  g894(.A1(new_n579), .A2(new_n561), .ZN(new_n1081));
  XNOR2_X1  g895(.A(new_n1081), .B(KEYINPUT127), .ZN(new_n1082));
  OAI211_X1 g896(.A(new_n963), .B(new_n1078), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g897(.A1(new_n1074), .A2(new_n1083), .ZN(G57));
endmodule


