//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT68), .A2(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT68), .A2(G119), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G116), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT67), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(KEYINPUT67), .A3(new_n195), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  OAI21_X1  g016(.A(G128), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(KEYINPUT65), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  AOI21_X1  g020(.A(G146), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n203), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT66), .B1(new_n200), .B2(G146), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n208), .A3(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n206), .A3(G146), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G137), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT11), .A3(G134), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(G137), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n221), .A2(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n223), .A2(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n214), .A2(new_n215), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n207), .B2(new_n209), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT11), .B1(new_n223), .B2(G134), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n229), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n225), .B1(new_n239), .B2(new_n224), .ZN(new_n240));
  INV_X1    g054(.A(new_n227), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n234), .B(new_n237), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n232), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT30), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT30), .ZN(new_n246));
  AOI211_X1 g060(.A(KEYINPUT64), .B(new_n246), .C1(new_n232), .C2(new_n242), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n199), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n243), .ZN(new_n254));
  INV_X1    g068(.A(new_n199), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n248), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n248), .A2(new_n259), .A3(new_n253), .A4(new_n256), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(KEYINPUT31), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n253), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n243), .A2(new_n199), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n256), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n243), .A2(new_n199), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT28), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n262), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n248), .A2(new_n269), .A3(new_n253), .A4(new_n256), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AOI211_X1 g085(.A(G472), .B(G902), .C1(new_n261), .C2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n187), .B1(new_n272), .B2(KEYINPUT70), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n271), .ZN(new_n274));
  INV_X1    g088(.A(G472), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT32), .ZN(new_n279));
  INV_X1    g093(.A(new_n248), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(new_n266), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n281), .B2(new_n253), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n262), .C1(new_n280), .C2(new_n266), .ZN(new_n285));
  OR3_X1    g099(.A1(new_n265), .A2(new_n262), .A3(new_n267), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n282), .A2(new_n283), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n287), .B(new_n276), .C1(new_n283), .C2(new_n286), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n273), .A2(new_n279), .B1(G472), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G217), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(G234), .B2(new_n276), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(G902), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n292), .B(KEYINPUT76), .Z(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n295));
  XNOR2_X1  g109(.A(G125), .B(G140), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT16), .ZN(new_n297));
  INV_X1    g111(.A(G125), .ZN(new_n298));
  OR3_X1    g112(.A1(new_n298), .A2(KEYINPUT16), .A3(G140), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(G146), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n296), .A2(new_n208), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n216), .A2(KEYINPUT23), .A3(G119), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT72), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n188), .A2(new_n189), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n216), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n188), .A2(G128), .A3(new_n189), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n306), .A2(new_n307), .B1(KEYINPUT23), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n216), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G110), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n308), .B1(new_n314), .B2(G128), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT24), .B(G110), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n302), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n300), .ZN(new_n319));
  AOI21_X1  g133(.A(G146), .B1(new_n297), .B2(new_n299), .ZN(new_n320));
  OAI22_X1  g134(.A1(new_n319), .A2(new_n320), .B1(new_n315), .B2(new_n316), .ZN(new_n321));
  INV_X1    g135(.A(new_n311), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(G110), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n295), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n315), .A2(new_n316), .ZN(new_n325));
  INV_X1    g139(.A(new_n320), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(new_n300), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n311), .B2(new_n312), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n311), .A2(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n328), .B(KEYINPUT74), .C1(new_n329), .C2(new_n302), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT22), .B(G137), .ZN(new_n331));
  INV_X1    g145(.A(G953), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(G221), .A3(G234), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n324), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n328), .B(new_n334), .C1(new_n329), .C2(new_n302), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n337), .B1(new_n336), .B2(new_n338), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n294), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n276), .A3(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT25), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n336), .A2(new_n345), .A3(new_n276), .A4(new_n338), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n291), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n341), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n289), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n350));
  OAI21_X1  g164(.A(G221), .B1(new_n350), .B2(G902), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n351), .B(KEYINPUT77), .Z(new_n352));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n240), .A2(new_n241), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G104), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G101), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G107), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT78), .A4(G104), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n360), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n361), .B1(new_n359), .B2(new_n363), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT79), .B1(new_n365), .B2(new_n367), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n210), .B(new_n218), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n214), .A2(new_n215), .ZN(new_n373));
  OAI21_X1  g187(.A(G128), .B1(new_n207), .B2(new_n202), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n365), .A2(new_n367), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n354), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n353), .B1(new_n378), .B2(KEYINPUT12), .ZN(new_n379));
  INV_X1    g193(.A(new_n354), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n362), .A2(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n364), .A2(new_n363), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n386), .A2(new_n387), .A3(G101), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n381), .B1(new_n388), .B2(new_n366), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n219), .B1(new_n389), .B2(new_n368), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n375), .A2(new_n376), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n380), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT12), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(KEYINPUT81), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n378), .A2(KEYINPUT12), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n379), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT10), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n375), .B2(new_n376), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n210), .B2(new_n218), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(new_n368), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n403), .B(G101), .C1(new_n386), .C2(new_n387), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n402), .A2(new_n234), .A3(new_n237), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n354), .B(KEYINPUT80), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G110), .B(G140), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n332), .A2(G227), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n406), .A2(KEYINPUT82), .A3(new_n380), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT82), .B1(new_n406), .B2(new_n380), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n408), .A2(new_n412), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n409), .A2(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G469), .B1(new_n418), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT83), .A3(new_n413), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n396), .A2(new_n417), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT83), .B1(new_n421), .B2(new_n413), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n420), .B(new_n276), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n352), .B1(new_n419), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n199), .A2(new_n404), .A3(new_n402), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G122), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n190), .A2(KEYINPUT5), .A3(new_n192), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G113), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n190), .A2(KEYINPUT5), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT84), .A3(G113), .A4(new_n432), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n196), .A2(new_n190), .A3(new_n192), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n389), .A2(new_n368), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n429), .B(new_n430), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n237), .A2(G125), .A3(new_n234), .ZN(new_n442));
  AOI21_X1  g256(.A(G125), .B1(new_n210), .B2(new_n218), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT7), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(KEYINPUT86), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT85), .B(G224), .Z(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G953), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n444), .A2(new_n446), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n445), .ZN(new_n450));
  OAI221_X1 g264(.A(new_n450), .B1(KEYINPUT86), .B2(new_n445), .C1(new_n442), .C2(new_n443), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n441), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n430), .B(KEYINPUT8), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n439), .A2(new_n376), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n438), .B1(new_n433), .B2(new_n434), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n440), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(G902), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n429), .B1(new_n439), .B2(new_n440), .ZN(new_n459));
  INV_X1    g273(.A(new_n430), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT6), .A3(new_n441), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n444), .B(new_n448), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n458), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n458), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n428), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G478), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n350), .A2(new_n290), .A3(G953), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n191), .A2(G122), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n191), .A2(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n358), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n204), .A2(new_n206), .A3(G128), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n216), .A2(G143), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n221), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n475), .A2(new_n476), .A3(G107), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n479), .A2(KEYINPUT92), .A3(new_n484), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n204), .A2(new_n206), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT13), .A3(G128), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n487), .A2(new_n488), .A3(new_n480), .A4(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n483), .B1(new_n491), .B2(G134), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n479), .A2(new_n480), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G134), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n481), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n358), .B1(new_n475), .B2(KEYINPUT14), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n496), .A2(new_n477), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n477), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n474), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n490), .A2(new_n488), .A3(new_n480), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n221), .B1(new_n502), .B2(new_n487), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n501), .B(new_n473), .C1(new_n503), .C2(new_n483), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n472), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n276), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT93), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(KEYINPUT93), .A3(new_n472), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n249), .A2(KEYINPUT87), .A3(G214), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT87), .B1(new_n249), .B2(G214), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n489), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G237), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n332), .A3(G214), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(new_n200), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n225), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n204), .A2(new_n206), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT87), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n525), .B2(new_n514), .ZN(new_n526));
  OAI21_X1  g340(.A(G131), .B1(new_n526), .B2(new_n520), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n225), .B1(new_n517), .B2(new_n521), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n319), .A2(new_n320), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n296), .B(new_n208), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n517), .A2(new_n521), .ZN(new_n535));
  AND2_X1   g349(.A1(KEYINPUT18), .A2(G131), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n537));
  OAI221_X1 g351(.A(new_n534), .B1(new_n535), .B2(new_n536), .C1(new_n537), .C2(new_n527), .ZN(new_n538));
  XOR2_X1   g352(.A(G113), .B(G122), .Z(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT90), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT89), .B(G104), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n533), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n533), .B2(new_n538), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n276), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(new_n276), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(G475), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G475), .A2(G902), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n526), .A2(G131), .A3(new_n520), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n530), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n522), .A2(new_n527), .A3(KEYINPUT88), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n296), .B(KEYINPUT19), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n319), .B1(new_n208), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n542), .B1(new_n558), .B2(new_n538), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n551), .B1(new_n544), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT20), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n551), .C1(new_n544), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n332), .A2(G952), .ZN(new_n565));
  NAND2_X1  g379(.A1(G234), .A2(G237), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(G902), .A3(G953), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT21), .B(G898), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n513), .A2(new_n550), .A3(new_n564), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n470), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n427), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n427), .A2(KEYINPUT94), .A3(new_n575), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n349), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  NOR2_X1   g395(.A1(new_n470), .A2(new_n572), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n509), .B2(new_n471), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n505), .A2(KEYINPUT97), .A3(G478), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n474), .B2(KEYINPUT95), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n500), .A2(new_n504), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n500), .B2(new_n504), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n471), .A2(G902), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT96), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  INV_X1    g409(.A(new_n593), .ZN(new_n596));
  NOR4_X1   g410(.A1(new_n590), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n587), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n550), .A2(new_n564), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT98), .B1(new_n583), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  INV_X1    g416(.A(new_n600), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n582), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n261), .B2(new_n271), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(new_n275), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n272), .ZN(new_n608));
  INV_X1    g422(.A(new_n348), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n427), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n561), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n560), .A2(KEYINPUT100), .A3(KEYINPUT20), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(KEYINPUT99), .A3(new_n563), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n550), .A2(new_n512), .A3(new_n511), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n563), .A2(KEYINPUT99), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n621), .A3(new_n616), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n618), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n583), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n610), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n324), .A2(new_n330), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n294), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n344), .B2(new_n347), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n628), .B1(new_n608), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n633), .ZN(new_n635));
  NOR4_X1   g449(.A1(new_n635), .A2(new_n607), .A3(new_n272), .A4(KEYINPUT101), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n578), .B(new_n579), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT102), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n637), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(new_n427), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n289), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n568), .B1(new_n570), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n618), .A2(new_n620), .A3(new_n622), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n428), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n458), .A2(new_n466), .ZN(new_n648));
  INV_X1    g462(.A(new_n467), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n458), .A2(new_n466), .A3(new_n467), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n633), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n642), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n216), .ZN(G30));
  AOI21_X1  g470(.A(new_n513), .B1(new_n564), .B2(new_n550), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n635), .A2(new_n428), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n273), .A2(new_n279), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n258), .A2(new_n260), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n253), .B1(new_n256), .B2(new_n264), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n276), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT103), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n650), .A2(new_n651), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n659), .A2(new_n666), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n644), .B(KEYINPUT39), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n641), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT40), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n671), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n523), .ZN(G45));
  NAND3_X1  g491(.A1(new_n598), .A2(new_n599), .A3(new_n645), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n653), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n642), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n208), .ZN(G48));
  INV_X1    g495(.A(new_n352), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n426), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n421), .A2(new_n413), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT83), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n422), .A3(new_n423), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n420), .B1(new_n688), .B2(new_n276), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n276), .B1(new_n424), .B2(new_n425), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(KEYINPUT106), .A3(G469), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n682), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n348), .A3(new_n289), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n605), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n624), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n691), .A2(G469), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n683), .A3(new_n426), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n692), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n682), .A3(new_n652), .A4(new_n633), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n288), .A2(G472), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n272), .A2(KEYINPUT70), .A3(new_n187), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT32), .B1(new_n277), .B2(new_n278), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n574), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n701), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g526(.A(new_n352), .B(new_n470), .C1(new_n703), .C2(new_n692), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n574), .B1(new_n660), .B2(new_n706), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n633), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NAND2_X1  g531(.A1(new_n274), .A2(new_n276), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(KEYINPUT108), .A3(G472), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n606), .B2(new_n275), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n652), .A2(new_n573), .A3(new_n657), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n609), .A4(new_n277), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT109), .B1(new_n694), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n352), .B1(new_n703), .B2(new_n692), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n272), .B(new_n348), .C1(new_n719), .C2(new_n721), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n726), .A2(new_n727), .A3(new_n728), .A4(new_n723), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  AOI211_X1 g545(.A(new_n272), .B(new_n678), .C1(new_n719), .C2(new_n721), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n726), .A2(new_n652), .A3(new_n732), .A4(new_n633), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NAND3_X1  g548(.A1(new_n650), .A2(new_n428), .A3(new_n651), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n352), .B(new_n735), .C1(new_n419), .C2(new_n426), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n709), .A2(new_n609), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n272), .A2(KEYINPUT32), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n277), .A2(new_n187), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n706), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n678), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n736), .A3(new_n609), .A4(new_n742), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n737), .A2(new_n738), .B1(new_n743), .B2(KEYINPUT42), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  INV_X1    g559(.A(new_n646), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n709), .A2(new_n609), .A3(new_n746), .A4(new_n736), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  NOR2_X1   g562(.A1(new_n608), .A2(new_n635), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n599), .B(KEYINPUT111), .Z(new_n751));
  INV_X1    g565(.A(new_n598), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n751), .A2(KEYINPUT112), .A3(new_n754), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n753), .B1(new_n752), .B2(new_n599), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT113), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT113), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n750), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT44), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n735), .B1(new_n763), .B2(KEYINPUT44), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n418), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(G469), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n426), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT110), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n774), .B(new_n426), .C1(new_n770), .C2(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n771), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n682), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n673), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n764), .A2(new_n765), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  NOR3_X1   g595(.A1(new_n609), .A2(new_n678), .A3(new_n735), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n777), .A2(KEYINPUT47), .A3(new_n682), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT47), .B1(new_n777), .B2(new_n682), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n289), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n788));
  INV_X1    g602(.A(new_n785), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n704), .B(KEYINPUT115), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n789), .B(new_n783), .C1(new_n682), .C2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n727), .A2(new_n568), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n760), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n735), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n794), .A2(new_n428), .A3(new_n669), .A4(new_n694), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT50), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n735), .A2(new_n567), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n726), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n660), .A2(new_n665), .A3(new_n609), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n800), .A2(KEYINPUT119), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n599), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT119), .B1(new_n800), .B2(new_n801), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n752), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n800), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n272), .B1(new_n719), .B2(new_n721), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n760), .A3(new_n633), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n798), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n788), .B1(new_n796), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n798), .A2(new_n808), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n792), .A2(new_n795), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(KEYINPUT51), .A4(new_n805), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n741), .A2(new_n609), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n806), .A2(new_n760), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT48), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n817));
  INV_X1    g631(.A(new_n713), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n794), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n760), .A2(new_n793), .A3(KEYINPUT120), .A4(new_n713), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n802), .A2(new_n603), .A3(new_n804), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n816), .A2(new_n821), .A3(new_n565), .A4(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT121), .Z(new_n824));
  NAND3_X1  g638(.A1(new_n810), .A2(new_n813), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n709), .B(new_n427), .C1(new_n654), .C2(new_n679), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n652), .A2(new_n657), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n427), .A2(new_n827), .A3(new_n635), .A4(new_n645), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n666), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n733), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n733), .A2(new_n826), .A3(new_n829), .A4(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT117), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n349), .B(new_n726), .C1(new_n605), .C2(new_n624), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n716), .A2(new_n730), .A3(new_n744), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n600), .B1(new_n599), .B2(new_n513), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n610), .A2(new_n582), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n580), .A2(new_n637), .A3(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n550), .A2(new_n618), .A3(new_n513), .A4(new_n622), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n709), .A2(new_n841), .B1(new_n603), .B2(new_n807), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n736), .A2(new_n633), .A3(new_n645), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n747), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n832), .A2(new_n846), .A3(new_n833), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n835), .A2(new_n837), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n716), .A2(new_n730), .A3(new_n744), .A4(new_n836), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n840), .A3(new_n844), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n830), .A2(new_n854), .A3(new_n831), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n833), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT53), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT54), .B1(new_n850), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n849), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n851), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n730), .A2(new_n836), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(KEYINPUT118), .A3(new_n716), .A4(new_n744), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n840), .A2(new_n844), .A3(new_n849), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n856), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n858), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n825), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n791), .A2(KEYINPUT49), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n352), .A2(new_n647), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n609), .A2(new_n751), .A3(new_n598), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n873), .A2(KEYINPUT114), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(KEYINPUT114), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n666), .A4(new_n669), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n877), .B2(new_n790), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n869), .B1(new_n870), .B2(new_n878), .ZN(G75));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n832), .A2(new_n846), .A3(new_n833), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n846), .B1(new_n832), .B2(new_n833), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n883), .B2(new_n852), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n856), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n885));
  OAI211_X1 g699(.A(G210), .B(G902), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n462), .A2(new_n464), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(new_n465), .Z(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT55), .Z(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(new_n887), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n332), .A2(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n886), .B2(new_n887), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n880), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n887), .ZN(new_n897));
  INV_X1    g711(.A(new_n890), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(KEYINPUT122), .A3(new_n891), .A4(new_n893), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n900), .ZN(G51));
  NAND2_X1  g715(.A1(new_n859), .A2(new_n866), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n867), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n769), .B(KEYINPUT57), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n688), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n276), .B1(new_n859), .B2(new_n866), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(G469), .A3(new_n767), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n892), .B1(new_n906), .B2(new_n908), .ZN(G54));
  NAND3_X1  g723(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n544), .A2(new_n559), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n892), .ZN(G60));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n867), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n852), .A2(new_n856), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n849), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n883), .A2(new_n852), .A3(KEYINPUT53), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n860), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n917), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  INV_X1    g738(.A(new_n592), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n916), .B1(new_n858), .B2(new_n867), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT123), .B1(new_n927), .B2(new_n592), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n903), .A2(new_n867), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n916), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n892), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n926), .A2(new_n928), .A3(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n884), .B2(new_n885), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n339), .A2(new_n340), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n892), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n939));
  AND4_X1   g753(.A1(new_n939), .A2(new_n902), .A3(new_n631), .A4(new_n934), .ZN(new_n940));
  INV_X1    g754(.A(new_n934), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n859), .B2(new_n866), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n942), .B2(new_n631), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT61), .B(new_n938), .C1(new_n940), .C2(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(G66));
  INV_X1    g762(.A(new_n840), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n863), .A2(new_n716), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n332), .ZN(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n447), .B2(new_n571), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT125), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n888), .B1(G898), .B2(new_n332), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  INV_X1    g771(.A(new_n245), .ZN(new_n958));
  INV_X1    g772(.A(new_n247), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n556), .B(KEYINPUT126), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n960), .B(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(G900), .B2(G953), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n779), .A2(new_n827), .A3(new_n814), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n733), .A2(new_n744), .A3(new_n747), .A4(new_n826), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n780), .A2(new_n786), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n967), .B2(G953), .ZN(new_n968));
  INV_X1    g782(.A(new_n735), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n349), .A2(new_n674), .A3(new_n969), .A4(new_n838), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n780), .A2(new_n786), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n676), .A2(new_n733), .A3(new_n826), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  AOI21_X1  g787(.A(G953), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n963), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n968), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n332), .B1(G227), .B2(G900), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n979), .B(new_n968), .C1(new_n974), .C2(new_n975), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G72));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n967), .B2(new_n951), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n262), .A3(new_n281), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n893), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n282), .A2(new_n285), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n987), .B2(new_n661), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n920), .B2(new_n921), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n253), .B1(new_n280), .B2(new_n266), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n971), .A2(new_n950), .A3(new_n973), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n983), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n986), .A2(new_n989), .A3(new_n992), .ZN(G57));
endmodule


