

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(n733), .ZN(n738) );
  NAND2_X1 U551 ( .A1(G8), .A2(n733), .ZN(n830) );
  AND2_X1 U552 ( .A1(n525), .A2(n516), .ZN(n839) );
  NAND2_X1 U553 ( .A1(n519), .A2(n518), .ZN(n517) );
  AND2_X1 U554 ( .A1(n523), .A2(n521), .ZN(n520) );
  NOR2_X1 U555 ( .A1(n780), .A2(n779), .ZN(n825) );
  AND2_X1 U556 ( .A1(n750), .A2(n730), .ZN(n731) );
  OR2_X1 U557 ( .A1(n548), .A2(n547), .ZN(n539) );
  INV_X1 U558 ( .A(KEYINPUT103), .ZN(n518) );
  INV_X1 U559 ( .A(G168), .ZN(n529) );
  NAND2_X1 U560 ( .A1(n535), .A2(n534), .ZN(n794) );
  NAND2_X1 U561 ( .A1(n546), .A2(n540), .ZN(n534) );
  AND2_X1 U562 ( .A1(n537), .A2(n536), .ZN(n535) );
  XNOR2_X1 U563 ( .A(n527), .B(n526), .ZN(n727) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n526) );
  NAND2_X1 U565 ( .A1(n528), .A2(n514), .ZN(n527) );
  INV_X1 U566 ( .A(G1384), .ZN(n543) );
  AND2_X1 U567 ( .A1(n543), .A2(KEYINPUT64), .ZN(n541) );
  AND2_X1 U568 ( .A1(n1013), .A2(KEYINPUT103), .ZN(n524) );
  AND2_X1 U569 ( .A1(n515), .A2(n522), .ZN(n521) );
  OR2_X1 U570 ( .A1(n1013), .A2(KEYINPUT103), .ZN(n522) );
  NOR2_X1 U571 ( .A1(n556), .A2(KEYINPUT88), .ZN(n547) );
  NOR2_X1 U572 ( .A1(n557), .A2(KEYINPUT88), .ZN(n548) );
  NAND2_X1 U573 ( .A1(n533), .A2(n553), .ZN(n532) );
  INV_X1 U574 ( .A(G2104), .ZN(n533) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n919) );
  OR2_X1 U576 ( .A1(n757), .A2(G171), .ZN(n514) );
  NOR2_X1 U577 ( .A1(n830), .A2(n821), .ZN(n515) );
  NAND2_X1 U578 ( .A1(n822), .A2(KEYINPUT33), .ZN(n516) );
  NAND2_X1 U579 ( .A1(n520), .A2(n517), .ZN(n525) );
  INV_X1 U580 ( .A(n783), .ZN(n519) );
  NAND2_X1 U581 ( .A1(n783), .A2(n524), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n724), .B(n531), .ZN(n530) );
  INV_X1 U584 ( .A(KEYINPUT100), .ZN(n531) );
  XNOR2_X2 U585 ( .A(n532), .B(KEYINPUT17), .ZN(n913) );
  INV_X1 U586 ( .A(n539), .ZN(n546) );
  NAND2_X1 U587 ( .A1(n542), .A2(n538), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n539), .A2(n538), .ZN(n537) );
  INV_X1 U589 ( .A(KEYINPUT64), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n546), .A2(n544), .ZN(G164) );
  AND2_X1 U591 ( .A1(n544), .A2(n541), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n544), .A2(n543), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n557), .A2(n545), .ZN(n544) );
  AND2_X1 U594 ( .A1(n556), .A2(KEYINPUT88), .ZN(n545) );
  INV_X1 U595 ( .A(KEYINPUT29), .ZN(n755) );
  XNOR2_X1 U596 ( .A(n756), .B(n755), .ZN(n759) );
  INV_X1 U597 ( .A(KEYINPUT99), .ZN(n760) );
  XNOR2_X1 U598 ( .A(KEYINPUT73), .B(KEYINPUT14), .ZN(n624) );
  XNOR2_X1 U599 ( .A(n625), .B(n624), .ZN(n626) );
  INV_X1 U600 ( .A(KEYINPUT87), .ZN(n551) );
  AND2_X1 U601 ( .A1(n553), .A2(G2104), .ZN(n915) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n561), .Z(n690) );
  AND2_X1 U603 ( .A1(G138), .A2(n913), .ZN(n550) );
  AND2_X1 U604 ( .A1(G114), .A2(n919), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n557) );
  INV_X1 U606 ( .A(G2105), .ZN(n553) );
  NOR2_X1 U607 ( .A1(G2104), .A2(n553), .ZN(n578) );
  AND2_X1 U608 ( .A1(n578), .A2(G126), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(n551), .ZN(n555) );
  AND2_X1 U610 ( .A1(n915), .A2(G102), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U612 ( .A1(G651), .A2(G543), .ZN(n677) );
  NAND2_X1 U613 ( .A1(G85), .A2(n677), .ZN(n559) );
  XOR2_X1 U614 ( .A(KEYINPUT0), .B(G543), .Z(n687) );
  INV_X1 U615 ( .A(G651), .ZN(n560) );
  NOR2_X1 U616 ( .A1(n687), .A2(n560), .ZN(n673) );
  NAND2_X1 U617 ( .A1(G72), .A2(n673), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n565) );
  NOR2_X1 U619 ( .A1(G543), .A2(n560), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G60), .A2(n690), .ZN(n563) );
  NOR2_X1 U621 ( .A1(G651), .A2(n687), .ZN(n683) );
  NAND2_X1 U622 ( .A1(G47), .A2(n683), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  OR2_X1 U624 ( .A1(n565), .A2(n564), .ZN(G290) );
  XOR2_X1 U625 ( .A(G2443), .B(KEYINPUT110), .Z(n567) );
  XNOR2_X1 U626 ( .A(G2451), .B(G2427), .ZN(n566) );
  XNOR2_X1 U627 ( .A(n567), .B(n566), .ZN(n571) );
  XOR2_X1 U628 ( .A(G2435), .B(G2438), .Z(n569) );
  XNOR2_X1 U629 ( .A(G2454), .B(G2430), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U631 ( .A(n571), .B(n570), .Z(n573) );
  XNOR2_X1 U632 ( .A(G2446), .B(KEYINPUT108), .ZN(n572) );
  XNOR2_X1 U633 ( .A(n573), .B(n572), .ZN(n576) );
  XOR2_X1 U634 ( .A(G1348), .B(G1341), .Z(n574) );
  XNOR2_X1 U635 ( .A(KEYINPUT109), .B(n574), .ZN(n575) );
  XOR2_X1 U636 ( .A(n576), .B(n575), .Z(n577) );
  AND2_X1 U637 ( .A1(G14), .A2(n577), .ZN(G401) );
  BUF_X1 U638 ( .A(n578), .Z(n922) );
  NAND2_X1 U639 ( .A1(G123), .A2(n922), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT18), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n919), .A2(G111), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G99), .A2(n915), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G135), .A2(n913), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U646 ( .A1(n585), .A2(n584), .ZN(n938) );
  XNOR2_X1 U647 ( .A(n938), .B(G2096), .ZN(n586) );
  XNOR2_X1 U648 ( .A(n586), .B(KEYINPUT79), .ZN(n587) );
  OR2_X1 U649 ( .A1(G2100), .A2(n587), .ZN(G156) );
  INV_X1 U650 ( .A(G57), .ZN(G237) );
  INV_X1 U651 ( .A(G132), .ZN(G219) );
  NAND2_X1 U652 ( .A1(G101), .A2(n915), .ZN(n588) );
  XOR2_X1 U653 ( .A(KEYINPUT23), .B(n588), .Z(n591) );
  NAND2_X1 U654 ( .A1(G113), .A2(n919), .ZN(n589) );
  XOR2_X1 U655 ( .A(KEYINPUT65), .B(n589), .Z(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U657 ( .A1(G125), .A2(n922), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n913), .A2(G137), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(G160) );
  NAND2_X1 U661 ( .A1(n683), .A2(G51), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n596), .B(KEYINPUT78), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G63), .A2(n690), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U665 ( .A(KEYINPUT6), .B(n599), .ZN(n607) );
  NAND2_X1 U666 ( .A1(G89), .A2(n677), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT4), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT76), .ZN(n603) );
  NAND2_X1 U669 ( .A1(G76), .A2(n673), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U671 ( .A(KEYINPUT77), .B(n604), .ZN(n605) );
  XNOR2_X1 U672 ( .A(KEYINPUT5), .B(n605), .ZN(n606) );
  NOR2_X1 U673 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U674 ( .A(KEYINPUT7), .B(n608), .Z(G168) );
  XOR2_X1 U675 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U676 ( .A1(G65), .A2(n690), .ZN(n610) );
  NAND2_X1 U677 ( .A1(G53), .A2(n683), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U679 ( .A(KEYINPUT70), .B(n611), .Z(n615) );
  NAND2_X1 U680 ( .A1(G91), .A2(n677), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G78), .A2(n673), .ZN(n612) );
  AND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(G299) );
  NAND2_X1 U684 ( .A1(G94), .A2(G452), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n616), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U686 ( .A1(G7), .A2(G661), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(KEYINPUT10), .ZN(n618) );
  XNOR2_X1 U688 ( .A(KEYINPUT72), .B(n618), .ZN(G223) );
  INV_X1 U689 ( .A(G223), .ZN(n859) );
  NAND2_X1 U690 ( .A1(n859), .A2(G567), .ZN(n619) );
  XOR2_X1 U691 ( .A(KEYINPUT11), .B(n619), .Z(G234) );
  NAND2_X1 U692 ( .A1(n677), .A2(G81), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n620), .B(KEYINPUT12), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G68), .A2(n673), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U696 ( .A(KEYINPUT13), .B(n623), .Z(n627) );
  NAND2_X1 U697 ( .A1(G56), .A2(n690), .ZN(n625) );
  NOR2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U699 ( .A(n628), .B(KEYINPUT74), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G43), .A2(n683), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n1024) );
  INV_X1 U702 ( .A(G860), .ZN(n653) );
  OR2_X1 U703 ( .A1(n1024), .A2(n653), .ZN(G153) );
  NAND2_X1 U704 ( .A1(n690), .A2(G64), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n631), .B(KEYINPUT66), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G52), .A2(n683), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U708 ( .A(KEYINPUT67), .B(n634), .Z(n639) );
  NAND2_X1 U709 ( .A1(G90), .A2(n677), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G77), .A2(n673), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U712 ( .A(KEYINPUT9), .B(n637), .Z(n638) );
  NOR2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U714 ( .A(KEYINPUT68), .B(n640), .ZN(G171) );
  XNOR2_X1 U715 ( .A(KEYINPUT75), .B(G171), .ZN(G301) );
  NAND2_X1 U716 ( .A1(G868), .A2(G301), .ZN(n649) );
  NAND2_X1 U717 ( .A1(G92), .A2(n677), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G79), .A2(n673), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G66), .A2(n690), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G54), .A2(n683), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT15), .B(n647), .Z(n1012) );
  INV_X1 U725 ( .A(n1012), .ZN(n884) );
  INV_X1 U726 ( .A(G868), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n884), .A2(n650), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(G284) );
  NOR2_X1 U729 ( .A1(G286), .A2(n650), .ZN(n652) );
  NOR2_X1 U730 ( .A1(G868), .A2(G299), .ZN(n651) );
  NOR2_X1 U731 ( .A1(n652), .A2(n651), .ZN(G297) );
  NAND2_X1 U732 ( .A1(n653), .A2(G559), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n654), .A2(n1012), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n655), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U735 ( .A1(G868), .A2(n1024), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n1012), .A2(G868), .ZN(n656) );
  NOR2_X1 U737 ( .A1(G559), .A2(n656), .ZN(n657) );
  NOR2_X1 U738 ( .A1(n658), .A2(n657), .ZN(G282) );
  NAND2_X1 U739 ( .A1(n1012), .A2(G559), .ZN(n701) );
  XNOR2_X1 U740 ( .A(n1024), .B(n701), .ZN(n659) );
  NOR2_X1 U741 ( .A1(n659), .A2(G860), .ZN(n666) );
  NAND2_X1 U742 ( .A1(G67), .A2(n690), .ZN(n661) );
  NAND2_X1 U743 ( .A1(G55), .A2(n683), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G93), .A2(n677), .ZN(n663) );
  NAND2_X1 U746 ( .A1(G80), .A2(n673), .ZN(n662) );
  NAND2_X1 U747 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U748 ( .A1(n665), .A2(n664), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n666), .B(n695), .ZN(G145) );
  NAND2_X1 U750 ( .A1(G88), .A2(n677), .ZN(n668) );
  NAND2_X1 U751 ( .A1(G75), .A2(n673), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G62), .A2(n690), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G50), .A2(n683), .ZN(n669) );
  NAND2_X1 U755 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U756 ( .A1(n672), .A2(n671), .ZN(G166) );
  INV_X1 U757 ( .A(G166), .ZN(G303) );
  NAND2_X1 U758 ( .A1(G73), .A2(n673), .ZN(n674) );
  XNOR2_X1 U759 ( .A(n674), .B(KEYINPUT2), .ZN(n682) );
  NAND2_X1 U760 ( .A1(G61), .A2(n690), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G48), .A2(n683), .ZN(n675) );
  NAND2_X1 U762 ( .A1(n676), .A2(n675), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n677), .A2(G86), .ZN(n678) );
  XOR2_X1 U764 ( .A(KEYINPUT82), .B(n678), .Z(n679) );
  NOR2_X1 U765 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n682), .A2(n681), .ZN(G305) );
  NAND2_X1 U767 ( .A1(G49), .A2(n683), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G74), .A2(G651), .ZN(n684) );
  NAND2_X1 U769 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U770 ( .A(KEYINPUT80), .B(n686), .Z(n692) );
  NAND2_X1 U771 ( .A1(G87), .A2(n687), .ZN(n688) );
  XNOR2_X1 U772 ( .A(KEYINPUT81), .B(n688), .ZN(n689) );
  NOR2_X1 U773 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U774 ( .A1(n692), .A2(n691), .ZN(G288) );
  NOR2_X1 U775 ( .A1(G868), .A2(n695), .ZN(n693) );
  XNOR2_X1 U776 ( .A(n693), .B(KEYINPUT83), .ZN(n704) );
  XNOR2_X1 U777 ( .A(KEYINPUT19), .B(G303), .ZN(n694) );
  XNOR2_X1 U778 ( .A(n694), .B(G305), .ZN(n698) );
  XNOR2_X1 U779 ( .A(n695), .B(G290), .ZN(n696) );
  XNOR2_X1 U780 ( .A(n696), .B(G299), .ZN(n697) );
  XNOR2_X1 U781 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U782 ( .A(n699), .B(G288), .ZN(n700) );
  XNOR2_X1 U783 ( .A(n1024), .B(n700), .ZN(n886) );
  XNOR2_X1 U784 ( .A(n886), .B(n701), .ZN(n702) );
  NAND2_X1 U785 ( .A1(G868), .A2(n702), .ZN(n703) );
  NAND2_X1 U786 ( .A1(n704), .A2(n703), .ZN(G295) );
  NAND2_X1 U787 ( .A1(G2084), .A2(G2078), .ZN(n705) );
  XOR2_X1 U788 ( .A(KEYINPUT20), .B(n705), .Z(n706) );
  NAND2_X1 U789 ( .A1(G2090), .A2(n706), .ZN(n707) );
  XNOR2_X1 U790 ( .A(KEYINPUT21), .B(n707), .ZN(n708) );
  NAND2_X1 U791 ( .A1(n708), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U792 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U793 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NAND2_X1 U794 ( .A1(G661), .A2(G483), .ZN(n718) );
  NOR2_X1 U795 ( .A1(G219), .A2(G220), .ZN(n709) );
  XOR2_X1 U796 ( .A(KEYINPUT22), .B(n709), .Z(n710) );
  XNOR2_X1 U797 ( .A(n710), .B(KEYINPUT84), .ZN(n711) );
  NOR2_X1 U798 ( .A1(G218), .A2(n711), .ZN(n712) );
  NAND2_X1 U799 ( .A1(G96), .A2(n712), .ZN(n864) );
  NAND2_X1 U800 ( .A1(G2106), .A2(n864), .ZN(n713) );
  XOR2_X1 U801 ( .A(KEYINPUT85), .B(n713), .Z(n717) );
  NAND2_X1 U802 ( .A1(G120), .A2(G69), .ZN(n714) );
  NOR2_X1 U803 ( .A1(G237), .A2(n714), .ZN(n715) );
  NAND2_X1 U804 ( .A1(G108), .A2(n715), .ZN(n863) );
  NAND2_X1 U805 ( .A1(G567), .A2(n863), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n866) );
  NOR2_X1 U807 ( .A1(n718), .A2(n866), .ZN(n719) );
  XNOR2_X1 U808 ( .A(n719), .B(KEYINPUT86), .ZN(n862) );
  NAND2_X1 U809 ( .A1(G36), .A2(n862), .ZN(G176) );
  NOR2_X1 U810 ( .A1(G1971), .A2(G303), .ZN(n720) );
  XOR2_X1 U811 ( .A(n720), .B(KEYINPUT102), .Z(n782) );
  NOR2_X1 U812 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  NAND2_X1 U813 ( .A1(G160), .A2(G40), .ZN(n795) );
  INV_X1 U814 ( .A(n795), .ZN(n721) );
  NAND2_X2 U815 ( .A1(n721), .A2(n794), .ZN(n733) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n830), .ZN(n778) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n733), .ZN(n773) );
  NOR2_X1 U818 ( .A1(n778), .A2(n773), .ZN(n722) );
  NAND2_X1 U819 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  XNOR2_X1 U821 ( .A(G2078), .B(KEYINPUT25), .ZN(n963) );
  NOR2_X1 U822 ( .A1(n733), .A2(n963), .ZN(n726) );
  INV_X1 U823 ( .A(G1961), .ZN(n984) );
  NOR2_X1 U824 ( .A1(n738), .A2(n984), .ZN(n725) );
  NOR2_X1 U825 ( .A1(n726), .A2(n725), .ZN(n757) );
  XNOR2_X1 U826 ( .A(n727), .B(KEYINPUT101), .ZN(n763) );
  AND2_X1 U827 ( .A1(n738), .A2(G2072), .ZN(n728) );
  XNOR2_X1 U828 ( .A(KEYINPUT27), .B(n728), .ZN(n750) );
  NAND2_X1 U829 ( .A1(G1956), .A2(n733), .ZN(n749) );
  INV_X1 U830 ( .A(G299), .ZN(n729) );
  AND2_X1 U831 ( .A1(n749), .A2(n729), .ZN(n730) );
  XOR2_X1 U832 ( .A(KEYINPUT98), .B(n731), .Z(n748) );
  XOR2_X1 U833 ( .A(G1996), .B(KEYINPUT95), .Z(n964) );
  NAND2_X1 U834 ( .A1(n738), .A2(n964), .ZN(n732) );
  XNOR2_X1 U835 ( .A(n732), .B(KEYINPUT26), .ZN(n736) );
  NAND2_X1 U836 ( .A1(n733), .A2(G1341), .ZN(n734) );
  XNOR2_X1 U837 ( .A(n734), .B(KEYINPUT96), .ZN(n735) );
  NAND2_X1 U838 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U839 ( .A1(n1024), .A2(n737), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n744), .A2(n1012), .ZN(n743) );
  AND2_X1 U841 ( .A1(n738), .A2(G2067), .ZN(n739) );
  XNOR2_X1 U842 ( .A(n739), .B(KEYINPUT97), .ZN(n741) );
  NAND2_X1 U843 ( .A1(n733), .A2(G1348), .ZN(n740) );
  NAND2_X1 U844 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U845 ( .A1(n743), .A2(n742), .ZN(n746) );
  OR2_X1 U846 ( .A1(n1012), .A2(n744), .ZN(n745) );
  NAND2_X1 U847 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U848 ( .A1(n748), .A2(n747), .ZN(n754) );
  NAND2_X1 U849 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U850 ( .A1(G299), .A2(n751), .ZN(n752) );
  XNOR2_X1 U851 ( .A(n752), .B(KEYINPUT28), .ZN(n753) );
  NAND2_X1 U852 ( .A1(n754), .A2(n753), .ZN(n756) );
  NAND2_X1 U853 ( .A1(n757), .A2(G171), .ZN(n758) );
  NAND2_X1 U854 ( .A1(n759), .A2(n758), .ZN(n761) );
  XNOR2_X1 U855 ( .A(n761), .B(n760), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n763), .A2(n762), .ZN(n775) );
  AND2_X1 U857 ( .A1(G286), .A2(G8), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n775), .A2(n764), .ZN(n771) );
  INV_X1 U859 ( .A(G8), .ZN(n769) );
  NOR2_X1 U860 ( .A1(G1971), .A2(n830), .ZN(n766) );
  NOR2_X1 U861 ( .A1(G2090), .A2(n733), .ZN(n765) );
  NOR2_X1 U862 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n767), .A2(G303), .ZN(n768) );
  OR2_X1 U864 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U866 ( .A(n772), .B(KEYINPUT32), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G8), .A2(n773), .ZN(n774) );
  XNOR2_X1 U868 ( .A(KEYINPUT94), .B(n774), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U871 ( .A1(n1011), .A2(n825), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  XOR2_X1 U874 ( .A(G1981), .B(G305), .Z(n1007) );
  NAND2_X1 U875 ( .A1(G104), .A2(n915), .ZN(n785) );
  NAND2_X1 U876 ( .A1(G140), .A2(n913), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G116), .A2(n919), .ZN(n788) );
  NAND2_X1 U880 ( .A1(G128), .A2(n922), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U882 ( .A(n789), .B(KEYINPUT35), .Z(n790) );
  NOR2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT36), .B(n792), .Z(n793) );
  XOR2_X1 U885 ( .A(KEYINPUT90), .B(n793), .Z(n929) );
  XNOR2_X1 U886 ( .A(G2067), .B(KEYINPUT37), .ZN(n850) );
  NOR2_X1 U887 ( .A1(n929), .A2(n850), .ZN(n941) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n841) );
  NAND2_X1 U889 ( .A1(n941), .A2(n841), .ZN(n796) );
  XNOR2_X1 U890 ( .A(n796), .B(KEYINPUT91), .ZN(n849) );
  INV_X1 U891 ( .A(n849), .ZN(n797) );
  AND2_X1 U892 ( .A1(n1007), .A2(n797), .ZN(n799) );
  XOR2_X1 U893 ( .A(G1986), .B(KEYINPUT89), .Z(n798) );
  XNOR2_X1 U894 ( .A(G290), .B(n798), .ZN(n1021) );
  NAND2_X1 U895 ( .A1(n841), .A2(n1021), .ZN(n834) );
  AND2_X1 U896 ( .A1(n799), .A2(n834), .ZN(n817) );
  NAND2_X1 U897 ( .A1(G129), .A2(n922), .ZN(n801) );
  NAND2_X1 U898 ( .A1(G141), .A2(n913), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n915), .A2(G105), .ZN(n802) );
  XOR2_X1 U901 ( .A(KEYINPUT38), .B(n802), .Z(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n919), .A2(G117), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n910) );
  NAND2_X1 U905 ( .A1(G1996), .A2(n910), .ZN(n814) );
  NAND2_X1 U906 ( .A1(G119), .A2(n922), .ZN(n808) );
  NAND2_X1 U907 ( .A1(G131), .A2(n913), .ZN(n807) );
  NAND2_X1 U908 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U909 ( .A1(G107), .A2(n919), .ZN(n810) );
  NAND2_X1 U910 ( .A1(G95), .A2(n915), .ZN(n809) );
  NAND2_X1 U911 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U912 ( .A1(n812), .A2(n811), .ZN(n897) );
  NAND2_X1 U913 ( .A1(G1991), .A2(n897), .ZN(n813) );
  NAND2_X1 U914 ( .A1(n814), .A2(n813), .ZN(n945) );
  NAND2_X1 U915 ( .A1(n945), .A2(n841), .ZN(n815) );
  XOR2_X1 U916 ( .A(KEYINPUT92), .B(n815), .Z(n844) );
  INV_X1 U917 ( .A(n844), .ZN(n816) );
  NAND2_X1 U918 ( .A1(n817), .A2(n816), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n1011), .A2(KEYINPUT33), .ZN(n818) );
  NOR2_X1 U920 ( .A1(n818), .A2(n830), .ZN(n819) );
  OR2_X1 U921 ( .A1(n820), .A2(n819), .ZN(n821) );
  INV_X1 U922 ( .A(n821), .ZN(n822) );
  NOR2_X1 U923 ( .A1(G2090), .A2(G303), .ZN(n823) );
  AND2_X1 U924 ( .A1(G8), .A2(n823), .ZN(n824) );
  OR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U926 ( .A1(n826), .A2(n830), .ZN(n832) );
  NOR2_X1 U927 ( .A1(G1981), .A2(G305), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n827), .B(KEYINPUT24), .ZN(n828) );
  XNOR2_X1 U929 ( .A(KEYINPUT93), .B(n828), .ZN(n829) );
  OR2_X1 U930 ( .A1(n830), .A2(n829), .ZN(n831) );
  AND2_X1 U931 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U932 ( .A1(n849), .A2(n833), .ZN(n837) );
  INV_X1 U933 ( .A(n834), .ZN(n835) );
  NOR2_X1 U934 ( .A1(n835), .A2(n844), .ZN(n836) );
  NAND2_X1 U935 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U937 ( .A(KEYINPUT104), .B(n840), .Z(n857) );
  INV_X1 U938 ( .A(n841), .ZN(n854) );
  NOR2_X1 U939 ( .A1(G1996), .A2(n910), .ZN(n952) );
  NOR2_X1 U940 ( .A1(G1986), .A2(G290), .ZN(n842) );
  NOR2_X1 U941 ( .A1(G1991), .A2(n897), .ZN(n939) );
  NOR2_X1 U942 ( .A1(n842), .A2(n939), .ZN(n843) );
  NOR2_X1 U943 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U944 ( .A1(n952), .A2(n845), .ZN(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT39), .B(n846), .ZN(n847) );
  XNOR2_X1 U946 ( .A(KEYINPUT105), .B(n847), .ZN(n848) );
  NOR2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n852) );
  AND2_X1 U948 ( .A1(n929), .A2(n850), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n851), .B(KEYINPUT106), .ZN(n959) );
  NOR2_X1 U950 ( .A1(n852), .A2(n959), .ZN(n853) );
  NOR2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U952 ( .A(KEYINPUT107), .B(n855), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U954 ( .A(KEYINPUT40), .B(n858), .ZN(G329) );
  NAND2_X1 U955 ( .A1(G2106), .A2(n859), .ZN(G217) );
  AND2_X1 U956 ( .A1(G15), .A2(G2), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G661), .A2(n860), .ZN(G259) );
  NAND2_X1 U958 ( .A1(G3), .A2(G1), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(G188) );
  XNOR2_X1 U960 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U962 ( .A(G120), .ZN(G236) );
  NOR2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n865), .B(KEYINPUT112), .ZN(G325) );
  INV_X1 U965 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U966 ( .A(KEYINPUT113), .B(n866), .ZN(G319) );
  XOR2_X1 U967 ( .A(G2100), .B(G2096), .Z(n868) );
  XNOR2_X1 U968 ( .A(KEYINPUT42), .B(G2678), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT43), .B(G2090), .Z(n870) );
  XNOR2_X1 U971 ( .A(G2067), .B(G2072), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(n872), .B(n871), .Z(n874) );
  XNOR2_X1 U974 ( .A(G2084), .B(G2078), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(G227) );
  XOR2_X1 U976 ( .A(G1976), .B(G1981), .Z(n876) );
  XNOR2_X1 U977 ( .A(G1986), .B(G1961), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U979 ( .A(n877), .B(G2474), .Z(n879) );
  XNOR2_X1 U980 ( .A(G1966), .B(G1971), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT41), .B(G1956), .Z(n881) );
  XNOR2_X1 U983 ( .A(G1996), .B(G1991), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(G229) );
  XNOR2_X1 U986 ( .A(G286), .B(G171), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U989 ( .A1(G37), .A2(n888), .ZN(G397) );
  NAND2_X1 U990 ( .A1(n922), .A2(G124), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n889), .B(KEYINPUT44), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G136), .A2(n913), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U994 ( .A(KEYINPUT114), .B(n892), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G112), .A2(n919), .ZN(n894) );
  NAND2_X1 U996 ( .A1(G100), .A2(n915), .ZN(n893) );
  NAND2_X1 U997 ( .A1(n894), .A2(n893), .ZN(n895) );
  NOR2_X1 U998 ( .A1(n896), .A2(n895), .ZN(G162) );
  XNOR2_X1 U999 ( .A(G162), .B(G164), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1001 ( .A(n899), .B(KEYINPUT48), .Z(n901) );
  XNOR2_X1 U1002 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n900) );
  XNOR2_X1 U1003 ( .A(n901), .B(n900), .ZN(n912) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n915), .ZN(n903) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n913), .ZN(n902) );
  NAND2_X1 U1006 ( .A1(n903), .A2(n902), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(G115), .A2(n919), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(G127), .A2(n922), .ZN(n904) );
  NAND2_X1 U1009 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1010 ( .A(KEYINPUT47), .B(n906), .Z(n907) );
  NOR2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n946) );
  XOR2_X1 U1012 ( .A(n946), .B(n938), .Z(n909) );
  XNOR2_X1 U1013 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1014 ( .A(n912), .B(n911), .Z(n928) );
  NAND2_X1 U1015 ( .A1(n913), .A2(G142), .ZN(n914) );
  XNOR2_X1 U1016 ( .A(n914), .B(KEYINPUT116), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(G106), .A2(n915), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT45), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(G118), .A2(n919), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(G130), .A2(n922), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(KEYINPUT115), .B(n923), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(G160), .B(n926), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(G37), .A2(n931), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(KEYINPUT118), .B(n932), .ZN(G395) );
  NOR2_X1 U1030 ( .A1(G227), .A2(G229), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT49), .B(n933), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(G401), .A2(n934), .ZN(n935) );
  AND2_X1 U1033 ( .A1(G319), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(G397), .A2(G395), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(G225) );
  INV_X1 U1036 ( .A(G225), .ZN(G308) );
  INV_X1 U1037 ( .A(G108), .ZN(G238) );
  INV_X1 U1038 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1039 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1045) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n1036) );
  NOR2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n943) );
  XOR2_X1 U1042 ( .A(G160), .B(G2084), .Z(n940) );
  NOR2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n957) );
  XNOR2_X1 U1046 ( .A(G2072), .B(n946), .ZN(n949) );
  XOR2_X1 U1047 ( .A(G2078), .B(KEYINPUT119), .Z(n947) );
  XNOR2_X1 U1048 ( .A(G164), .B(n947), .ZN(n948) );
  NAND2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(n950), .B(KEYINPUT50), .ZN(n955) );
  XOR2_X1 U1051 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1053 ( .A(KEYINPUT51), .B(n953), .ZN(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(KEYINPUT52), .B(n960), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n1036), .A2(n961), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n962), .A2(G29), .ZN(n1043) );
  XNOR2_X1 U1060 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n976) );
  XOR2_X1 U1061 ( .A(n963), .B(G27), .Z(n966) );
  XNOR2_X1 U1062 ( .A(n964), .B(G32), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT120), .B(n967), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(G33), .B(G2072), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1069 ( .A(G1991), .B(G25), .Z(n972) );
  NAND2_X1 U1070 ( .A1(G28), .A2(n972), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(n976), .B(n975), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G2084), .B(G34), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(n977), .B(KEYINPUT54), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(G35), .B(G2090), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n1037) );
  NOR2_X1 U1078 ( .A1(G29), .A2(KEYINPUT55), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n1037), .A2(n982), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(G11), .A2(n983), .ZN(n1041) );
  XNOR2_X1 U1081 ( .A(G5), .B(n984), .ZN(n1002) );
  XNOR2_X1 U1082 ( .A(KEYINPUT59), .B(G4), .ZN(n985) );
  XNOR2_X1 U1083 ( .A(n985), .B(KEYINPUT125), .ZN(n986) );
  XNOR2_X1 U1084 ( .A(G1348), .B(n986), .ZN(n988) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n987) );
  NOR2_X1 U1086 ( .A1(n988), .A2(n987), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n990) );
  XNOR2_X1 U1088 ( .A(G1956), .B(G20), .ZN(n989) );
  NOR2_X1 U1089 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1090 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1091 ( .A(n993), .B(KEYINPUT60), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n995) );
  XNOR2_X1 U1093 ( .A(G23), .B(G1976), .ZN(n994) );
  NOR2_X1 U1094 ( .A1(n995), .A2(n994), .ZN(n997) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n996) );
  NAND2_X1 U1096 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n998), .ZN(n999) );
  NOR2_X1 U1098 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1099 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1003) );
  NOR2_X1 U1101 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1005), .Z(n1006) );
  NOR2_X1 U1103 ( .A1(G16), .A2(n1006), .ZN(n1034) );
  XOR2_X1 U1104 ( .A(G16), .B(KEYINPUT56), .Z(n1031) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G168), .ZN(n1008) );
  NAND2_X1 U1106 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1107 ( .A(n1009), .B(KEYINPUT57), .ZN(n1028) );
  XNOR2_X1 U1108 ( .A(G1961), .B(G171), .ZN(n1023) );
  XOR2_X1 U1109 ( .A(G1971), .B(G166), .Z(n1010) );
  NOR2_X1 U1110 ( .A1(n1011), .A2(n1010), .ZN(n1019) );
  XNOR2_X1 U1111 ( .A(G1348), .B(n1012), .ZN(n1014) );
  NAND2_X1 U1112 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1113 ( .A(G1956), .B(G299), .ZN(n1015) );
  XNOR2_X1 U1114 ( .A(KEYINPUT122), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1115 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1116 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1117 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1118 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XNOR2_X1 U1119 ( .A(G1341), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1120 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1121 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1122 ( .A(n1029), .B(KEYINPUT123), .ZN(n1030) );
  NOR2_X1 U1123 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1124 ( .A(n1032), .B(KEYINPUT124), .ZN(n1033) );
  NOR2_X1 U1125 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1126 ( .A(KEYINPUT126), .B(n1035), .ZN(n1039) );
  OR2_X1 U1127 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1128 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1129 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1130 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XNOR2_X1 U1131 ( .A(n1045), .B(n1044), .ZN(G311) );
  INV_X1 U1132 ( .A(G311), .ZN(G150) );
endmodule

