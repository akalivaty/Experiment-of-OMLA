

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575;

  XNOR2_X1 U321 ( .A(n340), .B(n307), .ZN(n308) );
  AND2_X1 U322 ( .A1(n445), .A2(n454), .ZN(n556) );
  XNOR2_X1 U323 ( .A(n427), .B(n289), .ZN(n445) );
  XNOR2_X1 U324 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U325 ( .A(n361), .B(n566), .ZN(n542) );
  XNOR2_X1 U326 ( .A(KEYINPUT124), .B(KEYINPUT55), .ZN(n289) );
  XOR2_X1 U327 ( .A(KEYINPUT75), .B(KEYINPUT13), .Z(n290) );
  XOR2_X1 U328 ( .A(G92GAT), .B(G218GAT), .Z(n291) );
  INV_X1 U329 ( .A(KEYINPUT76), .ZN(n349) );
  XNOR2_X1 U330 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U331 ( .A(n352), .B(n351), .ZN(n360) );
  XOR2_X1 U332 ( .A(KEYINPUT36), .B(n533), .Z(n573) );
  XOR2_X1 U333 ( .A(KEYINPUT82), .B(n551), .Z(n533) );
  XOR2_X1 U334 ( .A(n468), .B(KEYINPUT28), .Z(n523) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n446) );
  XNOR2_X1 U336 ( .A(n447), .B(n446), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(G50GAT), .B(KEYINPUT78), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n292), .B(G162GAT), .ZN(n424) );
  XNOR2_X1 U339 ( .A(G99GAT), .B(G106GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n293), .B(G85GAT), .ZN(n348) );
  XNOR2_X1 U341 ( .A(n424), .B(n348), .ZN(n311) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n291), .B(n294), .ZN(n382) );
  XOR2_X1 U344 ( .A(KEYINPUT79), .B(n382), .Z(n296) );
  NAND2_X1 U345 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n309) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(KEYINPUT73), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n297), .B(G29GAT), .ZN(n298) );
  XOR2_X1 U349 ( .A(n298), .B(KEYINPUT7), .Z(n300) );
  XNOR2_X1 U350 ( .A(KEYINPUT8), .B(KEYINPUT74), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n340) );
  XOR2_X1 U352 ( .A(KEYINPUT66), .B(KEYINPUT80), .Z(n302) );
  XNOR2_X1 U353 ( .A(KEYINPUT9), .B(KEYINPUT81), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U355 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n304) );
  XNOR2_X1 U356 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(n306), .B(n305), .Z(n307) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n551) );
  XNOR2_X1 U360 ( .A(G22GAT), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n312), .B(G78GAT), .ZN(n416) );
  XNOR2_X1 U362 ( .A(G71GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n290), .B(n313), .ZN(n345) );
  XNOR2_X1 U364 ( .A(n416), .B(n345), .ZN(n328) );
  XOR2_X1 U365 ( .A(KEYINPUT83), .B(G211GAT), .Z(n315) );
  XNOR2_X1 U366 ( .A(G8GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n378) );
  XOR2_X1 U368 ( .A(n378), .B(G64GAT), .Z(n317) );
  XOR2_X1 U369 ( .A(G15GAT), .B(G127GAT), .Z(n428) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(n428), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U372 ( .A(KEYINPUT12), .B(KEYINPUT85), .Z(n319) );
  NAND2_X1 U373 ( .A1(G231GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U375 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U376 ( .A(KEYINPUT86), .B(KEYINPUT15), .Z(n323) );
  XNOR2_X1 U377 ( .A(KEYINPUT14), .B(KEYINPUT84), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n324), .B(KEYINPUT87), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U381 ( .A(n328), .B(n327), .Z(n570) );
  XOR2_X1 U382 ( .A(n570), .B(KEYINPUT114), .Z(n557) );
  XOR2_X1 U383 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n363) );
  XOR2_X1 U384 ( .A(KEYINPUT29), .B(KEYINPUT71), .Z(n330) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(KEYINPUT70), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n344) );
  XOR2_X1 U387 ( .A(G15GAT), .B(G197GAT), .Z(n332) );
  XNOR2_X1 U388 ( .A(G141GAT), .B(G22GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U390 ( .A(n333), .B(G50GAT), .Z(n335) );
  XOR2_X1 U391 ( .A(G113GAT), .B(G1GAT), .Z(n390) );
  XNOR2_X1 U392 ( .A(n390), .B(G36GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U394 ( .A(KEYINPUT72), .B(G8GAT), .Z(n337) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U397 ( .A(n339), .B(n338), .Z(n342) );
  XNOR2_X1 U398 ( .A(n340), .B(KEYINPUT30), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(n344), .B(n343), .Z(n563) );
  INV_X1 U401 ( .A(n563), .ZN(n553) );
  XNOR2_X1 U402 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n361) );
  XOR2_X1 U403 ( .A(G176GAT), .B(G64GAT), .Z(n375) );
  XOR2_X1 U404 ( .A(n375), .B(n345), .Z(n347) );
  NAND2_X1 U405 ( .A1(G230GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n348), .B(KEYINPUT31), .ZN(n350) );
  XOR2_X1 U408 ( .A(G92GAT), .B(G204GAT), .Z(n354) );
  XNOR2_X1 U409 ( .A(G148GAT), .B(G78GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U411 ( .A(KEYINPUT33), .B(KEYINPUT77), .Z(n356) );
  XNOR2_X1 U412 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U414 ( .A(n358), .B(n357), .Z(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n566) );
  NAND2_X1 U416 ( .A1(n553), .A2(n542), .ZN(n362) );
  XOR2_X1 U417 ( .A(n363), .B(n362), .Z(n364) );
  NOR2_X1 U418 ( .A1(n557), .A2(n364), .ZN(n365) );
  NAND2_X1 U419 ( .A1(n551), .A2(n365), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n366), .B(KEYINPUT47), .ZN(n371) );
  NOR2_X1 U421 ( .A1(n573), .A2(n570), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n367), .B(KEYINPUT45), .ZN(n368) );
  NAND2_X1 U423 ( .A1(n368), .A2(n566), .ZN(n369) );
  NOR2_X1 U424 ( .A1(n553), .A2(n369), .ZN(n370) );
  NOR2_X1 U425 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n372), .B(KEYINPUT48), .ZN(n521) );
  XOR2_X1 U427 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n374) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n429) );
  XOR2_X1 U430 ( .A(KEYINPUT99), .B(n375), .Z(n377) );
  NAND2_X1 U431 ( .A1(G226GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n379) );
  XOR2_X1 U433 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U434 ( .A(G204GAT), .B(KEYINPUT21), .Z(n381) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(KEYINPUT94), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n415) );
  XNOR2_X1 U437 ( .A(n415), .B(n382), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n429), .B(n385), .ZN(n515) );
  XOR2_X1 U440 ( .A(n515), .B(KEYINPUT123), .Z(n386) );
  NOR2_X1 U441 ( .A1(n521), .A2(n386), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n387), .B(KEYINPUT54), .ZN(n410) );
  XOR2_X1 U443 ( .A(G120GAT), .B(KEYINPUT90), .Z(n389) );
  XNOR2_X1 U444 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n432) );
  XOR2_X1 U446 ( .A(n432), .B(n390), .Z(n392) );
  NAND2_X1 U447 ( .A1(G225GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U449 ( .A(n393), .B(KEYINPUT6), .Z(n397) );
  XOR2_X1 U450 ( .A(G148GAT), .B(KEYINPUT3), .Z(n395) );
  XNOR2_X1 U451 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n423) );
  XNOR2_X1 U453 ( .A(n423), .B(KEYINPUT5), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U455 ( .A(G85GAT), .B(G155GAT), .Z(n399) );
  XNOR2_X1 U456 ( .A(G29GAT), .B(G162GAT), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U458 ( .A(n401), .B(n400), .Z(n409) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n403) );
  XNOR2_X1 U460 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n405) );
  XNOR2_X1 U463 ( .A(G127GAT), .B(G57GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n512) );
  NAND2_X1 U467 ( .A1(n410), .A2(n512), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n411), .B(KEYINPUT65), .ZN(n561) );
  XOR2_X1 U469 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n413) );
  NAND2_X1 U470 ( .A1(G228GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U472 ( .A(n414), .B(G211GAT), .Z(n418) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U475 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n420) );
  XNOR2_X1 U476 ( .A(G218GAT), .B(G106GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U478 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n467) );
  NAND2_X1 U481 ( .A1(n561), .A2(n467), .ZN(n427) );
  XOR2_X1 U482 ( .A(n429), .B(n428), .Z(n431) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(G190GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n436) );
  XOR2_X1 U485 ( .A(n432), .B(G113GAT), .Z(n434) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U488 ( .A(n436), .B(n435), .Z(n444) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n438) );
  XNOR2_X1 U490 ( .A(G99GAT), .B(KEYINPUT67), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U492 ( .A(G176GAT), .B(G71GAT), .Z(n440) );
  XNOR2_X1 U493 ( .A(KEYINPUT20), .B(G183GAT), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U496 ( .A(n444), .B(n443), .Z(n454) );
  INV_X1 U497 ( .A(n454), .ZN(n525) );
  NAND2_X1 U498 ( .A1(n556), .A2(n533), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n556), .A2(n542), .ZN(n450) );
  XOR2_X1 U500 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n448) );
  XNOR2_X1 U501 ( .A(n448), .B(G176GAT), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  OR2_X1 U503 ( .A1(n533), .A2(n570), .ZN(n453) );
  XNOR2_X1 U504 ( .A(KEYINPUT16), .B(KEYINPUT89), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n451), .B(KEYINPUT88), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n475) );
  NOR2_X1 U507 ( .A1(n467), .A2(n454), .ZN(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT102), .B(KEYINPUT26), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n562) );
  XOR2_X1 U510 ( .A(n515), .B(KEYINPUT100), .Z(n457) );
  XOR2_X1 U511 ( .A(n457), .B(KEYINPUT27), .Z(n469) );
  INV_X1 U512 ( .A(n469), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n562), .A2(n458), .ZN(n459) );
  XNOR2_X1 U514 ( .A(KEYINPUT103), .B(n459), .ZN(n464) );
  OR2_X1 U515 ( .A1(n515), .A2(n525), .ZN(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT104), .B(n460), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n461), .A2(n467), .ZN(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT25), .B(n462), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U520 ( .A(KEYINPUT105), .B(n465), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n466), .A2(n512), .ZN(n474) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT69), .ZN(n468) );
  INV_X1 U523 ( .A(n523), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n469), .A2(n512), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT101), .ZN(n522) );
  NOR2_X1 U526 ( .A1(n471), .A2(n522), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n525), .A2(n472), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n474), .A2(n473), .ZN(n487) );
  NAND2_X1 U529 ( .A1(n475), .A2(n487), .ZN(n476) );
  XNOR2_X1 U530 ( .A(KEYINPUT106), .B(n476), .ZN(n501) );
  NAND2_X1 U531 ( .A1(n553), .A2(n566), .ZN(n490) );
  OR2_X1 U532 ( .A1(n501), .A2(n490), .ZN(n484) );
  NOR2_X1 U533 ( .A1(n512), .A2(n484), .ZN(n478) );
  XNOR2_X1 U534 ( .A(KEYINPUT107), .B(KEYINPUT34), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n515), .A2(n484), .ZN(n480) );
  XOR2_X1 U538 ( .A(KEYINPUT108), .B(n480), .Z(n481) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n481), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n525), .A2(n484), .ZN(n483) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U543 ( .A1(n523), .A2(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(KEYINPUT109), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1327GAT) );
  XNOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n493) );
  NAND2_X1 U547 ( .A1(n570), .A2(n487), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n488), .A2(n573), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n489), .B(KEYINPUT37), .ZN(n511) );
  NOR2_X1 U550 ( .A1(n511), .A2(n490), .ZN(n491) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n491), .Z(n498) );
  NOR2_X1 U552 ( .A1(n512), .A2(n498), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U554 ( .A1(n498), .A2(n515), .ZN(n494) );
  XOR2_X1 U555 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  XNOR2_X1 U556 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n525), .A2(n498), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n497), .Z(G1330GAT) );
  NOR2_X1 U560 ( .A1(n498), .A2(n523), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT111), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  NAND2_X1 U563 ( .A1(n563), .A2(n542), .ZN(n510) );
  OR2_X1 U564 ( .A1(n501), .A2(n510), .ZN(n507) );
  NOR2_X1 U565 ( .A1(n512), .A2(n507), .ZN(n502) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(n502), .Z(n503) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n515), .A2(n507), .ZN(n504) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n525), .A2(n507), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT112), .B(n505), .Z(n506) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  NOR2_X1 U573 ( .A1(n523), .A2(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  OR2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n512), .A2(n518), .ZN(n514) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n518), .ZN(n516) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n525), .A2(n518), .ZN(n517) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n523), .A2(n518), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n522), .ZN(n539) );
  NAND2_X1 U588 ( .A1(n539), .A2(n523), .ZN(n524) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n534), .A2(n553), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U593 ( .A1(n534), .A2(n542), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(n529), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n531) );
  NAND2_X1 U597 ( .A1(n534), .A2(n557), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT118), .Z(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n562), .A2(n539), .ZN(n550) );
  NOR2_X1 U606 ( .A1(n563), .A2(n550), .ZN(n540) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n540), .Z(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT120), .B(n541), .ZN(G1344GAT) );
  INV_X1 U609 ( .A(n542), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n543), .A2(n550), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(KEYINPUT53), .B(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n570), .A2(n550), .ZN(n549) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n552), .Z(G1347GAT) );
  XOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT125), .Z(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U625 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT60), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT126), .B(n560), .Z(n565) );
  NAND2_X1 U628 ( .A1(n561), .A2(n562), .ZN(n572) );
  OR2_X1 U629 ( .A1(n572), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1352GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n568) );
  OR2_X1 U632 ( .A1(n572), .A2(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(G204GAT), .B(n569), .Z(G1353GAT) );
  OR2_X1 U635 ( .A1(n572), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT62), .B(n574), .Z(n575) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(n575), .ZN(G1355GAT) );
endmodule

