//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(new_n454), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n464), .A2(new_n465), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n464), .B2(new_n465), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n464), .B2(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  OR2_X1    g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(new_n492), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n490), .B1(new_n494), .B2(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G88), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n507), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n505), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n514), .B(new_n521), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(G90), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n503), .A2(new_n529), .B1(new_n505), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n509), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(G171));
  AND2_X1   g109(.A1(new_n501), .A2(G56), .ZN(new_n535));
  AND2_X1   g110(.A1(G68), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(G651), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  INV_X1    g115(.A(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n518), .B2(new_n519), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n520), .A2(G81), .B1(new_n542), .B2(G43), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n505), .A2(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n542), .B(G53), .C1(new_n551), .C2(new_n552), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT72), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT5), .A2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n515), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(KEYINPUT73), .A3(G651), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(new_n567), .B1(G91), .B2(new_n520), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n558), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n542), .B2(G49), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n503), .ZN(G288));
  AND2_X1   g151(.A1(KEYINPUT6), .A2(G651), .ZN(new_n577));
  NOR2_X1   g152(.A1(KEYINPUT6), .A2(G651), .ZN(new_n578));
  OAI211_X1 g153(.A(G48), .B(G543), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n502), .A2(KEYINPUT75), .A3(G48), .A4(G543), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n581), .A2(new_n582), .B1(new_n520), .B2(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(G61), .B1(new_n560), .B2(new_n515), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT74), .B1(new_n586), .B2(G651), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n588));
  AOI211_X1 g163(.A(new_n588), .B(new_n509), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n583), .B1(new_n587), .B2(new_n589), .ZN(G305));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n503), .A2(new_n591), .B1(new_n505), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n509), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n501), .A2(new_n502), .A3(G92), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n561), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n542), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n558), .A2(new_n568), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NOR2_X1   g189(.A1(new_n605), .A2(G559), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n497), .A2(new_n471), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n476), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n478), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n463), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(KEYINPUT79), .ZN(new_n640));
  INV_X1    g215(.A(G1341), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(KEYINPUT79), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(G1348), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT78), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2451), .Z(new_n649));
  XOR2_X1   g224(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n639), .B(KEYINPUT79), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G1341), .ZN(new_n654));
  INV_X1    g229(.A(G1348), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n643), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n646), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n652), .B1(new_n646), .B2(new_n656), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  INV_X1    g243(.A(new_n661), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n668), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n678), .A2(KEYINPUT82), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(KEYINPUT82), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(new_n685), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n681), .B1(new_n679), .B2(new_n680), .ZN(new_n691));
  MUX2_X1   g266(.A(new_n685), .B(new_n690), .S(new_n691), .Z(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n689), .B1(new_n688), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n677), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(new_n692), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT83), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n700), .A2(new_n693), .A3(new_n676), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n696), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n698), .B1(new_n696), .B2(new_n701), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n675), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n704), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(new_n674), .A3(new_n702), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G32), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n471), .A2(G105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT90), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n476), .A2(G141), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n478), .A2(G129), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n711), .B1(new_n722), .B2(new_n710), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G1996), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n710), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n710), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT29), .B(G2090), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(new_n710), .ZN(new_n733));
  INV_X1    g308(.A(G160), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n710), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2084), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G5), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G171), .B2(new_n737), .ZN(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  NOR2_X1   g315(.A1(G164), .A2(new_n710), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G27), .B2(new_n710), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n736), .B1(G1961), .B2(new_n739), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n726), .A2(new_n730), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n737), .A2(G20), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT94), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n610), .B2(new_n737), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT95), .B(G1956), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G16), .A2(G19), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n544), .B2(G16), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT86), .B(G1341), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n737), .A2(G4), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n606), .B2(new_n737), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1348), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n710), .A2(G26), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT28), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n476), .A2(G140), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT88), .Z(new_n765));
  INV_X1    g340(.A(G116), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n470), .B1(new_n766), .B2(G2105), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(new_n767), .B1(new_n478), .B2(G128), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n760), .B1(new_n769), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2067), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n742), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G2078), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n710), .A2(G33), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(new_n463), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n476), .A2(G139), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n775), .B1(new_n784), .B2(new_n710), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2072), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n758), .A2(new_n772), .A3(new_n774), .A4(new_n786), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n744), .A2(new_n755), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT30), .B(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n710), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n631), .B2(new_n710), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n739), .B2(G1961), .ZN(new_n794));
  NOR2_X1   g369(.A1(G168), .A2(new_n737), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n737), .B2(G21), .ZN(new_n796));
  INV_X1    g371(.A(G1966), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n788), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n710), .A2(G25), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n476), .A2(G131), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT84), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(G107), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G2105), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n478), .B2(G119), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n802), .B1(new_n809), .B2(new_n710), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  XOR2_X1   g386(.A(new_n810), .B(new_n811), .Z(new_n812));
  INV_X1    g387(.A(KEYINPUT85), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n737), .A2(G24), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n596), .B2(new_n737), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1986), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n737), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n737), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(G6), .A2(G16), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G305), .B2(new_n737), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT32), .B(G1981), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n737), .A2(G23), .ZN(new_n830));
  INV_X1    g405(.A(G288), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n737), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT33), .B(G1976), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n823), .A2(new_n828), .A3(new_n829), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(KEYINPUT34), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n819), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n801), .B1(new_n839), .B2(new_n840), .ZN(G311));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n839), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n842), .A2(new_n800), .A3(new_n788), .ZN(G150));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n503), .A2(new_n844), .B1(new_n505), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(new_n509), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT96), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n544), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n846), .A2(new_n848), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(KEYINPUT96), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n852), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n606), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT97), .ZN(new_n864));
  AOI21_X1  g439(.A(G860), .B1(new_n861), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n853), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n869), .ZN(G145));
  NAND2_X1  g445(.A1(new_n494), .A2(new_n499), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n487), .B1(new_n495), .B2(new_n496), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n463), .A2(G114), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT99), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n486), .A2(new_n489), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n769), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n769), .A2(new_n879), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n783), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n783), .B1(new_n880), .B2(new_n881), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n883), .A2(new_n721), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n769), .B(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n784), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n722), .B1(new_n887), .B2(new_n882), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n804), .A2(new_n808), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n622), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n476), .A2(G142), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT100), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G118), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n893), .A2(new_n894), .B1(new_n896), .B2(G2105), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n478), .A2(G130), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n890), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n885), .A2(new_n888), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n631), .B(new_n734), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n482), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n721), .B1(new_n883), .B2(new_n884), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n890), .B(new_n899), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n887), .A2(new_n722), .A3(new_n882), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT102), .A4(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n885), .B2(new_n888), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n901), .A3(new_n909), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g492(.A1(new_n853), .A2(G868), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n858), .A2(new_n616), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n615), .B1(new_n851), .B2(new_n857), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(G299), .A2(new_n605), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n606), .A2(new_n558), .A3(new_n568), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n923), .A2(KEYINPUT103), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT103), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n927), .A3(KEYINPUT104), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  INV_X1    g504(.A(new_n924), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n606), .B1(new_n568), .B2(new_n558), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n924), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n921), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT104), .B1(new_n922), .B2(new_n927), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT106), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n934), .A4(new_n928), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n596), .B(G288), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G303), .B(G305), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n942), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n944), .A2(new_n942), .A3(new_n941), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT42), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n937), .A2(new_n940), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n935), .A2(new_n936), .ZN(new_n951));
  INV_X1    g526(.A(new_n949), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n939), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n918), .B1(new_n954), .B2(G868), .ZN(G295));
  AOI21_X1  g530(.A(new_n918), .B1(new_n954), .B2(G868), .ZN(G331));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g532(.A1(G286), .A2(G301), .ZN(new_n958));
  NAND2_X1  g533(.A1(G168), .A2(G171), .ZN(new_n959));
  AND4_X1   g534(.A1(new_n851), .A2(new_n958), .A3(new_n857), .A4(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n851), .A2(new_n857), .B1(new_n958), .B2(new_n959), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n932), .B(new_n933), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n959), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n858), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n851), .A2(new_n958), .A3(new_n857), .A4(new_n959), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(new_n923), .A3(new_n924), .A4(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n948), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n915), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n948), .B1(new_n962), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n957), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n965), .B(new_n964), .C1(new_n925), .C2(new_n926), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n962), .ZN(new_n972));
  INV_X1    g547(.A(new_n948), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n974), .A2(KEYINPUT43), .A3(new_n915), .A4(new_n967), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT44), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n968), .B2(new_n969), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n974), .A2(new_n957), .A3(new_n915), .A4(new_n967), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n970), .B2(new_n975), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT44), .B1(new_n978), .B2(new_n979), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT107), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(G397));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n879), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT108), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT45), .B1(new_n990), .B2(KEYINPUT108), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n468), .A2(new_n473), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n721), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n769), .A2(G2067), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n763), .A2(new_n771), .A3(new_n768), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n997), .A2(KEYINPUT111), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT111), .B1(new_n997), .B2(new_n1003), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1000), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n997), .A2(G1996), .A3(new_n721), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n809), .A2(new_n811), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n809), .A2(new_n811), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n997), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1986), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n596), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT109), .Z(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n1015), .B2(new_n596), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n997), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n583), .B(new_n1021), .C1(new_n587), .C2(new_n589), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n585), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n501), .B2(G61), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n588), .B1(new_n1025), .B2(new_n509), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n586), .A2(KEYINPUT74), .A3(G651), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1021), .B1(new_n1028), .B2(new_n583), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1020), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G305), .A2(G1981), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1022), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n872), .A2(new_n875), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1034), .A2(new_n877), .B1(new_n494), .B2(new_n499), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n1035), .B2(new_n876), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1036), .B2(new_n995), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1030), .A2(new_n1032), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT114), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1030), .A2(new_n1032), .A3(new_n1040), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1384), .B1(new_n871), .B2(new_n1034), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(KEYINPUT45), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n879), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT112), .B(new_n1047), .C1(G164), .C2(G1384), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1045), .A2(new_n995), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n822), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n871), .A2(new_n1034), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n989), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n996), .B1(new_n1052), .B2(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g628(.A(G2090), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n879), .A2(new_n1055), .A3(new_n989), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1050), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n879), .A2(new_n995), .A3(new_n989), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n574), .B(G1976), .C1(new_n575), .C2(new_n503), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(G8), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1066), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1063), .A2(new_n1064), .A3(G8), .A4(new_n1068), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n831), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1042), .A2(new_n1062), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n995), .C1(new_n1036), .C2(new_n1055), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1055), .B1(new_n879), .B2(new_n989), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT115), .B1(new_n1075), .B2(new_n996), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1052), .A2(KEYINPUT50), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1074), .A2(new_n1076), .A3(new_n1054), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1050), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1061), .B1(new_n1080), .B2(G8), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1072), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n996), .B1(KEYINPUT45), .B2(new_n1044), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n990), .A2(new_n1047), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT53), .A4(new_n740), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1056), .A2(new_n1086), .A3(new_n995), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT122), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1085), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1049), .B2(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1082), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1036), .A2(KEYINPUT45), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n995), .B1(new_n1052), .B2(new_n1047), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n797), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G2084), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1053), .A2(new_n1102), .A3(new_n1056), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1103), .A3(G168), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1104), .A2(new_n1105), .A3(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G286), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n1104), .A3(G8), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1106), .B1(new_n1109), .B2(KEYINPUT51), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1104), .A2(G8), .ZN(new_n1113));
  AOI21_X1  g688(.A(G168), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT51), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(KEYINPUT51), .B2(new_n1113), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1098), .A2(new_n1112), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1074), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1122));
  INV_X1    g697(.A(G1956), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1049), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n555), .B2(new_n556), .ZN(new_n1127));
  AOI22_X1  g702(.A1(G299), .A2(KEYINPUT57), .B1(new_n568), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1121), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1087), .A2(new_n655), .ZN(new_n1130));
  AND4_X1   g705(.A1(new_n989), .A2(new_n879), .A3(new_n995), .A4(new_n771), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n606), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n568), .A2(new_n1127), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n610), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n996), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1077), .B1(new_n1138), .B2(new_n1073), .ZN(new_n1139));
  AOI21_X1  g714(.A(G1956), .B1(new_n1139), .B2(new_n1076), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1125), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1049), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT117), .B(new_n1137), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1129), .A2(new_n1134), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1142), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(new_n1128), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  NOR4_X1   g724(.A1(new_n468), .A2(new_n473), .A3(new_n994), .A4(G1996), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .A4(new_n1150), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1063), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT118), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1151), .A2(new_n1156), .A3(new_n1153), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n544), .A2(KEYINPUT119), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1149), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1151), .A2(new_n1156), .A3(new_n1153), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1156), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1149), .B(new_n1159), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1137), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT61), .B1(new_n1166), .B2(new_n1147), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1131), .B1(new_n1087), .B2(new_n655), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n606), .B1(new_n1168), .B2(KEYINPUT60), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1168), .A2(new_n1170), .A3(KEYINPUT60), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1170), .B1(new_n1168), .B2(KEYINPUT60), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n605), .B1(new_n1133), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n1132), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1168), .A2(new_n1170), .A3(KEYINPUT60), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1165), .A2(new_n1167), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1126), .A2(KEYINPUT120), .A3(new_n1128), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1182), .A2(KEYINPUT61), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1147), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1183), .A2(new_n1129), .A3(new_n1143), .A4(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1148), .B1(new_n1181), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1094), .A2(G301), .A3(new_n1096), .ZN(new_n1188));
  INV_X1    g763(.A(new_n993), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n740), .A4(new_n995), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1096), .B(new_n1089), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1191), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1192));
  AOI21_X1  g767(.A(KEYINPUT123), .B1(new_n1191), .B2(G171), .ZN(new_n1193));
  OAI211_X1 g768(.A(KEYINPUT54), .B(new_n1188), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT54), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1191), .A2(G171), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1195), .B1(new_n1097), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1194), .A2(new_n1197), .A3(new_n1116), .A4(new_n1082), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1120), .B1(new_n1187), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1080), .A2(G8), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1061), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1071), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1203), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1204));
  NOR2_X1   g779(.A1(G286), .A2(new_n1033), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1107), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1202), .A2(new_n1062), .A3(new_n1204), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT63), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1072), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1061), .B1(new_n1058), .B2(G8), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1107), .A2(KEYINPUT63), .A3(new_n1205), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1209), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1062), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1204), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g792(.A1(G288), .A2(G1976), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1023), .B1(new_n1042), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1037), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(KEYINPUT116), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1215), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI22_X1  g799(.A1(new_n1207), .A2(new_n1208), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1225));
  OAI21_X1  g800(.A(KEYINPUT116), .B1(new_n1225), .B2(new_n1221), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1019), .B1(new_n1199), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT125), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1006), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1230), .A2(new_n1002), .ZN(new_n1231));
  AOI21_X1  g806(.A(new_n1229), .B1(new_n1231), .B2(new_n997), .ZN(new_n1232));
  INV_X1    g807(.A(new_n997), .ZN(new_n1233));
  AOI211_X1 g808(.A(KEYINPUT125), .B(new_n1233), .C1(new_n1230), .C2(new_n1002), .ZN(new_n1234));
  OAI21_X1  g809(.A(new_n997), .B1(new_n721), .B2(new_n1003), .ZN(new_n1235));
  XNOR2_X1  g810(.A(new_n1235), .B(KEYINPUT126), .ZN(new_n1236));
  INV_X1    g811(.A(KEYINPUT47), .ZN(new_n1237));
  XNOR2_X1  g812(.A(new_n999), .B(KEYINPUT46), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g814(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g815(.A(new_n1237), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g816(.A1(new_n1233), .A2(new_n1017), .ZN(new_n1242));
  XNOR2_X1  g817(.A(new_n1242), .B(KEYINPUT48), .ZN(new_n1243));
  OAI22_X1  g818(.A1(new_n1240), .A2(new_n1241), .B1(new_n1014), .B2(new_n1243), .ZN(new_n1244));
  NOR3_X1   g819(.A1(new_n1232), .A2(new_n1234), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1228), .A2(new_n1245), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g821(.A(new_n916), .B1(new_n978), .B2(new_n979), .ZN(new_n1248));
  NOR2_X1   g822(.A1(G227), .A2(new_n461), .ZN(new_n1249));
  INV_X1    g823(.A(new_n1249), .ZN(new_n1250));
  NOR2_X1   g824(.A1(G401), .A2(new_n1250), .ZN(new_n1251));
  AND3_X1   g825(.A1(new_n708), .A2(new_n1251), .A3(KEYINPUT127), .ZN(new_n1252));
  AOI21_X1  g826(.A(KEYINPUT127), .B1(new_n708), .B2(new_n1251), .ZN(new_n1253));
  OAI21_X1  g827(.A(new_n1248), .B1(new_n1252), .B2(new_n1253), .ZN(G225));
  INV_X1    g828(.A(G225), .ZN(G308));
endmodule


