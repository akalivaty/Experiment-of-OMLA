//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1224, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n207), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n203), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n209), .A3(new_n230), .ZN(new_n231));
  NOR4_X1   g0031(.A1(new_n218), .A2(new_n219), .A3(new_n228), .A4(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NOR2_X1   g0048(.A1(new_n202), .A2(new_n203), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G58), .A2(G68), .ZN(new_n250));
  OAI21_X1  g0050(.A(G20), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G159), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n209), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT7), .B1(new_n258), .B2(new_n209), .ZN(new_n260));
  OAI21_X1  g0060(.A(G68), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT79), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n263), .B(KEYINPUT16), .C1(new_n262), .C2(new_n261), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT16), .ZN(new_n265));
  INV_X1    g0065(.A(new_n261), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n255), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n230), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(G274), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n271), .A2(new_n275), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n278), .B2(new_n221), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT81), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT81), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n276), .B(new_n281), .C1(new_n278), .C2(new_n221), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT66), .B(G1698), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G87), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n285), .A2(new_n258), .B1(new_n253), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n271), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n279), .B1(new_n271), .B2(new_n287), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n283), .A2(new_n290), .B1(new_n291), .B2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G1), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT8), .B(G58), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(new_n208), .B2(G20), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n269), .B(new_n296), .C1(new_n298), .C2(KEYINPUT80), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(KEYINPUT80), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n299), .A2(new_n300), .B1(new_n296), .B2(new_n297), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n270), .A2(new_n292), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT17), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT17), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n270), .A2(new_n292), .A3(new_n304), .A4(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT83), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n306), .B(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(G179), .B1(new_n287), .B2(new_n271), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(new_n280), .A3(new_n282), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n291), .B2(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n270), .B2(new_n301), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT82), .B1(new_n312), .B2(KEYINPUT18), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(KEYINPUT18), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(KEYINPUT82), .A3(KEYINPUT18), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n204), .A2(G20), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n209), .A2(G33), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n319), .B1(new_n320), .B2(new_n254), .C1(new_n321), .C2(new_n297), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n322), .A2(new_n269), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n296), .A2(new_n201), .ZN(new_n324));
  INV_X1    g0124(.A(new_n269), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(G1), .B2(new_n209), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n326), .B2(new_n201), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT9), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n275), .ZN(new_n331));
  INV_X1    g0131(.A(G274), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n331), .A2(new_n271), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G226), .B2(new_n277), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT3), .B(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G223), .A2(G1698), .ZN(new_n336));
  INV_X1    g0136(.A(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT66), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G222), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n335), .B(new_n336), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n343), .B(new_n271), .C1(G77), .C2(new_n335), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n289), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(G200), .B2(new_n345), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT68), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n330), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n330), .A2(KEYINPUT68), .ZN(new_n352));
  AOI211_X1 g0152(.A(KEYINPUT69), .B(new_n346), .C1(G200), .C2(new_n345), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n354), .B2(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(new_n345), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n356), .A2(G169), .B1(new_n323), .B2(new_n327), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n357), .A2(KEYINPUT67), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(KEYINPUT67), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n335), .B1(new_n222), .B2(new_n337), .C1(new_n341), .C2(new_n221), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n271), .C1(G107), .C2(new_n335), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n333), .B1(G244), .B2(new_n277), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G190), .ZN(new_n367));
  INV_X1    g0167(.A(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n296), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n326), .B2(new_n368), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G20), .A2(G77), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n297), .B2(new_n254), .C1(new_n321), .C2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n269), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n367), .B(new_n374), .C1(new_n375), .C2(new_n366), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n374), .B1(new_n366), .B2(new_n359), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(G169), .B2(new_n366), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n362), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n355), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n318), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT14), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT13), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT71), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n338), .A2(new_n340), .A3(G226), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n221), .A2(new_n337), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n258), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT70), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n389), .B(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n384), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n389), .B(KEYINPUT70), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n386), .B1(new_n284), .B2(G226), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT71), .B(new_n393), .C1(new_n394), .C2(new_n258), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n271), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(KEYINPUT72), .A3(new_n271), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n276), .B1(new_n278), .B2(new_n222), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT73), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n383), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT72), .B1(new_n396), .B2(new_n271), .ZN(new_n405));
  AOI211_X1 g0205(.A(new_n398), .B(new_n272), .C1(new_n392), .C2(new_n395), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n403), .B(new_n383), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n382), .B(G169), .C1(new_n404), .C2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(G179), .A3(new_n407), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G169), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n411), .B2(new_n407), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT76), .B1(new_n415), .B2(new_n382), .ZN(new_n416));
  OAI21_X1  g0216(.A(G169), .B1(new_n404), .B2(new_n408), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT14), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n413), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n203), .B1(new_n326), .B2(KEYINPUT12), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT11), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n203), .A2(G20), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n423), .B1(new_n321), .B2(new_n368), .C1(new_n201), .C2(new_n254), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n269), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n421), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT12), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n423), .A2(new_n427), .A3(G1), .A4(new_n293), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n427), .B2(new_n295), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n426), .B(new_n429), .C1(new_n422), .C2(new_n425), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT74), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n420), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT75), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n411), .A2(G190), .A3(new_n407), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n432), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n375), .B1(new_n411), .B2(new_n407), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(G200), .B1(new_n404), .B2(new_n408), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(KEYINPUT75), .A3(new_n432), .A4(new_n438), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n381), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT78), .B1(new_n436), .B2(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n208), .B(G45), .C1(new_n273), .C2(KEYINPUT5), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(KEYINPUT5), .B2(new_n273), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n271), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G257), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(G274), .A3(new_n272), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n335), .A2(new_n284), .A3(G244), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT4), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n335), .A2(G250), .A3(G1698), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n456), .A2(new_n457), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n271), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n359), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n254), .A2(new_n368), .ZN(new_n466));
  INV_X1    g0266(.A(G107), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  XOR2_X1   g0271(.A(G97), .B(G107), .Z(new_n472));
  OAI211_X1 g0272(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(KEYINPUT6), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n466), .B1(new_n473), .B2(G20), .ZN(new_n474));
  OAI21_X1  g0274(.A(G107), .B1(new_n259), .B2(new_n260), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n325), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n296), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n325), .B(new_n295), .C1(G1), .C2(new_n253), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n477), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n455), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n414), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n465), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(G200), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n481), .C1(new_n289), .C2(new_n483), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n335), .A2(new_n209), .A3(G87), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n488), .B(KEYINPUT22), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT24), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT90), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G116), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(G20), .ZN(new_n493));
  OR3_X1    g0293(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n209), .A2(KEYINPUT90), .A3(G33), .A4(G116), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n496));
  AND4_X1   g0296(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n490), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n490), .B1(new_n489), .B2(new_n497), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n269), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n452), .A2(G264), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n454), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n214), .A2(new_n337), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n335), .A2(new_n504), .B1(G33), .B2(G294), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n335), .A2(new_n284), .A3(G250), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n272), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(G200), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n296), .A2(new_n467), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(KEYINPUT25), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n510), .B(new_n511), .C1(new_n467), .C2(new_n479), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n503), .A2(new_n507), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G190), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n501), .A2(new_n508), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n485), .A2(new_n487), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n501), .A2(new_n513), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT91), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n501), .A2(KEYINPUT91), .A3(new_n513), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n507), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n502), .A2(new_n524), .A3(G179), .A4(new_n454), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n514), .B2(new_n414), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n517), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT86), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n335), .A2(G244), .A3(G1698), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n529), .A2(KEYINPUT85), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(KEYINPUT85), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n335), .A2(G238), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n492), .B1(new_n533), .B2(new_n341), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n271), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n208), .A2(new_n332), .A3(G45), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n207), .B1(new_n274), .B2(G1), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n272), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n414), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n534), .B1(new_n530), .B2(new_n531), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n272), .ZN(new_n541));
  INV_X1    g0341(.A(new_n538), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n541), .A2(new_n359), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n528), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n535), .A2(G179), .A3(new_n538), .ZN(new_n545));
  OAI21_X1  g0345(.A(G169), .B1(new_n541), .B2(new_n542), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT86), .ZN(new_n547));
  NOR3_X1   g0347(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n391), .A2(KEYINPUT19), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n209), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n335), .A2(new_n209), .A3(G68), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n321), .A2(new_n477), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(KEYINPUT19), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n269), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n296), .A2(new_n372), .ZN(new_n555));
  INV_X1    g0355(.A(new_n479), .ZN(new_n556));
  INV_X1    g0356(.A(new_n372), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n544), .A2(new_n547), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(G200), .B1(new_n541), .B2(new_n542), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(G87), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n554), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G190), .B(new_n538), .C1(new_n540), .C2(new_n272), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT87), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT87), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n560), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n295), .A2(G116), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n556), .B2(G116), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n459), .B(new_n209), .C1(G33), .C2(new_n477), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n572), .B(new_n269), .C1(new_n209), .C2(G116), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n452), .A2(G270), .ZN(new_n577));
  INV_X1    g0377(.A(G303), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n272), .B1(new_n578), .B2(new_n258), .ZN(new_n579));
  OAI221_X1 g0379(.A(new_n335), .B1(new_n215), .B2(new_n337), .C1(new_n341), .C2(new_n214), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT88), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT88), .B1(new_n579), .B2(new_n580), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n454), .B(new_n577), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n576), .B1(new_n584), .B2(G200), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n289), .B2(new_n584), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n414), .B1(new_n571), .B2(new_n575), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n587), .A3(KEYINPUT21), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n359), .B1(new_n571), .B2(new_n575), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n579), .A2(new_n580), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT88), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n581), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n589), .A2(new_n593), .A3(new_n454), .A4(new_n577), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT21), .B1(new_n584), .B2(new_n587), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(KEYINPUT89), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT89), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n598), .B(KEYINPUT21), .C1(new_n584), .C2(new_n587), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n586), .B(new_n595), .C1(new_n597), .C2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n527), .A2(new_n567), .A3(new_n569), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n449), .A2(new_n602), .ZN(G372));
  INV_X1    g0403(.A(new_n362), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n306), .B(KEYINPUT83), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n444), .A2(new_n378), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(new_n436), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n270), .A2(new_n301), .ZN(new_n608));
  INV_X1    g0408(.A(new_n311), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT93), .A3(new_n314), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT93), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n312), .A2(KEYINPUT18), .ZN(new_n615));
  AOI211_X1 g0415(.A(new_n611), .B(new_n311), .C1(new_n270), .C2(new_n301), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n607), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n355), .B(KEYINPUT94), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n604), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n559), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n545), .B2(new_n546), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  INV_X1    g0424(.A(new_n485), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n518), .A2(new_n526), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n626), .B(new_n595), .C1(new_n597), .C2(new_n599), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n487), .A2(new_n516), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT92), .B1(new_n630), .B2(new_n623), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n559), .B1(new_n539), .B2(new_n543), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT92), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n565), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n624), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n485), .A2(new_n624), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n567), .A2(new_n569), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n623), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n621), .B1(new_n449), .B2(new_n639), .ZN(G369));
  NAND2_X1  g0440(.A1(new_n523), .A2(new_n526), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n294), .A2(new_n209), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(G213), .ZN(new_n645));
  XOR2_X1   g0445(.A(KEYINPUT95), .B(G343), .Z(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n641), .B(new_n516), .C1(new_n522), .C2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n595), .B1(new_n597), .B2(new_n599), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n648), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n518), .A2(new_n526), .A3(new_n648), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n576), .A2(new_n647), .ZN(new_n656));
  MUX2_X1   g0456(.A(new_n650), .B(new_n601), .S(new_n656), .Z(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n649), .B1(new_n641), .B2(new_n648), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n655), .A2(new_n661), .ZN(G399));
  NOR2_X1   g0462(.A1(new_n213), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(G116), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n548), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n663), .A2(new_n665), .A3(new_n208), .ZN(new_n666));
  INV_X1    g0466(.A(new_n663), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n666), .A2(KEYINPUT96), .B1(new_n229), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(KEYINPUT96), .B2(new_n666), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT28), .Z(new_n670));
  INV_X1    g0470(.A(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n636), .A2(new_n638), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n647), .B1(new_n672), .B2(new_n632), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n671), .B1(new_n673), .B2(KEYINPUT29), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  OAI211_X1 g0475(.A(KEYINPUT99), .B(new_n675), .C1(new_n639), .C2(new_n647), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n635), .A2(new_n517), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n650), .B1(new_n523), .B2(new_n526), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n632), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n567), .A2(new_n569), .A3(new_n625), .ZN(new_n680));
  INV_X1    g0480(.A(new_n635), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n680), .A2(new_n624), .B1(new_n681), .B2(new_n637), .ZN(new_n682));
  OAI211_X1 g0482(.A(KEYINPUT29), .B(new_n648), .C1(new_n679), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n674), .A2(new_n676), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT31), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n593), .A2(new_n577), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n541), .A2(new_n542), .ZN(new_n687));
  INV_X1    g0487(.A(new_n525), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(KEYINPUT97), .A3(KEYINPUT30), .A4(new_n464), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT97), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n686), .A2(new_n687), .A3(new_n464), .A4(new_n688), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n687), .A2(G179), .A3(new_n514), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n584), .A2(new_n483), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g0500(.A(new_n685), .B(new_n648), .C1(new_n695), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT98), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n695), .A2(new_n700), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT98), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n696), .A2(new_n699), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n694), .B2(new_n690), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n685), .B1(new_n708), .B2(new_n648), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n702), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n602), .A2(new_n647), .ZN(new_n711));
  OAI21_X1  g0511(.A(G330), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n684), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n670), .B1(new_n713), .B2(G1), .ZN(G364));
  NOR2_X1   g0514(.A1(new_n293), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n208), .B1(new_n715), .B2(G45), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n663), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n212), .A2(new_n335), .ZN(new_n719));
  INV_X1    g0519(.A(G355), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n719), .A2(new_n720), .B1(G116), .B2(new_n212), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n213), .A2(new_n335), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n229), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n274), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n244), .A2(G45), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT100), .Z(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n230), .B1(G20), .B2(new_n414), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n718), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n731), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n209), .A2(new_n289), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n375), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G87), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n335), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n209), .B1(new_n742), .B2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n741), .B1(G97), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n209), .A2(G190), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n742), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n252), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT32), .ZN(new_n749));
  NAND3_X1  g0549(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n289), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(G190), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G50), .A2(new_n751), .B1(new_n752), .B2(G68), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n359), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n746), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n746), .A2(new_n737), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n368), .A2(new_n755), .B1(new_n756), .B2(new_n467), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n736), .A2(new_n754), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(G58), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n745), .A2(new_n749), .A3(new_n753), .A4(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n258), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G326), .B2(new_n751), .ZN(new_n764));
  INV_X1    g0564(.A(new_n756), .ZN(new_n765));
  INV_X1    g0565(.A(new_n755), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G283), .A2(new_n765), .B1(new_n766), .B2(G311), .ZN(new_n767));
  INV_X1    g0567(.A(new_n747), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G303), .A2(new_n739), .B1(new_n768), .B2(G329), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n744), .A2(G294), .B1(new_n752), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n764), .A2(new_n767), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n735), .B1(new_n761), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n734), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n730), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n657), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n718), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n658), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n657), .A2(G330), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT101), .Z(G396));
  OAI21_X1  g0581(.A(new_n376), .B1(new_n374), .B2(new_n648), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n378), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n378), .A2(new_n647), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n673), .B(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n718), .B1(new_n788), .B2(new_n712), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n712), .B2(new_n788), .ZN(new_n790));
  INV_X1    g0590(.A(new_n751), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n258), .B1(new_n756), .B2(new_n286), .C1(new_n791), .C2(new_n578), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(G283), .B2(new_n752), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n758), .A2(new_n794), .B1(new_n743), .B2(new_n477), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT102), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n768), .A2(G311), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G107), .A2(new_n739), .B1(new_n766), .B2(G116), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n793), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G143), .A2(new_n759), .B1(new_n766), .B2(G159), .ZN(new_n800));
  INV_X1    g0600(.A(G137), .ZN(new_n801));
  INV_X1    g0601(.A(new_n752), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(new_n791), .B2(new_n801), .C1(new_n320), .C2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT103), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n335), .B1(new_n756), .B2(new_n203), .ZN(new_n806));
  INV_X1    g0606(.A(G132), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n738), .A2(new_n201), .B1(new_n747), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(G58), .C2(new_n744), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n799), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n731), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n731), .A2(new_n728), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n777), .B1(new_n368), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(new_n787), .C2(new_n729), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n790), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G384));
  NOR2_X1   g0618(.A1(new_n715), .A2(new_n208), .ZN(new_n819));
  INV_X1    g0619(.A(G330), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n602), .A2(new_n647), .B1(new_n704), .B2(KEYINPUT112), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT112), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n701), .B1(new_n709), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n787), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n441), .A2(new_n443), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n434), .A2(new_n647), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(new_n420), .C2(new_n435), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n420), .B2(new_n825), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT107), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(KEYINPUT107), .B(new_n826), .C1(new_n420), .C2(new_n825), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT108), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n826), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n409), .A2(new_n412), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n418), .B1(new_n417), .B2(KEYINPUT14), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n382), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n444), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT107), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT108), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n828), .A2(new_n829), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n827), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n824), .B1(new_n832), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n263), .B1(new_n262), .B2(new_n261), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n265), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(new_n269), .A3(new_n264), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n301), .ZN(new_n848));
  INV_X1    g0648(.A(new_n645), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n315), .A2(new_n316), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n605), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n848), .A2(new_n609), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n850), .A3(new_n302), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT37), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n645), .B1(new_n270), .B2(new_n301), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(new_n302), .A3(new_n610), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n844), .B1(new_n852), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT38), .B(new_n859), .C1(new_n318), .C2(new_n850), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT40), .B1(new_n843), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n610), .A2(new_n302), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT110), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT110), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n856), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n866), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT111), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n868), .A2(new_n873), .A3(new_n857), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n858), .A2(KEYINPUT111), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n613), .A2(new_n617), .B1(new_n303), .B2(new_n305), .ZN(new_n877));
  INV_X1    g0677(.A(new_n856), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n872), .A2(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n844), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n865), .B1(new_n880), .B2(new_n862), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n864), .B1(new_n843), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n823), .ZN(new_n883));
  INV_X1    g0683(.A(new_n821), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n449), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n820), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n882), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n618), .A2(new_n849), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n880), .A2(new_n862), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n889), .B1(KEYINPUT39), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n436), .A2(KEYINPUT109), .A3(new_n648), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n837), .A2(new_n434), .A3(new_n648), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n888), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n784), .B1(new_n673), .B2(new_n787), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n842), .B2(new_n832), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n863), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n621), .B1(new_n684), .B2(new_n449), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n819), .B1(new_n887), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n903), .B2(new_n887), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n230), .A2(new_n209), .A3(new_n664), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n473), .B(KEYINPUT104), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT35), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n909), .B2(new_n908), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT105), .ZN(new_n912));
  XNOR2_X1  g0712(.A(KEYINPUT106), .B(KEYINPUT36), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n249), .A2(new_n229), .A3(new_n368), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n203), .A2(G50), .ZN(new_n916));
  OAI211_X1 g0716(.A(G1), .B(new_n293), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n905), .A2(new_n914), .A3(new_n917), .ZN(G367));
  NOR2_X1   g0718(.A1(new_n738), .A2(new_n664), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(KEYINPUT46), .B1(G311), .B2(new_n751), .ZN(new_n920));
  OAI221_X1 g0720(.A(new_n920), .B1(KEYINPUT46), .B2(new_n919), .C1(new_n467), .C2(new_n743), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n768), .A2(G317), .ZN(new_n922));
  INV_X1    g0722(.A(G283), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n922), .B1(new_n923), .B2(new_n755), .C1(new_n578), .C2(new_n758), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n258), .B1(new_n756), .B2(new_n477), .C1(new_n802), .C2(new_n794), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n765), .A2(G77), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n801), .B2(new_n747), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n335), .B1(new_n743), .B2(new_n203), .C1(new_n320), .C2(new_n758), .ZN(new_n929));
  INV_X1    g0729(.A(G143), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n802), .A2(new_n252), .B1(new_n791), .B2(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n738), .A2(new_n202), .B1(new_n755), .B2(new_n201), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n928), .A2(new_n929), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT47), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n731), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n733), .B1(new_n213), .B2(new_n557), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n722), .A2(new_n240), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n777), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n681), .B1(new_n563), .B2(new_n648), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n632), .A2(new_n563), .A3(new_n648), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n936), .B(new_n939), .C1(new_n942), .C2(new_n775), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT113), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n625), .A2(new_n647), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n485), .B(new_n487), .C1(new_n481), .C2(new_n648), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n649), .A2(new_n948), .A3(new_n651), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n485), .B1(new_n641), .B2(new_n946), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n949), .A2(KEYINPUT42), .B1(new_n648), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(KEYINPUT42), .B2(new_n949), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n661), .A2(new_n948), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT44), .B1(new_n655), .B2(new_n947), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n654), .A2(new_n960), .A3(new_n948), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n652), .A2(new_n653), .A3(new_n947), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT45), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n659), .B(new_n660), .C1(new_n962), .C2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n963), .B(KEYINPUT45), .Z(new_n966));
  NAND4_X1  g0766(.A1(new_n966), .A2(new_n661), .A3(new_n959), .A4(new_n961), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n651), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n652), .B1(new_n660), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n659), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n713), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n713), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n663), .B(KEYINPUT41), .Z(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n717), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n944), .B1(new_n958), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n958), .A2(new_n976), .A3(new_n944), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n943), .B1(new_n978), .B2(new_n979), .ZN(G387));
  NAND2_X1  g0780(.A1(new_n971), .A2(new_n717), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n660), .A2(new_n775), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n237), .A2(G45), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT114), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n297), .A2(G50), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT50), .ZN(new_n986));
  AOI211_X1 g0786(.A(G45), .B(new_n665), .C1(G68), .C2(G77), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n723), .B(new_n984), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n665), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n719), .A2(new_n989), .B1(G107), .B2(new_n212), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n732), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n738), .A2(new_n368), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n758), .A2(new_n201), .B1(new_n755), .B2(new_n203), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G150), .C2(new_n768), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n335), .B1(new_n756), .B2(new_n477), .ZN(new_n995));
  INV_X1    g0795(.A(new_n297), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(new_n752), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n751), .A2(G159), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n744), .A2(new_n557), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n994), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n335), .B1(new_n768), .B2(G326), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n738), .A2(new_n794), .B1(new_n743), .B2(new_n923), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G317), .A2(new_n759), .B1(new_n766), .B2(G303), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n752), .A2(G311), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n762), .C2(new_n791), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT48), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1001), .B1(new_n664), .B2(new_n756), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1000), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n731), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n991), .A2(new_n718), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n972), .A2(new_n663), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n713), .A2(new_n971), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n981), .B1(new_n982), .B2(new_n1014), .C1(new_n1015), .C2(new_n1016), .ZN(G393));
  AND2_X1   g0817(.A1(new_n968), .A2(new_n972), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n663), .B1(new_n968), .B2(new_n972), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n965), .A2(new_n967), .A3(new_n717), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n759), .A2(G311), .B1(G317), .B2(new_n751), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT52), .Z(new_n1023));
  OAI22_X1  g0823(.A1(new_n738), .A2(new_n923), .B1(new_n747), .B2(new_n762), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G294), .B2(new_n766), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n743), .A2(new_n664), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n258), .B1(new_n756), .B2(new_n467), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G303), .C2(new_n752), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n791), .A2(new_n320), .B1(new_n758), .B2(new_n252), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n743), .A2(new_n368), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n335), .B1(new_n756), .B2(new_n286), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(G50), .C2(new_n752), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n738), .A2(new_n203), .B1(new_n747), .B2(new_n930), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n996), .B2(new_n766), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1031), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n735), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n723), .A2(new_n247), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n733), .B1(G97), .B2(new_n213), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n777), .B(new_n1038), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n947), .B2(new_n775), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1021), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1020), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  NAND2_X1  g0845(.A1(new_n884), .A2(new_n883), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n447), .A2(new_n1046), .A3(G330), .A4(new_n448), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n621), .B(new_n1047), .C1(new_n684), .C2(new_n449), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n832), .A2(new_n842), .ZN(new_n1049));
  OAI211_X1 g0849(.A(G330), .B(new_n787), .C1(new_n821), .C2(new_n823), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT116), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1049), .A2(KEYINPUT116), .A3(new_n1051), .ZN(new_n1055));
  OAI211_X1 g0855(.A(G330), .B(new_n787), .C1(new_n710), .C2(new_n711), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n832), .A2(new_n1056), .A3(new_n842), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n898), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n832), .A2(new_n842), .A3(new_n1050), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1056), .B1(new_n832), .B2(new_n842), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n648), .B(new_n783), .C1(new_n679), .C2(new_n682), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n785), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1048), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT39), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n880), .A2(new_n862), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n861), .B2(new_n862), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n899), .B2(new_n896), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1062), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1049), .A2(new_n1064), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT115), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n896), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n892), .A2(new_n895), .A3(KEYINPUT115), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1076), .A2(new_n890), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1072), .A2(new_n1073), .A3(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1072), .A2(new_n1079), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT117), .B1(new_n1067), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1072), .A2(new_n1079), .A3(new_n1073), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1049), .A2(new_n1059), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n896), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(new_n1071), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1053), .B(new_n1050), .C1(new_n842), .C2(new_n832), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT116), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1084), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT117), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1065), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1093), .C1(new_n1094), .C2(new_n1048), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1083), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n667), .B1(new_n1067), .B2(new_n1082), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1082), .A2(new_n717), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n777), .B1(new_n297), .B2(new_n814), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n335), .B(new_n1032), .C1(G87), .C2(new_n739), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n467), .B2(new_n802), .C1(new_n923), .C2(new_n791), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n203), .A2(new_n756), .B1(new_n755), .B2(new_n477), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n758), .A2(new_n664), .B1(new_n747), .B2(new_n794), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT119), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n759), .A2(G132), .B1(new_n766), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(G125), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n747), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n335), .B1(new_n743), .B2(new_n252), .C1(new_n201), .C2(new_n756), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G128), .A2(new_n751), .B1(new_n752), .B2(G137), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n738), .A2(new_n320), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1116));
  XOR2_X1   g0916(.A(new_n1115), .B(new_n1116), .Z(new_n1117));
  NAND3_X1  g0917(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1106), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(KEYINPUT119), .B2(new_n1105), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1100), .B1(new_n735), .B2(new_n1120), .C1(new_n891), .C2(new_n729), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1099), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1098), .A2(new_n1123), .ZN(G378));
  NAND2_X1  g0924(.A1(new_n1060), .A2(new_n1066), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1048), .B1(new_n1082), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n620), .A2(new_n362), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1128), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n620), .A2(new_n362), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n328), .A2(new_n645), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1133), .A3(new_n1131), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n824), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1049), .A2(new_n1138), .A3(new_n881), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(G330), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1137), .B1(new_n1140), .B2(new_n864), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1049), .A2(new_n863), .A3(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n865), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1137), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n820), .B1(new_n843), .B2(new_n881), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1141), .A2(new_n901), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n901), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT57), .B1(new_n1126), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n901), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1140), .A2(new_n864), .A3(new_n1137), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1144), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1141), .A2(new_n901), .A3(new_n1146), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(KEYINPUT122), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1048), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT122), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1141), .A2(new_n901), .A3(new_n1146), .A4(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n667), .B1(new_n1150), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1156), .A2(new_n717), .A3(new_n1161), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n814), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n718), .B1(G50), .B2(new_n1165), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n791), .A2(new_n664), .B1(new_n743), .B2(new_n203), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT121), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n258), .A2(new_n273), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1169), .B(new_n992), .C1(G97), .C2(new_n752), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G58), .A2(new_n765), .B1(new_n768), .B2(G283), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n759), .A2(G107), .B1(new_n766), .B2(new_n557), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(G33), .A2(G41), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT120), .Z(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(G50), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1173), .A2(new_n1174), .B1(new_n1169), .B2(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n791), .A2(new_n1110), .B1(new_n743), .B2(new_n320), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G128), .A2(new_n759), .B1(new_n739), .B2(new_n1108), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n801), .B2(new_n755), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(G132), .C2(new_n752), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G159), .A2(new_n765), .B1(new_n768), .B2(G124), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT59), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1177), .B(new_n1186), .C1(new_n1183), .C2(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1179), .B1(new_n1174), .B2(new_n1173), .C1(new_n1185), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1166), .B1(new_n1189), .B2(new_n731), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1137), .B2(new_n729), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1164), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1163), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(G375));
  AOI21_X1  g0994(.A(new_n898), .B1(new_n1091), .B2(new_n1057), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1157), .B1(new_n1195), .B2(new_n1065), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1094), .A2(new_n1048), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n975), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n718), .B1(G68), .B2(new_n1165), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G97), .A2(new_n739), .B1(new_n768), .B2(G303), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n467), .B2(new_n755), .C1(new_n923), .C2(new_n758), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G116), .A2(new_n752), .B1(new_n751), .B2(G294), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n927), .A2(new_n1202), .A3(new_n999), .A4(new_n258), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G159), .A2(new_n739), .B1(new_n768), .B2(G128), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n801), .B2(new_n758), .C1(new_n320), .C2(new_n755), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n258), .B1(new_n765), .B2(G58), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n744), .A2(G50), .B1(G132), .B2(new_n751), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n802), .C2(new_n1107), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1201), .A2(new_n1203), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1199), .B1(new_n1209), .B2(new_n731), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n728), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(new_n1049), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1094), .B2(new_n716), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1198), .A2(new_n1214), .ZN(G381));
  OR3_X1    g1015(.A1(new_n958), .A2(new_n976), .A3(new_n944), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n977), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n943), .A3(new_n1044), .ZN(new_n1218));
  OR2_X1    g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1218), .A2(G384), .A3(G381), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1122), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n1221), .A3(new_n1193), .ZN(G407));
  NAND2_X1  g1022(.A1(new_n646), .A2(G213), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1193), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G407), .A2(G213), .A3(new_n1225), .ZN(G409));
  NOR3_X1   g1026(.A1(new_n1163), .A2(new_n1221), .A3(new_n1192), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1156), .A2(new_n1158), .A3(new_n975), .A4(new_n1161), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1154), .A2(KEYINPUT123), .A3(new_n1155), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n717), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(new_n1232), .A3(new_n1191), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1233), .A2(new_n1221), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1223), .B1(new_n1227), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1065), .B(new_n1157), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1196), .B2(KEYINPUT60), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT60), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n663), .B1(new_n1197), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1236), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1197), .B1(new_n1067), .B2(new_n1239), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n667), .B1(new_n1237), .B2(KEYINPUT60), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1243), .A3(KEYINPUT124), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1245), .B2(new_n1214), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n817), .B(new_n1213), .C1(new_n1241), .C2(new_n1244), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1224), .A2(G2897), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1248), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1242), .A2(new_n1243), .A3(KEYINPUT124), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT124), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1214), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n817), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1245), .A2(G384), .A3(new_n1214), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1250), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1235), .B1(new_n1249), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT62), .B1(new_n1235), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1163), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1192), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(G378), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1233), .A2(new_n1221), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1223), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .A4(new_n1268), .ZN(new_n1269));
  XOR2_X1   g1069(.A(G393), .B(G396), .Z(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1044), .B1(new_n1217), .B2(new_n943), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n943), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1273), .B(G390), .C1(new_n1216), .C2(new_n977), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1271), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(G390), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1218), .A3(new_n1270), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1269), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1257), .A2(KEYINPUT125), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT63), .B1(new_n1235), .B2(new_n1258), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1265), .A2(new_n1266), .A3(new_n1282), .A4(new_n1223), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1285), .B(new_n1235), .C1(new_n1249), .C2(new_n1256), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1280), .A2(new_n1284), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(new_n1288), .ZN(G405));
  INV_X1    g1089(.A(KEYINPUT127), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1275), .A2(new_n1277), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1266), .A2(KEYINPUT126), .A3(new_n1263), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1258), .B1(new_n1295), .B2(new_n1227), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1193), .A2(G378), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1294), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1297), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1294), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1292), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(G402));
endmodule


