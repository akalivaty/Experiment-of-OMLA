//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n582, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n606, new_n607, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT64), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT64), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n464), .A2(KEYINPUT65), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT3), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT64), .B(G2105), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(G137), .A3(new_n463), .A4(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n475), .B2(new_n477), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n474), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n478), .A2(new_n463), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT66), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n479), .C2(G112), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n485), .A2(new_n479), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n478), .A2(G138), .A3(new_n463), .A4(new_n479), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n466), .A2(KEYINPUT4), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n470), .A2(new_n472), .A3(G138), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(KEYINPUT67), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n469), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(new_n497), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(G126), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n485), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n496), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n516), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n511), .A2(KEYINPUT68), .A3(new_n512), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n529), .A2(new_n530), .A3(G63), .A4(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n510), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n531), .B(new_n535), .C1(new_n536), .C2(new_n518), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT69), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(KEYINPUT69), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n525), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n539), .A2(new_n541), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n513), .A2(new_n517), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G89), .B1(G51), .B2(new_n534), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT70), .A4(new_n531), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n545), .A2(new_n552), .ZN(G168));
  NAND3_X1  g128(.A1(new_n529), .A2(new_n530), .A3(G64), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n515), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G90), .ZN(new_n557));
  INV_X1    g132(.A(G52), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n518), .A2(new_n557), .B1(new_n520), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(G171));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n529), .A2(new_n530), .A3(G56), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n565), .A2(new_n566), .A3(new_n515), .ZN(new_n567));
  INV_X1    g142(.A(G81), .ZN(new_n568));
  INV_X1    g143(.A(G43), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n518), .A2(new_n568), .B1(new_n520), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n561), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n562), .A2(new_n564), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n515), .B1(new_n572), .B2(KEYINPUT71), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n570), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(KEYINPUT72), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  NAND4_X1  g155(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g156(.A1(G1), .A2(G3), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND4_X1  g158(.A1(G319), .A2(G483), .A3(G661), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT73), .ZN(G188));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n527), .A2(new_n528), .ZN(new_n587));
  INV_X1    g162(.A(G65), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(G91), .A2(new_n550), .B1(new_n589), .B2(G651), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT9), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n534), .A2(new_n591), .A3(G53), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n593));
  AND2_X1   g168(.A1(KEYINPUT6), .A2(G651), .ZN(new_n594));
  NOR2_X1   g169(.A1(KEYINPUT6), .A2(G651), .ZN(new_n595));
  OAI211_X1 g170(.A(G53), .B(G543), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT9), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n592), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n593), .B1(new_n592), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n598), .B2(new_n599), .ZN(G299));
  NAND2_X1  g175(.A1(G171), .A2(KEYINPUT75), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n556), .B2(new_n559), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G301));
  AND3_X1   g180(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n552), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT76), .B1(new_n545), .B2(new_n552), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(G286));
  AND2_X1   g183(.A1(new_n529), .A2(new_n530), .ZN(new_n609));
  OAI21_X1  g184(.A(G651), .B1(new_n609), .B2(G74), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n550), .A2(G87), .B1(G49), .B2(new_n534), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G288));
  INV_X1    g187(.A(G61), .ZN(new_n613));
  INV_X1    g188(.A(G73), .ZN(new_n614));
  OAI22_X1  g189(.A1(new_n587), .A2(new_n613), .B1(new_n614), .B2(new_n510), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G651), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT77), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n613), .B1(new_n511), .B2(new_n512), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n614), .A2(new_n510), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n618), .B(G651), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n550), .A2(G86), .B1(G48), .B2(new_n534), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(G305));
  AOI22_X1  g198(.A1(new_n609), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(new_n515), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT78), .B(G85), .Z(new_n626));
  INV_X1    g201(.A(G47), .ZN(new_n627));
  OAI22_X1  g202(.A1(new_n518), .A2(new_n626), .B1(new_n520), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(G290));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n631));
  INV_X1    g206(.A(G92), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n518), .B2(new_n632), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n513), .A2(new_n517), .A3(KEYINPUT10), .A4(G92), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(G79), .A2(G543), .ZN(new_n636));
  INV_X1    g211(.A(G66), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n587), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n638), .A2(G651), .B1(G54), .B2(new_n534), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n604), .B2(G868), .ZN(G284));
  AOI21_X1  g217(.A(new_n641), .B1(new_n604), .B2(G868), .ZN(G321));
  MUX2_X1   g218(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g219(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g220(.A(new_n640), .ZN(new_n646));
  INV_X1    g221(.A(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(G860), .ZN(G148));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT79), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(G868), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT80), .Z(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(G868), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g229(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g230(.A(new_n466), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n481), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n486), .A2(G135), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n490), .A2(G123), .ZN(new_n662));
  OAI221_X1 g237(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n479), .C2(G111), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(G2096), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n665), .ZN(G156));
  XOR2_X1   g241(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n667));
  XOR2_X1   g242(.A(KEYINPUT15), .B(G2435), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2438), .ZN(new_n669));
  XOR2_X1   g244(.A(G2427), .B(G2430), .Z(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n669), .B2(new_n670), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2451), .B(G2454), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT16), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2443), .B(G2446), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n680), .A3(G14), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G401));
  INV_X1    g259(.A(KEYINPUT18), .ZN(new_n685));
  XOR2_X1   g260(.A(G2084), .B(G2090), .Z(new_n686));
  XNOR2_X1  g261(.A(G2067), .B(G2678), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(KEYINPUT17), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2100), .ZN(new_n692));
  XOR2_X1   g267(.A(G2072), .B(G2078), .Z(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n688), .B2(KEYINPUT18), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G2096), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n692), .B(new_n695), .ZN(G227));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT83), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1961), .B(G1966), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1971), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT19), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n698), .A2(new_n701), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n704), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n706), .B1(new_n704), .B2(new_n702), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(G1981), .B(G1986), .Z(new_n714));
  XNOR2_X1  g289(.A(G1991), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n713), .B(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(G229));
  NOR2_X1   g295(.A1(G29), .A2(G35), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G162), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT29), .ZN(new_n723));
  INV_X1    g298(.A(G2090), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n478), .A2(G139), .A3(new_n469), .A4(new_n463), .ZN(new_n727));
  AND2_X1   g302(.A1(G103), .A2(G2104), .ZN(new_n728));
  AOI21_X1  g303(.A(KEYINPUT25), .B1(new_n479), .B2(new_n728), .ZN(new_n729));
  AND4_X1   g304(.A1(KEYINPUT25), .A2(new_n470), .A3(new_n472), .A4(new_n728), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n470), .A2(new_n472), .A3(new_n728), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n479), .A2(KEYINPUT25), .A3(new_n728), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n737), .A2(new_n738), .A3(new_n727), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n656), .A2(G127), .ZN(new_n741));
  NAND2_X1  g316(.A1(G115), .A2(G2104), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n479), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n726), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  AOI211_X1 g320(.A(KEYINPUT91), .B(new_n743), .C1(new_n732), .C2(new_n739), .ZN(new_n746));
  OAI21_X1  g321(.A(G29), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G33), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(G29), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n725), .B1(new_n749), .B2(G2072), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G2072), .B2(new_n749), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n579), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n752), .B2(G19), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(G1341), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(G1341), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n752), .A2(G4), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n646), .B2(new_n752), .ZN(new_n759));
  INV_X1    g334(.A(G1348), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n486), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n490), .A2(G128), .ZN(new_n766));
  OAI221_X1 g341(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n479), .C2(G116), .ZN(new_n767));
  AND3_X1   g342(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n764), .B1(new_n768), .B2(new_n762), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n756), .A2(new_n757), .A3(new_n761), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G11), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  INV_X1    g352(.A(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n782), .B2(KEYINPUT24), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(KEYINPUT24), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n483), .B2(new_n762), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n781), .B1(new_n664), .B2(new_n762), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n752), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n752), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1961), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n787), .B(new_n790), .C1(new_n786), .C2(new_n785), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n762), .A2(G32), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n490), .A2(G129), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT26), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n481), .A2(G105), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n486), .A2(G141), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(KEYINPUT92), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n486), .A2(new_n800), .A3(G141), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n797), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n792), .B1(new_n802), .B2(new_n762), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT27), .B(G1996), .Z(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n762), .A2(G27), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G164), .B2(new_n762), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2078), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n803), .B2(new_n804), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n752), .A2(G20), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G299), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n752), .ZN(new_n814));
  INV_X1    g389(.A(G1956), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n791), .A2(new_n805), .A3(new_n809), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(G16), .A2(G21), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G168), .B2(G16), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT93), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT94), .B(G1966), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n751), .A2(new_n774), .A3(new_n775), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n752), .A2(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n752), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G1971), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n752), .A2(G23), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G288), .B2(G16), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT33), .B(G1976), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n827), .A2(G1971), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n828), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  MUX2_X1   g411(.A(G6), .B(G305), .S(G16), .Z(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT32), .B(G1981), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n752), .A2(G24), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n629), .B2(new_n752), .ZN(new_n844));
  INV_X1    g419(.A(G1986), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n762), .A2(G25), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n486), .A2(G131), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n490), .A2(G119), .ZN(new_n849));
  OAI221_X1 g424(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n479), .C2(G107), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n847), .B1(new_n852), .B2(new_n762), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G1991), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n842), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT88), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n841), .B2(new_n840), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(KEYINPUT36), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(KEYINPUT36), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n825), .B1(new_n860), .B2(new_n861), .ZN(G311));
  AND3_X1   g437(.A1(new_n751), .A2(new_n775), .A3(new_n824), .ZN(new_n863));
  INV_X1    g438(.A(new_n861), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n863), .B(new_n774), .C1(new_n864), .C2(new_n859), .ZN(G150));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n867));
  INV_X1    g442(.A(G93), .ZN(new_n868));
  INV_X1    g443(.A(G55), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n518), .A2(new_n868), .B1(new_n520), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n529), .A2(new_n530), .A3(G67), .ZN(new_n871));
  INV_X1    g446(.A(G80), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n510), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n873), .B2(G651), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n866), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(KEYINPUT97), .B(new_n874), .C1(new_n567), .C2(new_n570), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n571), .A2(new_n577), .A3(new_n875), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n640), .A2(new_n647), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT38), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n883), .B(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT99), .Z(new_n888));
  AOI21_X1  g463(.A(G860), .B1(new_n886), .B2(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n875), .A2(G860), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n891), .B(KEYINPUT37), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(G145));
  XNOR2_X1  g468(.A(new_n664), .B(new_n483), .ZN(new_n894));
  XOR2_X1   g469(.A(G162), .B(new_n894), .Z(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n799), .A2(new_n801), .ZN(new_n897));
  OAI22_X1  g472(.A1(new_n745), .A2(new_n746), .B1(new_n897), .B2(new_n797), .ZN(new_n898));
  INV_X1    g473(.A(new_n739), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n738), .B1(new_n737), .B2(new_n727), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n744), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT91), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n740), .A2(new_n726), .A3(new_n744), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n802), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n479), .B2(G118), .ZN(new_n906));
  INV_X1    g481(.A(G118), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n473), .A2(KEYINPUT100), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n478), .A2(new_n473), .A3(G130), .A4(new_n463), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n478), .A2(G142), .A3(new_n469), .A4(new_n463), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT101), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n911), .A2(new_n917), .A3(new_n913), .A4(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n658), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n918), .A3(new_n658), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n898), .A2(new_n904), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n898), .B2(new_n904), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n768), .A2(G164), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n494), .A2(new_n495), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n485), .ZN(new_n931));
  INV_X1    g506(.A(new_n506), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n931), .A2(new_n932), .B1(new_n504), .B2(new_n501), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n851), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n926), .A2(new_n851), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n924), .A2(new_n925), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n938), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(new_n936), .ZN(new_n942));
  INV_X1    g517(.A(new_n923), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n902), .A2(new_n802), .A3(new_n903), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n802), .B1(new_n902), .B2(new_n903), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n898), .A2(new_n904), .A3(new_n923), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n896), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n939), .B1(new_n924), .B2(new_n925), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n942), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n895), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT102), .B(G37), .Z(new_n954));
  AOI21_X1  g529(.A(KEYINPUT103), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n957));
  INV_X1    g532(.A(new_n954), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n957), .B(new_n958), .C1(new_n949), .C2(new_n952), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g537(.A1(new_n646), .A2(G299), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n592), .A2(new_n597), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT74), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n592), .A2(new_n597), .A3(new_n593), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n640), .A3(new_n968), .A4(new_n590), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT104), .B1(new_n646), .B2(G299), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(KEYINPUT105), .A3(KEYINPUT41), .A4(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(KEYINPUT41), .A3(new_n963), .A4(new_n969), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT41), .ZN(new_n976));
  INV_X1    g551(.A(new_n971), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n963), .A2(new_n969), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n972), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n883), .A2(new_n650), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n651), .B1(new_n881), .B2(new_n882), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(G303), .B(G288), .Z(new_n985));
  NAND2_X1  g560(.A1(new_n629), .A2(G305), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n629), .A2(G305), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT42), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n970), .A2(new_n971), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n981), .A2(new_n993), .A3(new_n982), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n984), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n984), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g571(.A(G868), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G868), .B2(new_n874), .ZN(G295));
  OAI21_X1  g573(.A(new_n997), .B1(G868), .B2(new_n874), .ZN(G331));
  AND3_X1   g574(.A1(new_n989), .A2(KEYINPUT106), .A3(new_n990), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT106), .B1(new_n989), .B2(new_n990), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT76), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G168), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n552), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(G171), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G168), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n604), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n881), .B2(new_n882), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n878), .A2(new_n880), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT98), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n878), .A2(new_n880), .A3(new_n879), .ZN(new_n1012));
  AOI22_X1  g587(.A1(G286), .A2(G171), .B1(G168), .B2(G301), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1009), .A2(new_n1014), .A3(new_n993), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n979), .A2(new_n973), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1002), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n980), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n881), .A2(new_n1008), .A3(new_n882), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1013), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1009), .A2(new_n1014), .A3(new_n993), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n991), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1018), .A2(new_n1024), .A3(new_n1025), .A4(new_n954), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n980), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1002), .B1(new_n1015), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G37), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1024), .A3(new_n1029), .ZN(new_n1030));
  AOI22_X1  g605(.A1(KEYINPUT107), .A2(new_n1026), .B1(new_n1030), .B2(KEYINPUT43), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1015), .A2(new_n1027), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n958), .B1(new_n1033), .B2(new_n991), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n1025), .A4(new_n1018), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1031), .A2(new_n1032), .A3(new_n1036), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1030), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT108), .B1(new_n1030), .B2(KEYINPUT43), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1018), .A2(new_n1024), .A3(new_n954), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT43), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1038), .B(new_n1039), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(KEYINPUT44), .B2(new_n1045), .ZN(G397));
  NAND2_X1  g621(.A1(G303), .A2(G8), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT55), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  INV_X1    g624(.A(G1384), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n496), .B2(new_n507), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n474), .A2(G40), .A3(new_n480), .A4(new_n482), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n934), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n1050), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT113), .B(G1971), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n934), .A2(new_n1060), .A3(new_n1050), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1051), .A2(KEYINPUT50), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1054), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n724), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(KEYINPUT117), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G8), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT117), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1048), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G8), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1069), .B(new_n1048), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1384), .B1(new_n930), .B2(new_n933), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1063), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n610), .A2(new_n611), .A3(G1976), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(G8), .A4(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(G8), .B(new_n1075), .C1(new_n1051), .C2(new_n1054), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT52), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1072), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(new_n1069), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n550), .A2(G86), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n534), .A2(G48), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n621), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n618), .B1(new_n615), .B2(G651), .ZN(new_n1085));
  OAI21_X1  g660(.A(G1981), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n1089));
  INV_X1    g664(.A(G1981), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n617), .A2(new_n1090), .A3(new_n621), .A4(new_n622), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1082), .A2(new_n621), .A3(new_n1083), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(KEYINPUT114), .A3(new_n1090), .A4(new_n617), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1088), .A2(new_n1089), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1081), .B1(new_n1096), .B2(KEYINPUT49), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1098), .A2(KEYINPUT49), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1079), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1070), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1068), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1071), .A2(KEYINPUT45), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1055), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n821), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1061), .A2(new_n1062), .A3(new_n786), .A4(new_n1063), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(G168), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1108), .A2(new_n1109), .A3(G8), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1007), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(G8), .A3(new_n1108), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1113), .B2(KEYINPUT51), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1103), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G2078), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1055), .A2(new_n1104), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1055), .A2(new_n1104), .A3(KEYINPUT121), .A4(new_n1116), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(KEYINPUT53), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1116), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  INV_X1    g698(.A(G1961), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1122), .A2(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n604), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT110), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT45), .B1(new_n1051), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1071), .A2(KEYINPUT110), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1054), .A2(new_n1123), .A3(G2078), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n1053), .A3(new_n1056), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1126), .A2(G301), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1128), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1121), .A2(new_n1126), .A3(G301), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1126), .A2(new_n1134), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1139), .B2(G171), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1125), .A2(new_n815), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n813), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n590), .A2(new_n1143), .A3(new_n964), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT56), .B(G2072), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1142), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1051), .A2(G2067), .A3(new_n1054), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1125), .B2(new_n760), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n640), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1146), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n646), .B(new_n1150), .C1(new_n1125), .C2(new_n760), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT60), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT119), .B(G1996), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT58), .B(G1341), .Z(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1072), .A2(KEYINPUT120), .A3(new_n1159), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1158), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n579), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT60), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1151), .A2(new_n1168), .A3(new_n646), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1164), .A2(KEYINPUT59), .A3(new_n579), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1156), .A2(new_n1167), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1173), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1142), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1153), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1154), .B1(new_n1171), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1115), .A2(new_n1141), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(G8), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1048), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1069), .B(G286), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1102), .A2(new_n1183), .A3(KEYINPUT63), .A4(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1068), .A2(new_n1102), .A3(new_n1184), .ZN(new_n1186));
  XOR2_X1   g761(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1187));
  OAI21_X1  g762(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT49), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1096), .A2(KEYINPUT49), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(new_n1192), .A3(new_n1081), .ZN(new_n1193));
  NOR2_X1   g768(.A1(G288), .A2(G1976), .ZN(new_n1194));
  AOI22_X1  g769(.A1(new_n1193), .A2(new_n1194), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1081), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1048), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1181), .A2(G8), .A3(new_n1197), .ZN(new_n1198));
  OAI22_X1  g773(.A1(new_n1195), .A2(new_n1196), .B1(new_n1198), .B2(new_n1101), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT116), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT116), .ZN(new_n1201));
  OAI221_X1 g776(.A(new_n1201), .B1(new_n1198), .B2(new_n1101), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1180), .A2(new_n1188), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(KEYINPUT122), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1180), .A2(new_n1188), .A3(new_n1206), .A4(new_n1203), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1114), .B(KEYINPUT62), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1103), .A2(new_n1128), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1205), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1130), .A2(new_n1131), .A3(new_n1063), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(G1996), .ZN(new_n1214));
  AOI21_X1  g789(.A(KEYINPUT111), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT111), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1212), .A2(new_n1216), .A3(G1996), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n802), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n927), .B(new_n770), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(new_n1214), .B2(new_n802), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1220), .A2(new_n1213), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n851), .B(new_n854), .ZN(new_n1222));
  OAI211_X1 g797(.A(new_n1218), .B(new_n1221), .C1(new_n1212), .C2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g798(.A(new_n629), .B(new_n845), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1223), .B1(new_n1213), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1211), .A2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g801(.A1(new_n1218), .A2(new_n854), .A3(new_n852), .A4(new_n1221), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n768), .A2(new_n770), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1212), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AND2_X1   g804(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1231));
  OR2_X1    g806(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n1233));
  NOR3_X1   g808(.A1(new_n1212), .A2(G1986), .A3(G290), .ZN(new_n1234));
  XNOR2_X1  g809(.A(new_n1234), .B(KEYINPUT48), .ZN(new_n1235));
  OR2_X1    g810(.A1(new_n1223), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g811(.A(new_n1212), .B1(new_n802), .B2(new_n1219), .ZN(new_n1237));
  XOR2_X1   g812(.A(new_n1237), .B(KEYINPUT124), .Z(new_n1238));
  OR3_X1    g813(.A1(new_n1215), .A2(KEYINPUT46), .A3(new_n1217), .ZN(new_n1239));
  OAI21_X1  g814(.A(KEYINPUT46), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g816(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1242));
  XNOR2_X1  g817(.A(new_n1241), .B(new_n1242), .ZN(new_n1243));
  NAND4_X1  g818(.A1(new_n1232), .A2(new_n1233), .A3(new_n1236), .A4(new_n1243), .ZN(new_n1244));
  OAI211_X1 g819(.A(new_n1243), .B(new_n1236), .C1(new_n1231), .C2(new_n1230), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1245), .A2(KEYINPUT126), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1226), .A2(new_n1247), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g823(.A(KEYINPUT127), .ZN(new_n1250));
  NOR2_X1   g824(.A1(G227), .A2(new_n459), .ZN(new_n1251));
  AND3_X1   g825(.A1(new_n719), .A2(new_n683), .A3(new_n1251), .ZN(new_n1252));
  OAI21_X1  g826(.A(new_n1252), .B1(new_n955), .B2(new_n959), .ZN(new_n1253));
  AOI211_X1 g827(.A(new_n1250), .B(new_n1253), .C1(new_n1031), .C2(new_n1036), .ZN(new_n1254));
  NAND2_X1  g828(.A1(new_n1030), .A2(KEYINPUT43), .ZN(new_n1255));
  NAND2_X1  g829(.A1(new_n1026), .A2(KEYINPUT107), .ZN(new_n1256));
  NAND3_X1  g830(.A1(new_n1036), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g831(.A(new_n1253), .ZN(new_n1258));
  AOI21_X1  g832(.A(KEYINPUT127), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g833(.A1(new_n1254), .A2(new_n1259), .ZN(G308));
  NAND2_X1  g834(.A1(new_n1257), .A2(new_n1258), .ZN(G225));
endmodule


