//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT84), .A2(G8gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n204), .B(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT84), .A2(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT14), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT81), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G43gat), .A2(G50gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G43gat), .A2(G50gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT15), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n216), .ZN(new_n222));
  NOR2_X1   g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT14), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n215), .A2(new_n219), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n216), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT81), .B(new_n213), .C1(new_n223), .C2(KEYINPUT14), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT14), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT15), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT82), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n225), .A2(new_n235), .A3(new_n229), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n225), .B2(new_n229), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n234), .B1(new_n238), .B2(new_n231), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(KEYINPUT82), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n229), .A3(new_n235), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n240), .A2(new_n234), .A3(new_n231), .A4(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n209), .B(new_n233), .C1(new_n239), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n208), .A2(new_n238), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n244), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n246), .B(KEYINPUT13), .Z(new_n248));
  INV_X1    g047(.A(new_n245), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n208), .A2(new_n238), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT18), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT11), .ZN(new_n258));
  INV_X1    g057(.A(G169gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G197gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n252), .B(new_n255), .C1(new_n256), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n256), .A3(new_n251), .ZN(new_n264));
  INV_X1    g063(.A(new_n262), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n251), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n240), .A2(new_n231), .A3(new_n241), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT83), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n232), .B1(new_n268), .B2(new_n242), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n249), .B1(new_n269), .B2(new_n209), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT18), .B1(new_n270), .B2(new_n246), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n274), .B1(KEYINPUT23), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT25), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT24), .ZN(new_n281));
  NOR2_X1   g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI211_X1 g082(.A(new_n276), .B(new_n279), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT65), .B(G176gat), .Z(new_n285));
  NOR2_X1   g084(.A1(new_n278), .A2(G169gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT66), .B1(new_n287), .B2(new_n276), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n276), .B1(new_n285), .B2(new_n286), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n282), .B(KEYINPUT64), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n281), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n284), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT27), .B(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT28), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n277), .A2(KEYINPUT68), .A3(KEYINPUT26), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n274), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n275), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT68), .B1(new_n277), .B2(KEYINPUT26), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n280), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n309), .B(KEYINPUT69), .Z(new_n310));
  NAND2_X1  g109(.A1(new_n296), .A2(new_n297), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n298), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G113gat), .B(G120gat), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n313), .A2(KEYINPUT1), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G227gat), .ZN(new_n318));
  INV_X1    g117(.A(G233gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n314), .B(new_n315), .Z(new_n321));
  NAND4_X1  g120(.A1(new_n298), .A2(new_n310), .A3(new_n321), .A4(new_n311), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT32), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT33), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G15gat), .B(G43gat), .Z(new_n327));
  XNOR2_X1  g126(.A(G71gat), .B(G99gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n323), .B(KEYINPUT32), .C1(new_n325), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n320), .B1(new_n317), .B2(new_n322), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT34), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI211_X1 g135(.A(KEYINPUT34), .B(new_n320), .C1(new_n317), .C2(new_n322), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340));
  XNOR2_X1  g139(.A(G197gat), .B(G204gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT71), .B(G218gat), .ZN(new_n342));
  INV_X1    g141(.A(G211gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT70), .B(KEYINPUT22), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G211gat), .B(G218gat), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n340), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT3), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n357));
  INV_X1    g156(.A(G141gat), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n358), .A2(G148gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(G148gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G155gat), .ZN(new_n362));
  INV_X1    g161(.A(G162gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT73), .B(G148gat), .Z(new_n368));
  AOI21_X1  g167(.A(new_n359), .B1(new_n368), .B2(G141gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n364), .B1(new_n357), .B2(new_n365), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n350), .A2(new_n348), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(KEYINPUT72), .ZN(new_n379));
  INV_X1    g178(.A(new_n376), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n340), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n372), .B1(new_n382), .B2(new_n375), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n373), .A2(new_n378), .B1(new_n374), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT77), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G50gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n387), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G22gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n385), .B(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n336), .A2(new_n337), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n330), .A3(new_n332), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n339), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n296), .A2(new_n309), .ZN(new_n397));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n340), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n312), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n401), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n312), .B2(new_n398), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n379), .A2(new_n402), .B1(new_n404), .B2(new_n377), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n405), .A2(new_n410), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n377), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n312), .A2(new_n401), .ZN(new_n414));
  INV_X1    g213(.A(new_n399), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n379), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n416), .A3(new_n410), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT30), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n411), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n372), .A2(new_n375), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n321), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n316), .A2(new_n372), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n422), .B(new_n425), .C1(new_n423), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n429), .A2(KEYINPUT5), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n423), .B2(new_n426), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(new_n422), .C1(new_n424), .C2(new_n423), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n321), .A2(new_n371), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n423), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n429), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(KEYINPUT5), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(G57gat), .B(G85gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  NAND3_X1  g240(.A1(new_n431), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n431), .B2(new_n437), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n443), .B(new_n441), .C1(new_n431), .C2(new_n437), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n419), .A2(new_n449), .ZN(new_n450));
  OR3_X1    g249(.A1(new_n396), .A2(new_n450), .A3(KEYINPUT35), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n452));
  AND4_X1   g251(.A1(new_n406), .A2(new_n413), .A3(new_n416), .A4(new_n410), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n406), .B1(new_n405), .B2(new_n410), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n413), .A2(new_n416), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n409), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n452), .B1(new_n457), .B2(new_n448), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n419), .A2(KEYINPUT75), .A3(new_n449), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n396), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT35), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n451), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n395), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n394), .B1(new_n332), .B2(new_n330), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT36), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n339), .A2(new_n466), .A3(new_n395), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n393), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n458), .A2(new_n469), .A3(new_n459), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n427), .A2(new_n429), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n471), .A2(KEYINPUT39), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n471), .B(KEYINPUT39), .C1(new_n429), .C2(new_n435), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n441), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n474), .A2(KEYINPUT80), .A3(new_n475), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n472), .A2(new_n473), .A3(new_n441), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n445), .B1(new_n480), .B2(KEYINPUT40), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n457), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n410), .B1(new_n405), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n402), .A2(new_n379), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n404), .A2(new_n377), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT37), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n455), .B2(KEYINPUT37), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n488), .A2(new_n489), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n448), .A2(new_n417), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n482), .B(new_n393), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n470), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n273), .B1(new_n462), .B2(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G183gat), .B(G211gat), .Z(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT88), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(G57gat), .A2(G64gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(G57gat), .A2(G64gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n500), .B(new_n501), .C1(new_n503), .C2(KEYINPUT9), .ZN(new_n504));
  NOR2_X1   g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT86), .B1(new_n503), .B2(new_n505), .ZN(new_n508));
  INV_X1    g307(.A(G71gat), .ZN(new_n509));
  INV_X1    g308(.A(G78gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT86), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n502), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(new_n515), .A3(new_n504), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n514), .B2(new_n504), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n507), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g319(.A1(G231gat), .A2(G233gat), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  XNOR2_X1  g322(.A(G127gat), .B(G155gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n522), .B2(new_n523), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n499), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n527), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n525), .A3(new_n498), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n208), .B1(new_n519), .B2(KEYINPUT21), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n528), .B2(new_n530), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n496), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n531), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(new_n538));
  INV_X1    g337(.A(new_n496), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n542));
  AND3_X1   g341(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544));
  INV_X1    g343(.A(G85gat), .ZN(new_n545));
  INV_X1    g344(.A(G92gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(KEYINPUT8), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  NAND3_X1  g348(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n551), .B(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n543), .B1(new_n238), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT89), .ZN(new_n556));
  INV_X1    g355(.A(new_n554), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n269), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n542), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(KEYINPUT90), .A3(new_n561), .ZN(new_n566));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n569), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n542), .B(new_n571), .C1(new_n562), .C2(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n541), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(KEYINPUT91), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(new_n541), .B2(new_n573), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT92), .ZN(new_n578));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n518), .A2(new_n557), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n554), .B(new_n507), .C1(new_n517), .C2(new_n516), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n554), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n581), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n589), .A2(new_n590), .A3(new_n581), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n578), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(KEYINPUT92), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n575), .A2(new_n577), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n495), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n599), .A2(new_n449), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT93), .B(G1gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(G1324gat));
  INV_X1    g401(.A(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n457), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT16), .B(G8gat), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(KEYINPUT42), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT42), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n604), .B2(G8gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n608), .B1(new_n607), .B2(new_n610), .ZN(G1325gat));
  OAI21_X1  g410(.A(G15gat), .B1(new_n599), .B2(new_n468), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n339), .A2(new_n395), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n613), .A2(G15gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n599), .B2(new_n614), .ZN(G1326gat));
  NAND2_X1  g414(.A1(new_n603), .A2(new_n469), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT94), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT43), .B(G22gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(G1327gat));
  INV_X1    g418(.A(new_n541), .ZN(new_n620));
  INV_X1    g419(.A(new_n573), .ZN(new_n621));
  INV_X1    g420(.A(new_n597), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT95), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n495), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n210), .A3(new_n448), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT45), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n458), .A2(new_n459), .ZN(new_n629));
  INV_X1    g428(.A(new_n396), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n461), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n396), .A2(new_n450), .A3(KEYINPUT35), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n451), .B(KEYINPUT99), .C1(new_n460), .C2(new_n461), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n470), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT98), .A4(new_n469), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n636), .A2(new_n468), .A3(new_n493), .A4(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n640), .A3(new_n621), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n573), .B1(new_n462), .B2(new_n494), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n630), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n632), .B1(new_n645), .B2(KEYINPUT35), .ZN(new_n646));
  INV_X1    g445(.A(new_n487), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n409), .B1(new_n455), .B2(KEYINPUT37), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n489), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n484), .A2(new_n490), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n492), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n481), .A2(new_n478), .A3(new_n479), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n393), .B1(new_n419), .B2(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n465), .B(new_n467), .C1(new_n651), .C2(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n458), .A2(new_n469), .A3(new_n459), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n621), .B1(new_n646), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(KEYINPUT97), .A3(KEYINPUT44), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n644), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n597), .A2(KEYINPUT96), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n597), .A2(KEYINPUT96), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n663), .A2(new_n541), .A3(new_n273), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n659), .A2(new_n448), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n627), .B1(new_n210), .B2(new_n665), .ZN(G1328gat));
  NAND3_X1  g465(.A1(new_n659), .A2(new_n457), .A3(new_n664), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n211), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(new_n668), .B2(new_n667), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n625), .A2(new_n211), .A3(new_n457), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT46), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(G1329gat));
  INV_X1    g472(.A(new_n468), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n674), .A3(new_n664), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n613), .A2(G43gat), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n675), .A2(G43gat), .B1(new_n625), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT47), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1330gat));
  NOR2_X1   g480(.A1(new_n393), .A2(G50gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n625), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT104), .Z(new_n685));
  NAND3_X1  g484(.A1(new_n659), .A2(new_n469), .A3(new_n664), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(G50gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(KEYINPUT48), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n684), .B(KEYINPUT103), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(G50gat), .B2(new_n686), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n690), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g490(.A1(new_n575), .A2(new_n577), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n273), .A3(new_n663), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n639), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n449), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT106), .B(G57gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1332gat));
  NAND3_X1  g497(.A1(new_n694), .A2(new_n457), .A3(new_n639), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  AND2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n700), .B2(new_n699), .ZN(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n695), .B2(new_n468), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n339), .A2(new_n509), .A3(new_n395), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n695), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g506(.A1(new_n695), .A2(new_n393), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(new_n510), .ZN(G1335gat));
  NOR3_X1   g508(.A1(new_n449), .A2(G85gat), .A3(new_n622), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n263), .A2(new_n272), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n541), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n639), .A2(new_n621), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n639), .A2(KEYINPUT51), .A3(new_n621), .A4(new_n712), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n715), .A2(KEYINPUT108), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT108), .B1(new_n715), .B2(new_n716), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n710), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n541), .A2(new_n711), .A3(new_n622), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n659), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n659), .B2(new_n720), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n721), .A2(new_n722), .A3(new_n449), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n723), .B2(new_n545), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT109), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n726), .B(new_n719), .C1(new_n723), .C2(new_n545), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1336gat));
  NAND2_X1  g527(.A1(new_n715), .A2(new_n716), .ZN(new_n729));
  AND4_X1   g528(.A1(new_n546), .A2(new_n729), .A3(new_n457), .A4(new_n663), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(KEYINPUT52), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n659), .A2(new_n720), .ZN(new_n732));
  OAI21_X1  g531(.A(G92gat), .B1(new_n732), .B2(new_n419), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n722), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n659), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n457), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n730), .B1(new_n737), .B2(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(G1337gat));
  NOR3_X1   g539(.A1(new_n613), .A2(G99gat), .A3(new_n622), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT110), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n717), .B2(new_n718), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n721), .A2(new_n722), .A3(new_n468), .ZN(new_n744));
  INV_X1    g543(.A(G99gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(G1338gat));
  OAI21_X1  g545(.A(G106gat), .B1(new_n732), .B2(new_n393), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n662), .A2(new_n393), .A3(G106gat), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT53), .B1(new_n729), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n469), .A3(new_n736), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n748), .B(KEYINPUT111), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G106gat), .B1(new_n729), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(G1339gat));
  NOR4_X1   g554(.A1(new_n575), .A2(new_n577), .A3(new_n711), .A4(new_n597), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n587), .A2(new_n588), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n582), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n587), .A2(new_n588), .A3(new_n583), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n759), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n581), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n589), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n589), .A2(new_n763), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT112), .B1(new_n766), .B2(new_n760), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n757), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n759), .A2(KEYINPUT54), .A3(new_n760), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n771), .A2(KEYINPUT55), .A3(new_n761), .A4(new_n764), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n768), .A2(new_n595), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n255), .A2(new_n251), .A3(new_n247), .A4(new_n262), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n270), .A2(new_n246), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n249), .A2(new_n250), .A3(new_n248), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n261), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n572), .A2(new_n570), .A3(new_n773), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n597), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n768), .A2(new_n595), .A3(new_n772), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n273), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n773), .A2(new_n711), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n785), .A3(new_n780), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n779), .B1(new_n787), .B2(new_n573), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n541), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n621), .B1(new_n783), .B2(new_n786), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n791), .B2(new_n779), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n756), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n457), .A2(new_n449), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n630), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n711), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G113gat), .ZN(G1340gat));
  INV_X1    g599(.A(G120gat), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n797), .A2(new_n801), .A3(new_n662), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n597), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n801), .B2(new_n803), .ZN(G1341gat));
  NOR2_X1   g603(.A1(new_n797), .A2(new_n620), .ZN(new_n805));
  XNOR2_X1  g604(.A(KEYINPUT115), .B(G127gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1342gat));
  AOI21_X1  g606(.A(new_n573), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n796), .A2(new_n630), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(new_n809), .B(KEYINPUT116), .Z(new_n810));
  NOR2_X1   g609(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(G1343gat));
  NOR2_X1   g611(.A1(new_n674), .A2(new_n795), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n788), .A2(new_n789), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n792), .A3(new_n620), .ZN(new_n816));
  INV_X1    g615(.A(new_n756), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n393), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(KEYINPUT57), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n782), .B(KEYINPUT118), .Z(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n573), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n620), .B1(new_n822), .B2(new_n779), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n817), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n393), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n819), .A2(KEYINPUT117), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n818), .B2(KEYINPUT57), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n814), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n358), .B1(new_n830), .B2(new_n711), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n674), .A2(new_n393), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n796), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n711), .A2(new_n358), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT119), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT58), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n835), .A2(KEYINPUT58), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n831), .B2(new_n837), .ZN(G1344gat));
  XOR2_X1   g637(.A(new_n813), .B(KEYINPUT120), .Z(new_n839));
  OAI21_X1  g638(.A(KEYINPUT57), .B1(new_n793), .B2(new_n393), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n621), .B2(new_n773), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n573), .A2(KEYINPUT121), .A3(new_n781), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n778), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n541), .B1(new_n821), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n825), .B(new_n469), .C1(new_n845), .C2(new_n756), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n839), .A2(new_n840), .A3(new_n597), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n848));
  INV_X1    g647(.A(new_n833), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n368), .A3(new_n597), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n368), .B1(new_n830), .B2(new_n597), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n848), .B(new_n850), .C1(new_n851), .C2(KEYINPUT59), .ZN(G1345gat));
  NAND2_X1  g651(.A1(new_n827), .A2(new_n829), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n813), .ZN(new_n854));
  OAI21_X1  g653(.A(G155gat), .B1(new_n854), .B2(new_n620), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n362), .A3(new_n541), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1346gat));
  OAI21_X1  g656(.A(G162gat), .B1(new_n854), .B2(new_n573), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n833), .A2(G162gat), .A3(new_n573), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n363), .B1(new_n830), .B2(new_n621), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT122), .B1(new_n863), .B2(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1347gat));
  INV_X1    g664(.A(new_n793), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n419), .A2(new_n448), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n396), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n273), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(new_n259), .ZN(G1348gat));
  NOR2_X1   g671(.A1(new_n870), .A2(new_n622), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n662), .A2(new_n285), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n873), .A2(G176gat), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT123), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n870), .A2(new_n620), .ZN(new_n877));
  MUX2_X1   g676(.A(G183gat), .B(new_n299), .S(new_n877), .Z(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g678(.A1(new_n866), .A2(new_n621), .A3(new_n869), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G190gat), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT61), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(G190gat), .B2(new_n880), .ZN(G1351gat));
  NOR2_X1   g682(.A1(new_n674), .A2(new_n868), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n818), .A2(new_n884), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n885), .A2(G197gat), .A3(new_n273), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n840), .A2(new_n846), .A3(new_n884), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n273), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G197gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n887), .A3(new_n273), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(G1352gat));
  OAI21_X1  g691(.A(G204gat), .B1(new_n888), .B2(new_n662), .ZN(new_n893));
  OR3_X1    g692(.A1(new_n885), .A2(G204gat), .A3(new_n622), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n894), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT125), .B1(new_n894), .B2(KEYINPUT62), .ZN(new_n896));
  OAI221_X1 g695(.A(new_n893), .B1(KEYINPUT62), .B2(new_n894), .C1(new_n895), .C2(new_n896), .ZN(G1353gat));
  NAND4_X1  g696(.A1(new_n818), .A2(new_n343), .A3(new_n541), .A4(new_n884), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n840), .A2(new_n541), .A3(new_n846), .A4(new_n884), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT63), .B1(new_n899), .B2(G211gat), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT126), .B(KEYINPUT63), .C1(new_n899), .C2(G211gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(KEYINPUT127), .B(new_n898), .C1(new_n903), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1354gat));
  NOR2_X1   g708(.A1(new_n885), .A2(new_n573), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n573), .A2(new_n342), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n910), .A2(G218gat), .B1(new_n888), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(G1355gat));
endmodule


