//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n201), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n206), .A2(new_n207), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n211), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n221), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n213), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n201), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT65), .B(G50), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT69), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT69), .ZN(new_n252));
  NAND4_X1  g0052(.A1(new_n252), .A2(new_n249), .A3(G13), .A4(G20), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n223), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n249), .A2(G20), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G50), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n251), .A2(new_n253), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(G50), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n256), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT68), .A2(G58), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n224), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(new_n266), .B1(G150), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n208), .A2(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OR3_X1    g0070(.A1(new_n261), .A2(KEYINPUT9), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT9), .B1(new_n261), .B2(new_n270), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  OAI211_X1 g0074(.A(G1), .B(G13), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n277), .A4(G274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n277), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G226), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n289), .A2(G223), .B1(new_n292), .B2(G77), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1698), .B1(new_n287), .B2(new_n288), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G222), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n282), .B(new_n285), .C1(new_n296), .C2(new_n275), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n271), .A2(new_n272), .B1(G200), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n298), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n261), .A2(new_n270), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n297), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT70), .B(G179), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n311), .B2(new_n297), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n289), .A2(G238), .B1(new_n292), .B2(G107), .ZN(new_n313));
  INV_X1    g0113(.A(new_n294), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n213), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n283), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n284), .A2(G244), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n282), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n310), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n265), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G77), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(new_n256), .B1(new_n326), .B2(new_n254), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n257), .A2(G77), .A3(new_n258), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n318), .A2(new_n308), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n320), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT71), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n319), .A2(G190), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n329), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(KEYINPUT71), .B1(G200), .B2(new_n318), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n306), .A2(new_n312), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n280), .A2(KEYINPUT73), .A3(new_n281), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G97), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n213), .A2(G1698), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G226), .B2(G1698), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n339), .B1(new_n341), .B2(new_n292), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n283), .B1(new_n284), .B2(G238), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT73), .B1(new_n280), .B2(new_n281), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT13), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n345), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n347), .A2(new_n348), .A3(new_n338), .A4(new_n343), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n344), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n348), .A4(new_n347), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(G169), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT14), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n351), .A2(new_n356), .A3(G169), .A4(new_n353), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n346), .A2(new_n349), .A3(G179), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n254), .A2(new_n202), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT12), .ZN(new_n361));
  INV_X1    g0161(.A(new_n267), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n207), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n265), .A2(new_n326), .B1(new_n224), .B2(G68), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n256), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT11), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n257), .A2(G68), .A3(new_n258), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n346), .A2(G190), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n370), .B2(new_n349), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n351), .A2(G200), .A3(new_n353), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n264), .A2(new_n258), .ZN(new_n375));
  INV_X1    g0175(.A(new_n264), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n257), .A2(new_n375), .B1(new_n254), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT3), .B(G33), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n379), .A2(new_n380), .A3(G20), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n292), .B2(new_n224), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(G20), .B1(G159), .B2(new_n267), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n262), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n378), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G226), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G1698), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(G223), .B2(G1698), .ZN(new_n393));
  INV_X1    g0193(.A(G87), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n292), .B1(new_n273), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n283), .B1(G232), .B2(new_n284), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n282), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G200), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(G190), .A3(new_n282), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n390), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g0202(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n390), .A2(new_n400), .A3(KEYINPUT75), .A4(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n397), .A2(new_n308), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n396), .A2(new_n282), .A3(new_n310), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT18), .B1(new_n390), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n388), .A2(new_n389), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n377), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  INV_X1    g0212(.A(new_n408), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n404), .A2(new_n405), .A3(new_n409), .A4(new_n414), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n337), .A2(new_n374), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n254), .A2(new_n214), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n249), .A2(G33), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n260), .A2(new_n262), .A3(G97), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g0220(.A(G97), .B(G107), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT6), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n422), .A2(new_n214), .A3(G107), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n427));
  OAI21_X1  g0227(.A(G107), .B1(new_n381), .B2(new_n382), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n420), .B1(new_n429), .B2(new_n256), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n276), .A2(G1), .ZN(new_n431));
  AND2_X1   g0231(.A1(KEYINPUT5), .A2(G41), .ZN(new_n432));
  NOR2_X1   g0232(.A1(KEYINPUT5), .A2(G41), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(G257), .A3(new_n275), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT5), .B(G41), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n436), .A2(new_n275), .A3(G274), .A4(new_n431), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n435), .A2(new_n437), .A3(KEYINPUT77), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT77), .B1(new_n435), .B2(new_n437), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(G250), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G283), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G244), .B(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT4), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(G1698), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(G244), .C1(new_n291), .C2(new_n290), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n379), .A2(KEYINPUT76), .A3(G244), .A4(new_n447), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n443), .A2(new_n446), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n283), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n440), .A2(new_n453), .A3(G190), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n430), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n450), .A2(new_n451), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n441), .A2(new_n442), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n445), .B2(new_n444), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n275), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n435), .A2(new_n437), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n435), .A2(new_n437), .A3(KEYINPUT77), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(G200), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT78), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n440), .A2(new_n453), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(KEYINPUT78), .A3(G200), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n455), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(G169), .B1(new_n459), .B2(new_n464), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n440), .A2(new_n453), .A3(new_n311), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n430), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n249), .A2(G45), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n275), .A2(G250), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n275), .A2(G274), .A3(new_n431), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(G244), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n479));
  OAI211_X1 g0279(.A(G238), .B(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G116), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n283), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G200), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT19), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n224), .B1(new_n339), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G107), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n394), .A2(new_n214), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n224), .B(G68), .C1(new_n290), .C2(new_n291), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n486), .B1(new_n265), .B2(new_n214), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n256), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n254), .A2(new_n324), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n260), .A2(new_n262), .A3(G87), .A4(new_n418), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n478), .A2(new_n483), .A3(G190), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n485), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n478), .A2(new_n483), .A3(new_n310), .ZN(new_n500));
  INV_X1    g0300(.A(new_n324), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n260), .A2(new_n262), .A3(new_n501), .A4(new_n418), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n494), .A2(new_n495), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n477), .B1(new_n283), .B2(new_n482), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n500), .B(new_n503), .C1(new_n504), .C2(G169), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n470), .A2(new_n473), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n224), .B2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n488), .A2(KEYINPUT23), .A3(G20), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n266), .A2(G116), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n224), .B(G87), .C1(new_n290), .C2(new_n291), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT82), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n379), .A2(KEYINPUT82), .A3(new_n224), .A4(G87), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT83), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n513), .B2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n512), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT83), .A4(KEYINPUT22), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT84), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT24), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n262), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT22), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n522), .B(new_n511), .C1(new_n526), .C2(new_n519), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n521), .A2(KEYINPUT84), .A3(new_n522), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(KEYINPUT24), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n254), .A2(new_n488), .ZN(new_n533));
  XOR2_X1   g0333(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n534));
  OR2_X1    g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n257), .A2(new_n418), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n488), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n542));
  OAI211_X1 g0342(.A(G250), .B(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n543));
  INV_X1    g0343(.A(G294), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n543), .C1(new_n273), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n283), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n434), .A2(G264), .A3(new_n275), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n437), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT86), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(G169), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n547), .B1(new_n283), .B2(new_n545), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n552), .A2(G179), .A3(new_n437), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n550), .B1(new_n549), .B2(G169), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n541), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G200), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G190), .B2(new_n549), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n529), .A2(KEYINPUT24), .A3(new_n530), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n256), .B1(new_n529), .B2(KEYINPUT24), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n540), .B(new_n561), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n507), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(G264), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n379), .A2(KEYINPUT79), .A3(G264), .A4(G1698), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n215), .B1(new_n287), .B2(new_n288), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n286), .B1(new_n292), .B2(G303), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n570), .A2(KEYINPUT80), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT80), .B1(new_n570), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n283), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n434), .A2(G270), .A3(new_n275), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n437), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G116), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n254), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n260), .A2(new_n262), .A3(G116), .A4(new_n418), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n255), .A2(new_n223), .B1(G20), .B2(new_n580), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n442), .B(new_n224), .C1(G33), .C2(new_n214), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n584), .A2(KEYINPUT20), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT20), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(G169), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT21), .B1(new_n579), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n570), .A2(new_n572), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT80), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n570), .A2(KEYINPUT80), .A3(new_n572), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n275), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(KEYINPUT21), .B(new_n590), .C1(new_n596), .C2(new_n577), .ZN(new_n597));
  INV_X1    g0397(.A(new_n583), .ZN(new_n598));
  INV_X1    g0398(.A(new_n588), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n576), .A2(new_n437), .A3(G179), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n575), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n591), .B1(new_n604), .B2(KEYINPUT81), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n602), .B1(new_n583), .B2(new_n588), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n594), .A2(new_n595), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n283), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n589), .B1(new_n575), .B2(new_n578), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(KEYINPUT21), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n600), .B1(new_n579), .B2(G200), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n299), .B2(new_n579), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n565), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n416), .A2(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n404), .A2(new_n405), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n373), .A2(new_n331), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n369), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n414), .A2(new_n409), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n306), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n312), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n416), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n459), .A2(new_n464), .A3(new_n310), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n308), .B1(new_n440), .B2(new_n453), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT87), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n471), .A2(new_n629), .A3(new_n472), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n424), .B1(new_n422), .B2(new_n421), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n633), .A2(new_n224), .B1(new_n326), .B2(new_n362), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n380), .B1(new_n379), .B2(G20), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n488), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n256), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n417), .A3(new_n419), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n499), .A2(new_n639), .A3(new_n505), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n631), .A2(new_n632), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n626), .B2(new_n627), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT26), .B1(new_n643), .B2(new_n506), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n505), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT78), .B1(new_n468), .B2(G200), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n466), .B(new_n559), .C1(new_n440), .C2(new_n453), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n430), .B(new_n454), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n506), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n564), .A2(new_n643), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n579), .A2(new_n590), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT21), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n558), .A2(new_n610), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n645), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n624), .B1(new_n625), .B2(new_n655), .ZN(G369));
  AOI21_X1  g0456(.A(new_n556), .B1(new_n532), .B2(new_n540), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n249), .A2(new_n224), .A3(G13), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT88), .Z(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n539), .B1(new_n525), .B2(new_n531), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n564), .B1(new_n669), .B2(new_n556), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n665), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n541), .A2(new_n664), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n558), .A2(new_n673), .A3(KEYINPUT89), .A4(new_n564), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT90), .B1(new_n558), .B2(new_n665), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT90), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n657), .A2(new_n677), .A3(new_n664), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n597), .A2(new_n611), .A3(new_n603), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n611), .B1(new_n597), .B2(new_n603), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n681), .A2(new_n682), .A3(new_n591), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n664), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n667), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n664), .A2(new_n600), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n604), .B2(new_n591), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n615), .B2(new_n686), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n680), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n227), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n489), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n222), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n694), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n471), .A2(new_n629), .A3(new_n472), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n629), .B1(new_n471), .B2(new_n472), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n641), .B(KEYINPUT26), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n632), .B1(new_n643), .B2(new_n506), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(KEYINPUT93), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n631), .A2(new_n705), .A3(KEYINPUT26), .A4(new_n641), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n704), .A2(new_n505), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n558), .A2(new_n612), .A3(new_n605), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n650), .ZN(new_n709));
  AOI211_X1 g0509(.A(KEYINPUT94), .B(new_n664), .C1(new_n707), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT94), .ZN(new_n711));
  INV_X1    g0511(.A(new_n505), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n632), .B(new_n640), .C1(new_n628), .C2(new_n630), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n705), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n653), .B1(new_n610), .B2(new_n611), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n715), .A2(new_n657), .A3(new_n681), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n564), .A2(new_n643), .A3(new_n648), .A4(new_n649), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n704), .B(new_n714), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n711), .B1(new_n718), .B2(new_n665), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT29), .B1(new_n710), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT95), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n717), .B1(new_n683), .B2(new_n558), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n704), .A2(new_n505), .A3(new_n706), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n665), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT94), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n718), .A2(new_n711), .A3(new_n665), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT95), .A3(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n654), .A2(new_n650), .ZN(new_n731));
  INV_X1    g0531(.A(new_n645), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n664), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT92), .B1(new_n733), .B2(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT92), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n735), .B(new_n736), .C1(new_n655), .C2(new_n664), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n273), .A2(new_n544), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n294), .B2(G250), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n275), .B1(new_n741), .B2(new_n542), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(new_n601), .A3(new_n547), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n453), .A3(new_n440), .A4(new_n504), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n739), .B1(new_n744), .B2(new_n596), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n549), .A2(new_n310), .A3(new_n484), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n746), .B(new_n468), .C1(new_n596), .C2(new_n577), .ZN(new_n747));
  INV_X1    g0547(.A(new_n468), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n504), .A2(new_n552), .A3(new_n602), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n575), .A3(new_n749), .A4(KEYINPUT30), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n745), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n752));
  AOI21_X1  g0552(.A(KEYINPUT31), .B1(new_n751), .B2(new_n664), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT91), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n664), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT91), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n565), .A2(new_n615), .A3(new_n664), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n730), .A2(new_n738), .B1(G330), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n699), .B1(new_n764), .B2(G1), .ZN(G364));
  NAND2_X1  g0565(.A1(new_n224), .A2(G13), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n249), .B1(new_n767), .B2(G45), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n693), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n379), .A2(new_n227), .ZN(new_n771));
  INV_X1    g0571(.A(G355), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n772), .B1(G116), .B2(new_n227), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n243), .A2(new_n276), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n692), .A2(new_n379), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n222), .B2(new_n276), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n773), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n223), .B1(G20), .B2(new_n308), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n770), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G179), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n559), .ZN(new_n787));
  OAI21_X1  g0587(.A(G20), .B1(new_n787), .B2(new_n299), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n214), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n311), .A2(G20), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n299), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n292), .B(new_n790), .C1(new_n792), .C2(G50), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n224), .A2(G190), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(new_n786), .A3(new_n559), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT96), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT96), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G159), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT97), .B(KEYINPUT32), .Z(new_n801));
  OAI21_X1  g0601(.A(new_n793), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n559), .A2(G179), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT98), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n794), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G107), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n224), .A2(new_n299), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n311), .A2(new_n559), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n311), .A2(new_n559), .A3(new_n794), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G58), .A2(new_n813), .B1(new_n815), .B2(G77), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n804), .A2(new_n811), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n394), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n791), .A2(G190), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(G68), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n810), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n802), .B(new_n821), .C1(new_n800), .C2(new_n801), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n809), .A2(G283), .ZN(new_n825));
  INV_X1    g0625(.A(G329), .ZN(new_n826));
  INV_X1    g0626(.A(G322), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n798), .A2(new_n826), .B1(new_n827), .B2(new_n812), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n292), .B1(new_n789), .B2(new_n544), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G311), .B2(new_n815), .ZN(new_n832));
  INV_X1    g0632(.A(new_n817), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(G303), .B1(new_n792), .B2(G326), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n825), .A2(new_n830), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n824), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n785), .B1(new_n837), .B2(new_n782), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n781), .B(KEYINPUT101), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n688), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n689), .A2(new_n770), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(G330), .B2(new_n688), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  NAND2_X1  g0644(.A1(new_n331), .A2(new_n665), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n335), .A2(new_n333), .B1(new_n329), .B2(new_n664), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n846), .B2(new_n331), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n733), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n847), .B(KEYINPUT104), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n733), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n763), .A2(G330), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n770), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  INV_X1    g0654(.A(new_n770), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n782), .A2(new_n779), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n326), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n379), .B(new_n790), .C1(new_n833), .C2(G107), .ZN(new_n858));
  INV_X1    g0658(.A(G311), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n544), .B2(new_n812), .C1(new_n859), .C2(new_n798), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n792), .A2(G303), .B1(new_n815), .B2(G116), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  INV_X1    g0662(.A(new_n819), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT102), .Z(new_n865));
  AOI211_X1 g0665(.A(new_n860), .B(new_n865), .C1(G87), .C2(new_n809), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT103), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n792), .A2(G137), .B1(new_n813), .B2(G143), .ZN(new_n868));
  INV_X1    g0668(.A(G150), .ZN(new_n869));
  INV_X1    g0669(.A(G159), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n868), .B1(new_n869), .B2(new_n863), .C1(new_n870), .C2(new_n814), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT34), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n808), .A2(new_n202), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n379), .B1(new_n201), .B2(new_n789), .C1(new_n817), .C2(new_n207), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(G132), .B2(new_n799), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n867), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(KEYINPUT103), .B2(new_n866), .ZN(new_n881));
  INV_X1    g0681(.A(new_n782), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n857), .B1(new_n780), .B2(new_n848), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n854), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G384));
  OR2_X1    g0685(.A1(new_n426), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n426), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n225), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n889));
  XNOR2_X1  g0689(.A(new_n888), .B(new_n889), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n222), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n207), .A2(G68), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n249), .B(G13), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n625), .B1(new_n734), .B2(new_n737), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n623), .B1(new_n730), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n411), .A2(new_n413), .ZN(new_n898));
  INV_X1    g0698(.A(new_n662), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n411), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n900), .A3(new_n401), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT37), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n898), .A2(new_n900), .A3(new_n903), .A4(new_n401), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n900), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n415), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n905), .A2(new_n907), .A3(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT106), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n897), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n369), .A2(new_n664), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n910), .A2(KEYINPUT106), .A3(KEYINPUT39), .A4(new_n911), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n849), .A2(new_n845), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n664), .A2(new_n368), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n369), .A2(new_n373), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n373), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n368), .B(new_n664), .C1(new_n359), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n918), .A2(new_n912), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n621), .A2(new_n662), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n917), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n896), .B(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n752), .A2(new_n753), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n762), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n847), .B1(new_n920), .B2(new_n922), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n912), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n930), .A2(new_n912), .A3(KEYINPUT40), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n416), .A2(new_n930), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(G330), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n927), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n249), .B2(new_n767), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n927), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n894), .B1(new_n942), .B2(new_n943), .ZN(G367));
  NOR2_X1   g0744(.A1(new_n665), .A2(new_n497), .ZN(new_n945));
  MUX2_X1   g0745(.A(new_n649), .B(new_n712), .S(new_n945), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n665), .A2(new_n430), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n631), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n648), .A2(new_n643), .ZN(new_n950));
  OAI22_X1  g0750(.A1(KEYINPUT107), .A2(new_n949), .B1(new_n950), .B2(new_n948), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n949), .A2(KEYINPUT107), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n643), .B1(new_n953), .B2(new_n558), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n665), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n672), .A2(new_n674), .B1(new_n676), .B2(new_n678), .ZN(new_n957));
  INV_X1    g0757(.A(new_n684), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n957), .A2(new_n958), .A3(new_n953), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT42), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n955), .B(new_n956), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n680), .A2(new_n684), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT42), .B1(new_n964), .B2(new_n953), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n956), .B1(new_n965), .B2(new_n955), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n947), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n953), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n689), .A2(new_n680), .A3(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT109), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n958), .B1(new_n675), .B2(new_n679), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n960), .B1(new_n974), .B2(new_n968), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n954), .A2(new_n665), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT108), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(new_n962), .A3(new_n961), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n947), .A3(new_n970), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n972), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n973), .ZN(new_n981));
  AND3_X1   g0781(.A1(new_n978), .A2(new_n947), .A3(new_n970), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n970), .B1(new_n978), .B2(new_n947), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n693), .B(new_n985), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n688), .A2(G330), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(KEYINPUT112), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n957), .A2(new_n958), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n988), .B1(new_n964), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n964), .A2(new_n989), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n987), .B(KEYINPUT112), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n685), .B2(new_n968), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n953), .B1(KEYINPUT111), .B2(KEYINPUT44), .C1(new_n974), .C2(new_n667), .ZN(new_n996));
  NAND2_X1  g0796(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n690), .A2(KEYINPUT113), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n666), .A4(new_n968), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n666), .B(new_n968), .C1(new_n957), .C2(new_n958), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n690), .A2(KEYINPUT113), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n998), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(new_n998), .B2(new_n1004), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n764), .B(new_n993), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n986), .B1(new_n1008), .B2(new_n764), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n980), .B(new_n984), .C1(new_n1009), .C2(new_n769), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n207), .A2(new_n814), .B1(new_n812), .B2(new_n869), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n379), .B1(new_n202), .B2(new_n789), .C1(new_n863), .C2(new_n870), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G143), .C2(new_n792), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n799), .A2(G137), .B1(new_n833), .B2(G58), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT114), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n809), .A2(G77), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(KEYINPUT114), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n792), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n859), .B1(new_n862), .B2(new_n814), .ZN(new_n1020));
  INV_X1    g0820(.A(G303), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n863), .A2(new_n544), .B1(new_n1021), .B2(new_n812), .ZN(new_n1022));
  INV_X1    g0822(.A(G317), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n292), .B1(new_n488), .B2(new_n789), .C1(new_n798), .C2(new_n1023), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n809), .A2(G97), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n833), .A2(G116), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT46), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1018), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT47), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n782), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n946), .A2(new_n839), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n784), .B1(new_n692), .B2(new_n501), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n238), .A2(new_n775), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n855), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1010), .A2(new_n1037), .ZN(G387));
  AOI21_X1  g0838(.A(KEYINPUT95), .B1(new_n728), .B2(KEYINPUT29), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n721), .B(new_n736), .C1(new_n726), .C2(new_n727), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n738), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n852), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n993), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n852), .A3(new_n993), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n693), .A3(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n680), .A2(new_n839), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n771), .A2(new_n695), .B1(G107), .B2(new_n227), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n235), .A2(new_n276), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n695), .ZN(new_n1050));
  AOI211_X1 g0850(.A(G45), .B(new_n1050), .C1(G68), .C2(G77), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n321), .A2(G50), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n776), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1048), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n770), .B1(new_n1055), .B2(new_n784), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n207), .A2(new_n812), .B1(new_n814), .B2(new_n202), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n379), .B1(new_n324), .B2(new_n789), .C1(new_n1019), .C2(new_n870), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n264), .C2(new_n819), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n817), .A2(new_n326), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n799), .B2(G150), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT115), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT115), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1059), .A2(new_n1026), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n817), .A2(new_n544), .B1(new_n862), .B2(new_n789), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n819), .A2(G311), .B1(new_n815), .B2(G303), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n1023), .B2(new_n812), .C1(new_n827), .C2(new_n1019), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n379), .B1(new_n799), .B2(G326), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n808), .B2(new_n580), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT116), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1064), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1056), .B1(new_n1077), .B2(new_n782), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n993), .A2(new_n769), .B1(new_n1047), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1046), .A2(new_n1079), .ZN(G393));
  INV_X1    g0880(.A(new_n1007), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n998), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n1045), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1008), .A2(new_n1083), .A3(new_n693), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n769), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n953), .A2(new_n781), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n247), .A2(new_n776), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n783), .B1(new_n214), .B2(new_n227), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n770), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n863), .A2(new_n207), .B1(new_n202), .B2(new_n817), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n322), .B2(new_n815), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n379), .B1(new_n789), .B2(new_n326), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n799), .B2(G143), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(new_n394), .C2(new_n808), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n792), .A2(G150), .B1(new_n813), .B2(G159), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n863), .A2(new_n1021), .B1(new_n862), .B2(new_n817), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G322), .B2(new_n799), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n292), .B1(new_n789), .B2(new_n580), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G294), .B2(new_n815), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n810), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n792), .A2(G317), .B1(new_n813), .B2(G311), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT52), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1095), .A2(new_n1097), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1090), .B1(new_n1105), .B2(new_n782), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1087), .A2(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1085), .A2(new_n1086), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1086), .B1(new_n1085), .B2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1084), .B1(new_n1108), .B2(new_n1109), .ZN(G390));
  OAI211_X1 g0910(.A(G330), .B(new_n848), .C1(new_n761), .C2(new_n762), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT119), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n923), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n930), .A2(G330), .A3(new_n931), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1112), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n918), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1111), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT118), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n923), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n920), .A2(KEYINPUT118), .A3(new_n922), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n850), .B(G330), .C1(new_n762), .C2(new_n929), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n923), .A2(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n726), .A2(new_n727), .A3(new_n845), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n846), .A2(new_n331), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1118), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n930), .A2(G330), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n416), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n896), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1122), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT118), .B1(new_n920), .B2(new_n922), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1126), .A2(new_n1127), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n915), .B1(new_n910), .B2(new_n911), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n914), .A2(new_n916), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n733), .A2(new_n1127), .B1(new_n331), .B2(new_n665), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1141), .A2(new_n1113), .B1(new_n369), .B2(new_n664), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1119), .A2(new_n923), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1139), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1137), .A2(new_n1138), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n1115), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n694), .B1(new_n1133), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n895), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n624), .A3(new_n1132), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n931), .A3(new_n1131), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n1153), .A3(new_n1145), .A4(new_n1130), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1140), .A2(new_n779), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n855), .B1(new_n376), .B2(new_n856), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1019), .A2(new_n862), .B1(new_n544), .B2(new_n798), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n379), .B(new_n818), .C1(G77), .C2(new_n788), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n488), .B2(new_n863), .C1(new_n580), .C2(new_n812), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(G97), .C2(new_n815), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n379), .B1(new_n789), .B2(new_n870), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n799), .A2(G125), .B1(new_n792), .B2(G128), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT54), .B(G143), .Z(new_n1164));
  AOI22_X1  g0964(.A1(new_n813), .A2(G132), .B1(new_n815), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1162), .B(new_n1166), .C1(G137), .C2(new_n819), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT53), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n817), .B2(new_n869), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n833), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n809), .A2(G50), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1161), .A2(new_n876), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1156), .B(new_n1157), .C1(new_n882), .C2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1147), .B2(new_n768), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1155), .A2(new_n1174), .ZN(G378));
  INV_X1    g0975(.A(KEYINPUT120), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1150), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n896), .A2(KEYINPUT120), .A3(new_n1132), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n1133), .C2(new_n1147), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n934), .A2(G330), .A3(new_n935), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n307), .A2(new_n662), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n306), .B2(new_n312), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n306), .A2(new_n312), .A3(new_n1183), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1181), .A2(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1192), .A2(new_n934), .A3(G330), .A4(new_n935), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n926), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1191), .A2(new_n1193), .A3(new_n926), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1180), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n694), .B1(new_n1179), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT121), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1191), .A2(new_n1193), .A3(new_n926), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n926), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT120), .B1(new_n896), .B2(new_n1132), .ZN(new_n1204));
  AND4_X1   g1004(.A1(KEYINPUT120), .A2(new_n1149), .A3(new_n624), .A4(new_n1132), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1203), .B1(new_n1206), .B2(new_n1154), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1199), .A2(new_n1200), .B1(new_n1207), .B2(KEYINPUT57), .ZN(new_n1208));
  AOI211_X1 g1008(.A(KEYINPUT121), .B(new_n694), .C1(new_n1179), .C2(new_n1198), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1203), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1190), .A2(new_n779), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n863), .A2(new_n214), .B1(new_n862), .B2(new_n798), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G107), .B2(new_n813), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n809), .A2(G58), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n292), .A2(new_n274), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1216), .B(new_n1060), .C1(G68), .C2(new_n788), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n792), .A2(G116), .B1(new_n815), .B2(new_n501), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1216), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n833), .A2(new_n1164), .B1(new_n792), .B2(G125), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G128), .A2(new_n813), .B1(new_n815), .B2(G137), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n819), .A2(G132), .B1(G150), .B2(new_n788), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n809), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1223), .B1(new_n1220), .B2(new_n1219), .C1(new_n1228), .C2(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1233), .A2(new_n782), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n855), .B(new_n1234), .C1(new_n207), .C2(new_n856), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n1211), .A2(new_n769), .B1(new_n1212), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1210), .A2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT119), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(new_n1115), .A3(new_n1114), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1240), .A2(new_n918), .B1(new_n1128), .B2(new_n1125), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1150), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n986), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1133), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n855), .B1(new_n202), .B2(new_n856), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n799), .A2(G303), .B1(G107), .B2(new_n815), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n214), .B2(new_n817), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n292), .B1(new_n324), .B2(new_n789), .C1(new_n863), .C2(new_n580), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n1019), .A2(new_n544), .B1(new_n862), .B2(new_n812), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n799), .A2(G128), .B1(new_n819), .B2(new_n1164), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n870), .B2(new_n817), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n792), .A2(G132), .B1(new_n813), .B2(G137), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n292), .B1(new_n788), .B2(G50), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n869), .C2(new_n814), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1250), .A2(new_n1016), .B1(new_n1256), .B2(new_n1215), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1245), .B1(new_n882), .B2(new_n1257), .C1(new_n1136), .C2(new_n780), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1130), .B2(new_n769), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1244), .A2(new_n1260), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1261), .B(KEYINPUT122), .ZN(G381));
  NOR2_X1   g1062(.A1(new_n1155), .A2(new_n1174), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n768), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1107), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT117), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1085), .A2(new_n1086), .A3(new_n1107), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1045), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n694), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1266), .A2(new_n1267), .B1(new_n1270), .B2(new_n1083), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1263), .A2(new_n884), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G387), .A2(G375), .A3(G381), .A4(new_n1273), .ZN(G407));
  AND2_X1   g1074(.A1(new_n1210), .A2(new_n1236), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1275), .A2(G213), .A3(new_n663), .A4(new_n1263), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G407), .A2(G213), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT123), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(G407), .A2(new_n1279), .A3(G213), .A4(new_n1276), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(G409));
  NAND2_X1  g1081(.A1(new_n984), .A2(new_n980), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1045), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1243), .B1(new_n1283), .B2(new_n1042), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1284), .B2(new_n768), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1037), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1271), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1010), .A2(G390), .A3(new_n1037), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n843), .B1(new_n1046), .B2(new_n1079), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1272), .A2(new_n1289), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G378), .B(new_n1236), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1207), .A2(new_n1243), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1236), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1263), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n663), .A2(G213), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT124), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT60), .B1(new_n1150), .B2(new_n1241), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1242), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n1241), .ZN(new_n1305));
  AND4_X1   g1105(.A1(new_n1302), .A2(new_n1304), .A3(new_n693), .A4(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n694), .B1(new_n1303), .B2(new_n1242), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1302), .B1(new_n1307), .B2(new_n1305), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1260), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n884), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1304), .A2(new_n693), .A3(new_n1305), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(KEYINPUT124), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1307), .A2(new_n1302), .A3(new_n1305), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(G384), .A3(new_n1260), .ZN(new_n1315));
  INV_X1    g1115(.A(G2897), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1300), .A2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1310), .A2(new_n1315), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1310), .B2(new_n1315), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1301), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1295), .A2(new_n1298), .B1(G213), .B2(new_n663), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1310), .A2(new_n1315), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT127), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1320), .B(new_n1321), .C1(new_n1325), .C2(KEYINPUT62), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1294), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT125), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1329));
  AOI21_X1  g1129(.A(G384), .B1(new_n1314), .B2(new_n1260), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1260), .ZN(new_n1331));
  AOI211_X1 g1131(.A(new_n884), .B(new_n1331), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1332));
  OAI22_X1  g1132(.A1(new_n1330), .A2(new_n1332), .B1(new_n1316), .B2(new_n1300), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1310), .A2(new_n1315), .A3(new_n1317), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1329), .A2(new_n1336), .A3(new_n1301), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT63), .B1(new_n1322), .B2(new_n1324), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1292), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1321), .A3(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1310), .A2(new_n1315), .A3(KEYINPUT63), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1342), .B1(new_n1322), .B2(new_n1344), .ZN(new_n1345));
  AND4_X1   g1145(.A1(KEYINPUT126), .A2(new_n1337), .A3(new_n1339), .A4(new_n1345), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1291), .A2(new_n1292), .A3(KEYINPUT61), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1347), .B1(new_n1301), .B2(new_n1343), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1348), .A2(new_n1338), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT126), .B1(new_n1349), .B2(new_n1337), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1328), .B1(new_n1346), .B2(new_n1350), .ZN(G405));
  NAND2_X1  g1151(.A1(G375), .A2(new_n1263), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1295), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1324), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1352), .A2(new_n1323), .A3(new_n1295), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1294), .ZN(G402));
endmodule


