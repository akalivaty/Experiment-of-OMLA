//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n202), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G97), .C2(G257), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G1), .B2(G20), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n207), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  AOI211_X1 g0026(.A(new_n210), .B(new_n222), .C1(new_n224), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT65), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  OAI211_X1 g0045(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G232), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT78), .ZN(new_n253));
  INV_X1    g0053(.A(G179), .ZN(new_n254));
  OR2_X1    g0054(.A1(G223), .A2(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n216), .A2(G1698), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n255), .B(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G87), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n248), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT78), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(new_n246), .C1(new_n250), .C2(new_n251), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n253), .A2(new_n254), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G169), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n248), .B1(new_n259), .B2(new_n260), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n252), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n272), .A2(new_n223), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n257), .A2(new_n258), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT7), .B1(new_n274), .B2(new_n207), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT7), .ZN(new_n276));
  NOR4_X1   g0076(.A1(new_n257), .A2(new_n258), .A3(new_n276), .A4(G20), .ZN(new_n277));
  OAI21_X1  g0077(.A(G68), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G58), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(new_n217), .ZN(new_n280));
  OAI21_X1  g0080(.A(G20), .B1(new_n280), .B2(new_n201), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G159), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT16), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n273), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n257), .A2(new_n258), .A3(G20), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT75), .B1(new_n289), .B2(KEYINPUT7), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  INV_X1    g0091(.A(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n207), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT75), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(new_n276), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n277), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT16), .B(new_n285), .C1(new_n298), .C2(new_n217), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT76), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n288), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n288), .B2(new_n299), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT8), .B(G58), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n272), .A2(new_n223), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n206), .B2(G20), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n308), .B1(new_n311), .B2(new_n305), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT77), .B1(new_n303), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n295), .A2(new_n296), .A3(new_n276), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n296), .B1(new_n295), .B2(new_n276), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI211_X1 g0118(.A(new_n287), .B(new_n284), .C1(new_n318), .C2(G68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n295), .A2(new_n276), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n217), .B1(new_n320), .B2(new_n315), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n287), .B1(new_n321), .B2(new_n284), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n309), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT76), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n288), .A2(new_n299), .A3(new_n300), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT77), .A4(new_n313), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n271), .B1(new_n314), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT18), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT17), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n253), .A2(new_n331), .A3(new_n263), .A4(new_n265), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n268), .B2(new_n252), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT79), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(KEYINPUT79), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n339), .A2(new_n324), .A3(new_n313), .A4(new_n325), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n330), .B1(new_n340), .B2(KEYINPUT80), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n301), .A2(new_n302), .A3(new_n312), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT80), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT17), .A4(new_n339), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n324), .A2(new_n313), .A3(new_n325), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n326), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n271), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n329), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n293), .A2(new_n294), .ZN(new_n354));
  INV_X1    g0154(.A(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G222), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT67), .B(G223), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n354), .B(new_n356), .C1(new_n357), .C2(new_n355), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n262), .C1(G77), .C2(new_n354), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n246), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n248), .A2(new_n249), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G226), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n267), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n203), .A2(G20), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  INV_X1    g0166(.A(new_n282), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n207), .A2(G33), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n365), .B1(new_n366), .B2(new_n367), .C1(new_n304), .C2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n309), .B1(new_n202), .B2(new_n307), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n202), .B2(new_n311), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT68), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n363), .A2(G179), .ZN(new_n374));
  XOR2_X1   g0174(.A(new_n374), .B(KEYINPUT69), .Z(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n360), .A2(G190), .A3(new_n362), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT72), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n363), .A2(G200), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n371), .B(KEYINPUT9), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n379), .A2(KEYINPUT10), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT10), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G77), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n367), .A2(new_n202), .B1(new_n368), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n207), .A2(G68), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n309), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n389), .A2(new_n390), .B1(new_n311), .B2(new_n217), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n206), .A3(G13), .ZN(new_n393));
  XOR2_X1   g0193(.A(new_n393), .B(KEYINPUT12), .Z(new_n394));
  OR3_X1    g0194(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  INV_X1    g0196(.A(new_n246), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n216), .A2(new_n355), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n398), .B1(G232), .B2(new_n355), .C1(new_n257), .C2(new_n258), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G97), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n401), .B2(new_n262), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n361), .A2(G238), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n400), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n293), .A2(new_n294), .B1(new_n251), .B2(G1698), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n246), .B(new_n403), .C1(new_n407), .C2(new_n248), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n395), .B1(new_n410), .B2(G190), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n333), .B2(new_n410), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n376), .A2(new_n382), .A3(new_n385), .A4(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(KEYINPUT73), .B(G169), .C1(new_n404), .C2(new_n409), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT14), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n402), .A2(new_n396), .A3(new_n403), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n408), .A2(KEYINPUT13), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(KEYINPUT73), .A3(new_n419), .A4(G169), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT74), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n410), .A2(new_n421), .A3(G179), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT74), .B1(new_n418), .B2(new_n254), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n415), .A2(new_n420), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n424), .A2(new_n395), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n304), .B(KEYINPUT71), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT15), .B(G87), .Z(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n426), .A2(new_n367), .B1(new_n368), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n207), .A2(new_n386), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n309), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n307), .A2(new_n386), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n310), .A2(G77), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G238), .A2(G1698), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n354), .B(new_n436), .C1(new_n251), .C2(G1698), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT70), .B(G107), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n262), .C1(new_n354), .C2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G244), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n246), .C1(new_n440), .C2(new_n250), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G200), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n435), .B(new_n442), .C1(new_n331), .C2(new_n441), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n267), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n434), .B(new_n444), .C1(G179), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n425), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n353), .A2(new_n413), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n354), .B2(G250), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n355), .ZN(new_n453));
  OAI21_X1  g0253(.A(G244), .B1(new_n257), .B2(new_n258), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n451), .A2(G1698), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(G244), .C1(new_n258), .C2(new_n257), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n262), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n462), .B(G274), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n462), .B1(new_n464), .B2(new_n463), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n466), .A2(new_n248), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G257), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n460), .A2(G190), .A3(new_n465), .A4(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n460), .A2(new_n465), .A3(new_n468), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(new_n333), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n306), .A2(G97), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n438), .B1(new_n275), .B2(new_n277), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT81), .B1(new_n282), .B2(G77), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT6), .ZN(new_n475));
  AND2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G97), .A2(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G107), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(KEYINPUT6), .A3(G97), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n474), .B1(new_n481), .B2(G20), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n282), .A2(KEYINPUT81), .A3(G77), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n473), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n472), .B1(new_n484), .B2(new_n309), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n206), .A2(G33), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n273), .A2(new_n306), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G97), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT82), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n471), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n454), .A2(new_n451), .B1(G33), .B2(G283), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n458), .C1(new_n355), .C2(new_n452), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(new_n262), .B1(G257), .B2(new_n467), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n267), .B1(new_n497), .B2(new_n465), .ZN(new_n498));
  AND4_X1   g0298(.A1(G179), .A2(new_n460), .A3(new_n465), .A4(new_n468), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n207), .B(G68), .C1(new_n257), .C2(new_n258), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n502), .A2(new_n503), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  INV_X1    g0306(.A(G87), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n507), .B(new_n508), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n400), .A2(new_n207), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n400), .A2(KEYINPUT19), .A3(G20), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n504), .B(new_n505), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n309), .B1(new_n307), .B2(new_n428), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n462), .A2(G274), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n248), .B(G250), .C1(G1), .C2(new_n461), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n293), .A2(new_n294), .B1(new_n440), .B2(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n218), .A2(new_n355), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n519), .A2(new_n520), .B1(G33), .B2(G116), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n517), .B(new_n518), .C1(new_n521), .C2(new_n248), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G190), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(G200), .ZN(new_n525));
  OR3_X1    g0325(.A1(new_n487), .A2(KEYINPUT84), .A3(new_n507), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT84), .B1(new_n487), .B2(new_n507), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n516), .A2(new_n524), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n505), .A2(new_n504), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n507), .A2(new_n508), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n512), .B1(new_n438), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n514), .B1(new_n532), .B2(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n309), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n428), .A2(new_n307), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n488), .A2(new_n427), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n522), .A2(new_n267), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n523), .A2(new_n254), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n529), .A2(new_n540), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n494), .A2(new_n501), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n354), .B1(G257), .B2(new_n355), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G250), .A2(G1698), .ZN(new_n544));
  INV_X1    g0344(.A(G294), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n543), .A2(new_n544), .B1(new_n292), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(new_n262), .B1(G264), .B2(new_n467), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n267), .B1(new_n547), .B2(new_n465), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n465), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n550), .B2(G179), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT90), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n487), .A2(new_n479), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n207), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT87), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT22), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(KEYINPUT22), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n354), .A2(new_n207), .A3(G87), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT88), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n565));
  OR2_X1    g0365(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n565), .B(new_n566), .C1(new_n438), .C2(new_n207), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n560), .A2(new_n562), .A3(new_n564), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n567), .A2(new_n564), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n562), .A4(new_n560), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n554), .B1(new_n573), .B2(new_n309), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n307), .A2(new_n479), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT25), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n553), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n273), .B1(new_n569), .B2(new_n572), .ZN(new_n579));
  NOR4_X1   g0379(.A1(new_n579), .A2(KEYINPUT90), .A3(new_n554), .A4(new_n576), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n552), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT85), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n487), .B2(new_n212), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n307), .A2(new_n309), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(KEYINPUT85), .A3(G116), .A4(new_n486), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n456), .B(new_n207), .C1(G33), .C2(new_n508), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n212), .A2(G20), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n309), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n306), .A2(G116), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT86), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n586), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n355), .A2(G257), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n354), .B(new_n595), .C1(new_n229), .C2(new_n355), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n262), .C1(G303), .C2(new_n354), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n467), .A2(G270), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n465), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(G169), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT21), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n594), .A2(new_n602), .A3(G169), .A4(new_n599), .ZN(new_n603));
  INV_X1    g0403(.A(new_n594), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n599), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n601), .A2(new_n603), .B1(new_n605), .B2(G179), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n599), .A2(G200), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n604), .B(new_n607), .C1(new_n331), .C2(new_n599), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n550), .A2(G190), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n549), .A2(G200), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n574), .A2(new_n577), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n542), .A2(new_n581), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n450), .A2(new_n613), .ZN(G372));
  AND3_X1   g0414(.A1(new_n347), .A2(KEYINPUT18), .A3(new_n271), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT18), .B1(new_n347), .B2(new_n271), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT93), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n445), .B(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n425), .B1(new_n412), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n620), .B2(new_n345), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n385), .A2(new_n382), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n623), .A2(new_n376), .ZN(new_n624));
  INV_X1    g0424(.A(new_n471), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n485), .A2(new_n492), .A3(new_n489), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n492), .B1(new_n485), .B2(new_n489), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT91), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n534), .A2(new_n528), .A3(new_n535), .ZN(new_n630));
  INV_X1    g0430(.A(new_n525), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n516), .A2(KEYINPUT91), .A3(new_n525), .A4(new_n528), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n524), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n628), .A2(new_n612), .A3(new_n500), .A4(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n579), .A2(new_n554), .A3(new_n576), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n551), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n601), .A2(new_n603), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n605), .A2(G179), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n626), .A2(new_n627), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n497), .A2(new_n465), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G169), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n470), .A2(G179), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n634), .A2(new_n643), .A3(new_n540), .A4(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n541), .A2(new_n500), .ZN(new_n650));
  XNOR2_X1  g0450(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n540), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n642), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n624), .B1(new_n450), .B2(new_n654), .ZN(G369));
  INV_X1    g0455(.A(G13), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G20), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n206), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n594), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n609), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n606), .B2(new_n664), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n578), .A2(new_n580), .ZN(new_n668));
  INV_X1    g0468(.A(new_n663), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n581), .B(new_n612), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n581), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n606), .A2(new_n663), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT94), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n671), .A2(new_n674), .B1(new_n637), .B2(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n208), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n511), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n225), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n683));
  XNOR2_X1  g0483(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n635), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n581), .A2(new_n606), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n650), .A2(new_n651), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n634), .A2(new_n643), .A3(KEYINPUT26), .A4(new_n647), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n663), .B1(new_n689), .B2(new_n540), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n648), .A2(new_n649), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n650), .A2(new_n651), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n494), .A2(new_n501), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n606), .B1(new_n636), .B2(new_n551), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n612), .A4(new_n634), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n696), .A3(new_n540), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n669), .ZN(new_n698));
  XNOR2_X1  g0498(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n690), .A2(KEYINPUT29), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n550), .A2(G179), .A3(new_n523), .ZN(new_n702));
  INV_X1    g0502(.A(new_n599), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n497), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n549), .A2(new_n254), .A3(new_n522), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n703), .A4(new_n497), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n703), .A2(G179), .A3(new_n523), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n549), .A3(new_n644), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n663), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n713), .B(new_n714), .C1(new_n613), .C2(new_n663), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n700), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n684), .B1(new_n718), .B2(G1), .ZN(G364));
  NAND2_X1  g0519(.A1(new_n657), .A2(G45), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n679), .A2(G1), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT97), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n667), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n666), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n677), .A2(new_n354), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n226), .B2(new_n461), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n244), .B2(new_n461), .ZN(new_n728));
  INV_X1    g0528(.A(G355), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n354), .A2(new_n208), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n728), .B1(G116), .B2(new_n208), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n223), .B1(G20), .B2(new_n267), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n722), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n254), .A2(G200), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT99), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n207), .A2(new_n331), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n207), .A2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n507), .A2(new_n744), .B1(new_n748), .B2(new_n479), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n207), .B1(new_n750), .B2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n749), .B1(G97), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n254), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n741), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n254), .A2(new_n333), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n745), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G58), .A2(new_n756), .B1(new_n759), .B2(G68), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n741), .A2(new_n757), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n202), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n745), .A2(new_n754), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(G77), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n745), .A2(new_n750), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT98), .B(KEYINPUT32), .Z(new_n769));
  XNOR2_X1  g0569(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n753), .A2(new_n354), .A3(new_n765), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n354), .B1(new_n743), .B2(G303), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT100), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT100), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n747), .A2(G283), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  INV_X1    g0576(.A(G329), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n763), .A2(new_n776), .B1(new_n766), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT33), .B(G317), .Z(new_n779));
  OAI22_X1  g0579(.A1(new_n779), .A2(new_n758), .B1(new_n751), .B2(new_n545), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(G322), .C2(new_n756), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n773), .A2(new_n774), .A3(new_n775), .A4(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n761), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(G326), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n771), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n738), .B1(new_n785), .B2(new_n735), .ZN(new_n786));
  INV_X1    g0586(.A(new_n734), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n737), .B(new_n786), .C1(new_n666), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n724), .A2(new_n788), .ZN(G396));
  INV_X1    g0589(.A(new_n698), .ZN(new_n790));
  INV_X1    g0590(.A(new_n446), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n435), .A2(new_n669), .ZN(new_n792));
  MUX2_X1   g0592(.A(new_n791), .B(new_n619), .S(new_n792), .Z(new_n793));
  OR2_X1    g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n697), .A2(new_n793), .A3(new_n669), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n716), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(new_n717), .A3(new_n795), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n738), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n735), .A2(new_n732), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n386), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G143), .A2(new_n756), .B1(new_n759), .B2(G150), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n803), .B2(new_n761), .C1(new_n767), .C2(new_n763), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT34), .Z(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n354), .B1(new_n806), .B2(new_n766), .C1(new_n744), .C2(new_n202), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n748), .A2(new_n217), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n751), .A2(new_n279), .ZN(new_n809));
  OR3_X1    g0609(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G303), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n761), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n758), .A2(new_n813), .B1(new_n763), .B2(new_n212), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT101), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n747), .A2(G87), .B1(new_n743), .B2(G107), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n274), .B1(new_n766), .B2(new_n776), .C1(new_n545), .C2(new_n755), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G97), .B2(new_n752), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n805), .A2(new_n810), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n738), .B1(new_n820), .B2(new_n735), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n801), .B(new_n821), .C1(new_n793), .C2(new_n733), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n799), .A2(new_n822), .ZN(G384));
  INV_X1    g0623(.A(G330), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n711), .A2(KEYINPUT105), .A3(new_n712), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n712), .A2(KEYINPUT105), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n710), .A2(new_n663), .A3(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(new_n613), .C2(new_n663), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n395), .A2(new_n663), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n424), .A2(new_n830), .A3(new_n395), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n424), .B2(new_n395), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n412), .B(new_n829), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n425), .A2(new_n663), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n828), .A2(new_n835), .A3(new_n793), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n285), .B1(new_n298), .B2(new_n217), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n839), .A2(KEYINPUT104), .A3(new_n287), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n287), .A2(KEYINPUT104), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n285), .B(new_n841), .C1(new_n298), .C2(new_n217), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n840), .A2(new_n309), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n313), .ZN(new_n844));
  INV_X1    g0644(.A(new_n661), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n271), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n838), .B1(new_n846), .B2(new_n340), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n314), .A2(new_n327), .B1(new_n271), .B2(new_n845), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n340), .A2(new_n838), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n844), .A2(new_n845), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n837), .B(new_n851), .C1(new_n353), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n661), .B1(new_n349), .B2(new_n326), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n340), .B1(new_n342), .B2(new_n270), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n349), .A2(new_n326), .B1(new_n270), .B2(new_n661), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n849), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n341), .B(new_n344), .C1(new_n615), .C2(new_n616), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n855), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT38), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT40), .B(new_n836), .C1(new_n854), .C2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n828), .A2(new_n835), .A3(new_n793), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n351), .B1(new_n350), .B2(new_n271), .ZN(new_n865));
  AOI211_X1 g0665(.A(KEYINPUT18), .B(new_n270), .C1(new_n349), .C2(new_n326), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n852), .B1(new_n867), .B2(new_n346), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n837), .B1(new_n868), .B2(new_n851), .ZN(new_n869));
  INV_X1    g0669(.A(new_n851), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n865), .A2(new_n866), .A3(new_n345), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT38), .B(new_n870), .C1(new_n871), .C2(new_n852), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n864), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n863), .B1(new_n873), .B2(KEYINPUT40), .ZN(new_n874));
  INV_X1    g0674(.A(new_n413), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n828), .A2(new_n871), .A3(new_n875), .A4(new_n447), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n824), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT106), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n876), .B2(new_n874), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n854), .B2(new_n862), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n831), .A2(new_n832), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n669), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n880), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n835), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n445), .A2(new_n663), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n795), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n353), .A2(new_n853), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n891), .B2(new_n870), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n892), .B2(new_n854), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n617), .A2(new_n845), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n623), .A2(new_n376), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n700), .B2(new_n449), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n879), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n206), .B2(new_n657), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n481), .B(KEYINPUT102), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n212), .B1(new_n902), .B2(KEYINPUT35), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(new_n224), .C1(KEYINPUT35), .C2(new_n902), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT36), .ZN(new_n905));
  OAI21_X1  g0705(.A(G77), .B1(new_n279), .B2(new_n217), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n906), .A2(new_n225), .B1(G50), .B2(new_n217), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G1), .A3(new_n656), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n901), .A2(new_n905), .A3(new_n908), .ZN(G367));
  INV_X1    g0709(.A(new_n672), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n643), .A2(new_n663), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n694), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n643), .A2(new_n647), .A3(new_n663), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n671), .A2(new_n674), .A3(new_n914), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n581), .B1(new_n912), .B2(new_n913), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n669), .B1(new_n918), .B2(new_n501), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n630), .A2(new_n663), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n634), .A2(new_n540), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n540), .B2(new_n921), .ZN(new_n923));
  XOR2_X1   g0723(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n917), .A2(new_n919), .A3(new_n920), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT108), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(KEYINPUT43), .B2(new_n923), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(KEYINPUT109), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT109), .B1(new_n927), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n915), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n933), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n935), .A2(new_n910), .A3(new_n914), .A4(new_n931), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n678), .B(KEYINPUT41), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n675), .A2(new_n914), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT45), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT44), .B1(new_n675), .B2(new_n914), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n675), .A2(KEYINPUT44), .A3(new_n914), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n910), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n667), .B(new_n671), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n674), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n946), .A2(new_n718), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n940), .A2(new_n672), .A3(new_n941), .A4(new_n942), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n938), .B1(new_n949), .B2(new_n718), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n720), .A2(G1), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n934), .B(new_n936), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n736), .B1(new_n208), .B2(new_n428), .C1(new_n232), .C2(new_n726), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT110), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n738), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G294), .A2(new_n759), .B1(new_n756), .B2(G303), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n813), .B2(new_n763), .C1(new_n776), .C2(new_n761), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n354), .B(new_n957), .C1(new_n438), .C2(new_n752), .ZN(new_n958));
  INV_X1    g0758(.A(new_n766), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(G317), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n743), .A2(G116), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT46), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n747), .A2(G97), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n958), .A2(new_n960), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n748), .A2(new_n386), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n279), .B2(new_n744), .C1(new_n217), .C2(new_n751), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G150), .A2(new_n756), .B1(new_n959), .B2(G137), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n202), .B2(new_n763), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G159), .B2(new_n759), .ZN(new_n970));
  INV_X1    g0770(.A(G143), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n970), .B(new_n354), .C1(new_n971), .C2(new_n761), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n964), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT47), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n735), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n955), .B1(new_n787), .B2(new_n923), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT111), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n952), .A2(new_n979), .ZN(G387));
  NOR2_X1   g0780(.A1(new_n671), .A2(new_n787), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n755), .A2(new_n982), .B1(new_n763), .B2(new_n811), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n983), .A2(KEYINPUT113), .B1(G311), .B2(new_n759), .ZN(new_n984));
  INV_X1    g0784(.A(G322), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(KEYINPUT113), .B2(new_n983), .C1(new_n985), .C2(new_n761), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT48), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n813), .B2(new_n751), .C1(new_n545), .C2(new_n744), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT49), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n959), .A2(G326), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n354), .B1(new_n747), .B2(G116), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n963), .B1(new_n428), .B2(new_n751), .C1(new_n744), .C2(new_n386), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G68), .A2(new_n764), .B1(new_n959), .B2(G150), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n202), .B2(new_n755), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G159), .B2(new_n783), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n354), .C1(new_n304), .C2(new_n758), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n994), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n735), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n722), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n426), .A2(G50), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT50), .Z(new_n1004));
  OAI211_X1 g0804(.A(new_n680), .B(new_n461), .C1(new_n217), .C2(new_n386), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT112), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n725), .B1(new_n461), .B2(new_n236), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(G107), .B2(new_n208), .C1(new_n680), .C2(new_n730), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n981), .B(new_n1002), .C1(new_n736), .C2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n946), .B2(new_n951), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n678), .B1(new_n946), .B2(new_n718), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n947), .B2(new_n1011), .ZN(G393));
  INV_X1    g0812(.A(KEYINPUT114), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n944), .A2(new_n1013), .A3(new_n948), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n1013), .B2(new_n948), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n678), .B(new_n949), .C1(new_n1015), .C2(new_n947), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n912), .A2(new_n734), .A3(new_n913), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n736), .B1(new_n508), .B2(new_n208), .C1(new_n241), .C2(new_n726), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n744), .A2(new_n217), .B1(new_n426), .B2(new_n763), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G150), .A2(new_n783), .B1(new_n756), .B2(G159), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(KEYINPUT51), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n354), .B1(new_n758), .B2(new_n202), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n971), .A2(new_n766), .B1(new_n751), .B2(new_n386), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n747), .C2(G87), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(KEYINPUT51), .C2(new_n1020), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n761), .A2(new_n982), .B1(new_n755), .B2(new_n776), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT52), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n763), .A2(new_n545), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n274), .B1(new_n766), .B2(new_n985), .C1(new_n811), .C2(new_n758), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(G116), .C2(new_n752), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n747), .A2(G107), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n813), .C2(new_n744), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1025), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n738), .B1(new_n1034), .B2(new_n735), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1017), .A2(new_n1018), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1015), .B2(new_n951), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1016), .A2(new_n1037), .ZN(G390));
  AOI21_X1  g0838(.A(new_n888), .B1(new_n690), .B2(new_n793), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n884), .B1(new_n854), .B2(new_n862), .C1(new_n1039), .C2(new_n887), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n715), .A2(new_n835), .A3(G330), .A4(new_n793), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n845), .B1(new_n314), .B2(new_n327), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n856), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n838), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n858), .A2(new_n849), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n861), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n837), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT39), .B1(new_n872), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n892), .A2(new_n854), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1048), .B1(new_n1049), .B2(KEYINPUT39), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n890), .A2(new_n885), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1040), .B(new_n1041), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1040), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n828), .A2(new_n835), .A3(G330), .A4(new_n793), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n880), .A2(new_n882), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1051), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1061), .A2(KEYINPUT115), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n828), .A2(G330), .A3(new_n793), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n887), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n688), .B1(new_n650), .B2(new_n651), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n574), .A2(new_n577), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT90), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n580), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n640), .B1(new_n1069), .B2(new_n552), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n540), .B(new_n1065), .C1(new_n1070), .C2(new_n635), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1071), .A2(new_n669), .A3(new_n793), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1041), .A2(new_n889), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n715), .A2(G330), .A3(new_n793), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n887), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n1056), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n795), .A2(new_n889), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1064), .A2(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT116), .B1(new_n876), .B2(new_n824), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT116), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n449), .A2(new_n1080), .A3(G330), .A4(new_n828), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n898), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1054), .A2(new_n1058), .A3(new_n1062), .A4(new_n1084), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1054), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n699), .B1(new_n654), .B2(new_n663), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1071), .A2(KEYINPUT29), .A3(new_n669), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n449), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n624), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1064), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT117), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n678), .B(new_n1085), .C1(new_n1086), .C2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n354), .B(new_n808), .C1(new_n438), .C2(new_n759), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G116), .A2(new_n756), .B1(new_n959), .B2(G294), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n508), .B2(new_n763), .C1(new_n813), .C2(new_n761), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G77), .B2(new_n752), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1098), .B(new_n1101), .C1(new_n507), .C2(new_n744), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n783), .A2(G128), .B1(new_n959), .B2(G125), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n806), .B2(new_n755), .C1(new_n803), .C2(new_n758), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n274), .B(new_n1104), .C1(G159), .C2(new_n752), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n743), .A2(G150), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT53), .Z(new_n1107));
  OAI211_X1 g0907(.A(new_n1105), .B(new_n1107), .C1(new_n202), .C2(new_n748), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n763), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1102), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n738), .B1(new_n1111), .B2(new_n735), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1050), .B2(new_n733), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n304), .B2(new_n800), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1086), .B2(new_n951), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1097), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(G378));
  NAND2_X1  g0917(.A1(new_n622), .A2(new_n376), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT55), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n371), .A2(new_n845), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT56), .Z(new_n1121));
  XNOR2_X1  g0921(.A(new_n1119), .B(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n732), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n800), .A2(new_n202), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n763), .A2(new_n803), .ZN(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n761), .A2(new_n1126), .B1(new_n758), .B2(new_n806), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G150), .C2(new_n752), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n744), .B2(new_n1109), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G128), .B2(new_n756), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT59), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G41), .B1(new_n747), .B2(G159), .ZN(new_n1132));
  AOI21_X1  g0932(.A(G33), .B1(new_n959), .B2(G124), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n202), .B1(new_n257), .B2(G41), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G116), .A2(new_n783), .B1(new_n759), .B2(G97), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n813), .B2(new_n766), .C1(new_n744), .C2(new_n386), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n748), .A2(new_n279), .ZN(new_n1138));
  OR3_X1    g0938(.A1(new_n755), .A2(KEYINPUT118), .A3(new_n479), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT118), .B1(new_n755), .B2(new_n479), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n217), .C2(new_n751), .ZN(new_n1141));
  INV_X1    g0941(.A(G41), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n274), .B(new_n1142), .C1(new_n428), .C2(new_n763), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .A4(new_n1143), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT58), .Z(new_n1145));
  NAND3_X1  g0945(.A1(new_n1134), .A2(new_n1135), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n735), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n722), .B1(new_n1148), .B2(KEYINPUT119), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(KEYINPUT119), .B2(new_n1148), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1123), .A2(new_n1124), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G330), .B(new_n863), .C1(new_n873), .C2(KEYINPUT40), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n896), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1153), .A2(new_n895), .A3(new_n886), .A4(new_n893), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1122), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1155), .A2(new_n1122), .A3(new_n1156), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1152), .B1(new_n1161), .B2(new_n951), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1160), .A2(new_n1159), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n678), .B1(new_n1163), .B2(KEYINPUT57), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1162), .B1(new_n1164), .B2(new_n1168), .ZN(G375));
  AOI211_X1 g0969(.A(new_n938), .B(new_n1096), .C1(new_n1083), .C2(new_n1078), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G116), .A2(new_n759), .B1(new_n959), .B2(G303), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n813), .B2(new_n755), .C1(new_n545), .C2(new_n761), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n427), .B2(new_n752), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n743), .A2(G97), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n354), .B1(new_n764), .B2(new_n438), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1173), .A2(new_n966), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT120), .Z(new_n1177));
  AOI22_X1  g0977(.A1(new_n743), .A2(G159), .B1(G128), .B2(new_n959), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT121), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n756), .A2(G137), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n758), .B2(new_n1109), .C1(new_n806), .C2(new_n761), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n354), .B1(new_n751), .B2(new_n202), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1138), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1179), .B(new_n1183), .C1(new_n366), .C2(new_n763), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n738), .B1(new_n1185), .B2(new_n735), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n800), .A2(new_n217), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n733), .C2(new_n835), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n951), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1078), .B2(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1170), .A2(new_n1190), .ZN(G381));
  INV_X1    g0991(.A(new_n1160), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1122), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n951), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1097), .A2(new_n1115), .A3(new_n1194), .A4(new_n1151), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1163), .A2(KEYINPUT57), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n679), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1199), .A2(G396), .A3(G393), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n952), .A2(new_n1016), .A3(new_n979), .A4(new_n1037), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(G381), .A2(new_n1201), .A3(G384), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(G407));
  OAI211_X1 g1003(.A(G407), .B(G213), .C1(G343), .C2(new_n1199), .ZN(G409));
  INV_X1    g1004(.A(G213), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(G343), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  AND4_X1   g1007(.A1(new_n1207), .A2(new_n1161), .A3(new_n937), .A4(new_n1165), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1195), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1161), .A2(new_n1165), .A3(new_n937), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT122), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1206), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(G375), .A2(G378), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1216), .A2(new_n678), .A3(new_n1095), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1078), .A2(new_n1083), .A3(KEYINPUT60), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT123), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1078), .A2(new_n1083), .A3(KEYINPUT123), .A4(KEYINPUT60), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1217), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1190), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G384), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1226), .B(new_n1190), .C1(new_n1217), .C2(new_n1222), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1214), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1216), .A2(new_n678), .A3(new_n1095), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1226), .B1(new_n1230), .B2(new_n1190), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1223), .A2(G384), .A3(new_n1224), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(KEYINPUT124), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1228), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1212), .A2(new_n1213), .A3(KEYINPUT63), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT125), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT63), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1206), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1161), .A2(new_n1165), .A3(new_n1207), .A4(new_n937), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1116), .A2(new_n1211), .A3(new_n1162), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1194), .A2(new_n1151), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1238), .B(new_n1240), .C1(new_n1242), .C2(new_n1116), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1234), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1237), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1236), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1206), .A2(G2897), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1234), .B2(new_n1247), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT126), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1197), .A2(new_n1196), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1116), .B1(new_n1251), .B2(new_n1162), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1239), .A2(new_n1162), .A3(new_n1115), .A4(new_n1097), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1211), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1238), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1249), .B(new_n1250), .C1(new_n1252), .C2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(KEYINPUT125), .B(new_n1237), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1246), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n952), .A2(new_n979), .B1(new_n1016), .B2(new_n1037), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(G396), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(KEYINPUT127), .A3(new_n1201), .A4(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1263), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1201), .A2(KEYINPUT127), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1266), .B2(new_n1261), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT62), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1212), .A2(new_n1213), .A3(new_n1270), .A4(new_n1234), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1257), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1268), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1268), .A2(new_n1250), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1260), .A2(new_n1268), .B1(new_n1274), .B2(new_n1275), .ZN(G405));
  OAI22_X1  g1076(.A1(new_n1252), .A2(new_n1198), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1213), .A2(new_n1199), .A3(new_n1234), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(new_n1268), .Z(G402));
endmodule


