

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745;

  AND2_X1 U365 ( .A1(n364), .A2(n362), .ZN(n343) );
  OR2_X1 U366 ( .A1(n705), .A2(G902), .ZN(n415) );
  AND2_X1 U367 ( .A1(n354), .A2(KEYINPUT19), .ZN(n353) );
  NOR2_X1 U368 ( .A1(n529), .A2(n530), .ZN(n531) );
  XNOR2_X2 U369 ( .A(n715), .B(n448), .ZN(n382) );
  XNOR2_X2 U370 ( .A(n454), .B(n371), .ZN(n715) );
  XNOR2_X2 U371 ( .A(n585), .B(n584), .ZN(n719) );
  INV_X1 U372 ( .A(G953), .ZN(n735) );
  NOR2_X2 U373 ( .A1(n540), .A2(n547), .ZN(n541) );
  NOR2_X2 U374 ( .A1(n676), .A2(n578), .ZN(n558) );
  XNOR2_X2 U375 ( .A(n556), .B(n555), .ZN(n676) );
  XNOR2_X2 U376 ( .A(G116), .B(G113), .ZN(n368) );
  XNOR2_X2 U377 ( .A(n409), .B(KEYINPUT4), .ZN(n443) );
  NOR2_X1 U378 ( .A1(n357), .A2(n389), .ZN(n352) );
  AND2_X1 U379 ( .A1(n359), .A2(n358), .ZN(n357) );
  NOR2_X1 U380 ( .A1(n524), .A2(n500), .ZN(n526) );
  AND2_X1 U381 ( .A1(n678), .A2(n516), .ZN(n575) );
  AND2_X1 U382 ( .A1(n678), .A2(n552), .ZN(n573) );
  NOR2_X1 U383 ( .A1(n353), .A2(n352), .ZN(n351) );
  BUF_X1 U384 ( .A(n552), .Z(n679) );
  XNOR2_X1 U385 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U386 ( .A(n481), .B(n480), .ZN(n505) );
  NOR2_X2 U387 ( .A1(n528), .A2(n527), .ZN(n656) );
  XNOR2_X2 U388 ( .A(n382), .B(n381), .ZN(n610) );
  XNOR2_X2 U389 ( .A(n443), .B(n442), .ZN(n730) );
  XNOR2_X2 U390 ( .A(n730), .B(G146), .ZN(n460) );
  XNOR2_X1 U391 ( .A(n516), .B(KEYINPUT1), .ZN(n552) );
  XNOR2_X1 U392 ( .A(G134), .B(G116), .ZN(n406) );
  NOR2_X1 U393 ( .A1(n363), .A2(n513), .ZN(n362) );
  NOR2_X1 U394 ( .A1(n453), .A2(n566), .ZN(n363) );
  NAND2_X1 U395 ( .A1(n361), .A2(KEYINPUT104), .ZN(n360) );
  BUF_X1 U396 ( .A(n505), .Z(n682) );
  NOR2_X1 U397 ( .A1(n388), .A2(KEYINPUT19), .ZN(n350) );
  NAND2_X1 U398 ( .A1(n386), .A2(n595), .ZN(n358) );
  NOR2_X1 U399 ( .A1(n679), .A2(KEYINPUT104), .ZN(n365) );
  OR2_X1 U400 ( .A1(n620), .A2(G902), .ZN(n452) );
  XNOR2_X1 U401 ( .A(n368), .B(G119), .ZN(n370) );
  OR2_X1 U402 ( .A1(n602), .A2(G902), .ZN(n462) );
  BUF_X1 U403 ( .A(n557), .Z(n578) );
  XNOR2_X1 U404 ( .A(n413), .B(n412), .ZN(n705) );
  XNOR2_X1 U405 ( .A(n610), .B(n612), .ZN(n613) );
  AND2_X1 U406 ( .A1(n605), .A2(G953), .ZN(n714) );
  XNOR2_X1 U407 ( .A(n564), .B(n563), .ZN(n633) );
  NAND2_X1 U408 ( .A1(n343), .A2(n360), .ZN(n569) );
  INV_X1 U409 ( .A(n679), .ZN(n453) );
  XNOR2_X1 U410 ( .A(n370), .B(n369), .ZN(n454) );
  AND2_X1 U411 ( .A1(n633), .A2(n565), .ZN(n344) );
  AND2_X1 U412 ( .A1(n582), .A2(n581), .ZN(n345) );
  NAND2_X1 U413 ( .A1(n351), .A2(n348), .ZN(n518) );
  XNOR2_X1 U414 ( .A(n540), .B(KEYINPUT105), .ZN(n636) );
  NAND2_X1 U415 ( .A1(n634), .A2(n344), .ZN(n347) );
  NAND2_X1 U416 ( .A1(n346), .A2(n345), .ZN(n585) );
  XNOR2_X1 U417 ( .A(n347), .B(n572), .ZN(n346) );
  NAND2_X1 U418 ( .A1(n571), .A2(n570), .ZN(n634) );
  NAND2_X1 U419 ( .A1(n357), .A2(n355), .ZN(n500) );
  NAND2_X1 U420 ( .A1(n357), .A2(n349), .ZN(n348) );
  AND2_X1 U421 ( .A1(n355), .A2(n350), .ZN(n349) );
  NAND2_X1 U422 ( .A1(n355), .A2(n668), .ZN(n354) );
  OR2_X2 U423 ( .A1(n610), .A2(n356), .ZN(n355) );
  OR2_X1 U424 ( .A1(n386), .A2(n595), .ZN(n356) );
  NAND2_X1 U425 ( .A1(n610), .A2(n386), .ZN(n359) );
  NAND2_X1 U426 ( .A1(n366), .A2(n453), .ZN(n567) );
  INV_X1 U427 ( .A(n366), .ZN(n361) );
  NAND2_X1 U428 ( .A1(n366), .A2(n365), .ZN(n364) );
  INV_X1 U429 ( .A(n485), .ZN(n366) );
  XNOR2_X2 U430 ( .A(n472), .B(n471), .ZN(n729) );
  XOR2_X1 U431 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n367) );
  INV_X1 U432 ( .A(KEYINPUT48), .ZN(n545) );
  XNOR2_X1 U433 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n502) );
  INV_X1 U434 ( .A(KEYINPUT44), .ZN(n572) );
  INV_X1 U435 ( .A(KEYINPUT19), .ZN(n389) );
  XNOR2_X1 U436 ( .A(n411), .B(n410), .ZN(n412) );
  INV_X1 U437 ( .A(n636), .ZN(n650) );
  XNOR2_X1 U438 ( .A(G101), .B(KEYINPUT3), .ZN(n369) );
  INV_X1 U439 ( .A(G122), .ZN(n631) );
  XNOR2_X1 U440 ( .A(n631), .B(G107), .ZN(n402) );
  XNOR2_X1 U441 ( .A(n402), .B(KEYINPUT16), .ZN(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT87), .B(G110), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n372), .B(G104), .ZN(n716) );
  XNOR2_X1 U444 ( .A(n716), .B(KEYINPUT74), .ZN(n448) );
  XNOR2_X2 U445 ( .A(KEYINPUT77), .B(G143), .ZN(n374) );
  INV_X1 U446 ( .A(G128), .ZN(n373) );
  XNOR2_X2 U447 ( .A(n374), .B(n373), .ZN(n409) );
  XNOR2_X2 U448 ( .A(G146), .B(G125), .ZN(n418) );
  XNOR2_X1 U449 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n375) );
  XNOR2_X1 U450 ( .A(n418), .B(n375), .ZN(n379) );
  XNOR2_X1 U451 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n377) );
  NAND2_X1 U452 ( .A1(n735), .A2(G224), .ZN(n376) );
  XNOR2_X1 U453 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U454 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U455 ( .A(n443), .B(n380), .ZN(n381) );
  XNOR2_X1 U456 ( .A(G902), .B(KEYINPUT15), .ZN(n590) );
  INV_X1 U457 ( .A(n590), .ZN(n595) );
  INV_X1 U458 ( .A(G902), .ZN(n428) );
  INV_X1 U459 ( .A(G237), .ZN(n383) );
  NAND2_X1 U460 ( .A1(n428), .A2(n383), .ZN(n387) );
  NAND2_X1 U461 ( .A1(n387), .A2(G210), .ZN(n385) );
  INV_X1 U462 ( .A(KEYINPUT89), .ZN(n384) );
  XNOR2_X1 U463 ( .A(n385), .B(n384), .ZN(n386) );
  NAND2_X1 U464 ( .A1(n387), .A2(G214), .ZN(n668) );
  INV_X1 U465 ( .A(n668), .ZN(n388) );
  NAND2_X1 U466 ( .A1(G234), .A2(G237), .ZN(n390) );
  XNOR2_X1 U467 ( .A(n390), .B(KEYINPUT14), .ZN(n393) );
  NAND2_X1 U468 ( .A1(G952), .A2(n393), .ZN(n696) );
  NOR2_X1 U469 ( .A1(n696), .A2(G953), .ZN(n392) );
  INV_X1 U470 ( .A(KEYINPUT90), .ZN(n391) );
  XNOR2_X1 U471 ( .A(n392), .B(n391), .ZN(n492) );
  NAND2_X1 U472 ( .A1(G902), .A2(n393), .ZN(n489) );
  NOR2_X1 U473 ( .A1(G898), .A2(n735), .ZN(n394) );
  XNOR2_X1 U474 ( .A(KEYINPUT91), .B(n394), .ZN(n717) );
  NOR2_X1 U475 ( .A1(n489), .A2(n717), .ZN(n396) );
  INV_X1 U476 ( .A(KEYINPUT92), .ZN(n395) );
  XNOR2_X1 U477 ( .A(n396), .B(n395), .ZN(n397) );
  NAND2_X1 U478 ( .A1(n492), .A2(n397), .ZN(n398) );
  NAND2_X1 U479 ( .A1(n518), .A2(n398), .ZN(n401) );
  INV_X1 U480 ( .A(KEYINPUT83), .ZN(n399) );
  XNOR2_X1 U481 ( .A(n399), .B(KEYINPUT0), .ZN(n400) );
  XNOR2_X1 U482 ( .A(n401), .B(n400), .ZN(n557) );
  INV_X1 U483 ( .A(n557), .ZN(n438) );
  XOR2_X1 U484 ( .A(n402), .B(KEYINPUT100), .Z(n405) );
  NAND2_X1 U485 ( .A1(G234), .A2(n735), .ZN(n403) );
  XOR2_X1 U486 ( .A(KEYINPUT8), .B(n403), .Z(n473) );
  NAND2_X1 U487 ( .A1(G217), .A2(n473), .ZN(n404) );
  XNOR2_X1 U488 ( .A(n405), .B(n404), .ZN(n413) );
  XNOR2_X1 U489 ( .A(n367), .B(n406), .ZN(n408) );
  XOR2_X1 U490 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n407) );
  XNOR2_X1 U491 ( .A(n408), .B(n407), .ZN(n411) );
  INV_X1 U492 ( .A(n409), .ZN(n410) );
  INV_X1 U493 ( .A(G478), .ZN(n414) );
  XNOR2_X2 U494 ( .A(n415), .B(n414), .ZN(n560) );
  XOR2_X1 U495 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n417) );
  NOR2_X1 U496 ( .A1(G953), .A2(G237), .ZN(n455) );
  NAND2_X1 U497 ( .A1(G214), .A2(n455), .ZN(n416) );
  XNOR2_X1 U498 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U499 ( .A(n418), .B(KEYINPUT10), .ZN(n470) );
  XNOR2_X1 U500 ( .A(n419), .B(n470), .ZN(n427) );
  XOR2_X1 U501 ( .A(G140), .B(G104), .Z(n421) );
  XNOR2_X1 U502 ( .A(G143), .B(G131), .ZN(n420) );
  XNOR2_X1 U503 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U504 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n423) );
  XNOR2_X1 U505 ( .A(G113), .B(G122), .ZN(n422) );
  XNOR2_X1 U506 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U507 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U508 ( .A(n427), .B(n426), .ZN(n626) );
  NAND2_X1 U509 ( .A1(n626), .A2(n428), .ZN(n432) );
  XOR2_X1 U510 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n430) );
  XNOR2_X1 U511 ( .A(KEYINPUT98), .B(G475), .ZN(n429) );
  XOR2_X1 U512 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U513 ( .A(n432), .B(n431), .ZN(n520) );
  INV_X1 U514 ( .A(n520), .ZN(n559) );
  NAND2_X1 U515 ( .A1(n560), .A2(n559), .ZN(n671) );
  NAND2_X1 U516 ( .A1(n590), .A2(G234), .ZN(n433) );
  XNOR2_X1 U517 ( .A(n433), .B(KEYINPUT20), .ZN(n477) );
  AND2_X1 U518 ( .A1(n477), .A2(G221), .ZN(n436) );
  INV_X1 U519 ( .A(KEYINPUT94), .ZN(n434) );
  XNOR2_X1 U520 ( .A(n434), .B(KEYINPUT21), .ZN(n435) );
  XNOR2_X1 U521 ( .A(n436), .B(n435), .ZN(n504) );
  NOR2_X1 U522 ( .A1(n671), .A2(n504), .ZN(n437) );
  NAND2_X1 U523 ( .A1(n438), .A2(n437), .ZN(n439) );
  XNOR2_X1 U524 ( .A(n439), .B(KEYINPUT22), .ZN(n485) );
  XOR2_X1 U525 ( .A(G137), .B(KEYINPUT71), .Z(n441) );
  XNOR2_X1 U526 ( .A(G131), .B(G134), .ZN(n440) );
  XNOR2_X1 U527 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U528 ( .A(KEYINPUT70), .B(G140), .Z(n471) );
  INV_X1 U529 ( .A(G101), .ZN(n444) );
  XNOR2_X1 U530 ( .A(n444), .B(G107), .ZN(n446) );
  NAND2_X1 U531 ( .A1(G227), .A2(n735), .ZN(n445) );
  XNOR2_X1 U532 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n471), .B(n447), .ZN(n449) );
  XNOR2_X1 U534 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U535 ( .A(n460), .B(n450), .ZN(n620) );
  XOR2_X1 U536 ( .A(KEYINPUT73), .B(G469), .Z(n451) );
  XNOR2_X2 U537 ( .A(n452), .B(n451), .ZN(n516) );
  XOR2_X1 U538 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n457) );
  NAND2_X1 U539 ( .A1(n455), .A2(G210), .ZN(n456) );
  XNOR2_X1 U540 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U541 ( .A(n454), .B(n458), .ZN(n459) );
  XNOR2_X1 U542 ( .A(n460), .B(n459), .ZN(n602) );
  XNOR2_X1 U543 ( .A(G472), .B(KEYINPUT75), .ZN(n461) );
  XNOR2_X2 U544 ( .A(n462), .B(n461), .ZN(n576) );
  INV_X1 U545 ( .A(KEYINPUT6), .ZN(n463) );
  XNOR2_X1 U546 ( .A(n576), .B(n463), .ZN(n553) );
  XNOR2_X1 U547 ( .A(G137), .B(G110), .ZN(n465) );
  INV_X1 U548 ( .A(KEYINPUT24), .ZN(n464) );
  XNOR2_X1 U549 ( .A(n465), .B(n464), .ZN(n467) );
  XOR2_X1 U550 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n466) );
  XNOR2_X1 U551 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U552 ( .A(G128), .B(G119), .ZN(n468) );
  XOR2_X1 U553 ( .A(n469), .B(n468), .Z(n476) );
  INV_X1 U554 ( .A(n470), .ZN(n472) );
  NAND2_X1 U555 ( .A1(G221), .A2(n473), .ZN(n474) );
  XNOR2_X1 U556 ( .A(n729), .B(n474), .ZN(n475) );
  XNOR2_X1 U557 ( .A(n476), .B(n475), .ZN(n710) );
  NOR2_X1 U558 ( .A1(n710), .A2(G902), .ZN(n481) );
  XOR2_X1 U559 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n479) );
  AND2_X1 U560 ( .A1(G217), .A2(n477), .ZN(n478) );
  XNOR2_X1 U561 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U562 ( .A1(n553), .A2(n682), .ZN(n482) );
  OR2_X1 U563 ( .A1(n567), .A2(n482), .ZN(n581) );
  XNOR2_X1 U564 ( .A(n581), .B(G101), .ZN(G3) );
  XNOR2_X1 U565 ( .A(n679), .B(KEYINPUT85), .ZN(n528) );
  INV_X1 U566 ( .A(n682), .ZN(n570) );
  NAND2_X1 U567 ( .A1(n553), .A2(n570), .ZN(n483) );
  OR2_X1 U568 ( .A1(n528), .A2(n483), .ZN(n484) );
  OR2_X1 U569 ( .A1(n485), .A2(n484), .ZN(n488) );
  INV_X1 U570 ( .A(KEYINPUT65), .ZN(n486) );
  XNOR2_X1 U571 ( .A(n486), .B(KEYINPUT32), .ZN(n487) );
  XNOR2_X1 U572 ( .A(n488), .B(n487), .ZN(n565) );
  XNOR2_X1 U573 ( .A(n565), .B(G119), .ZN(G21) );
  NAND2_X1 U574 ( .A1(n560), .A2(n520), .ZN(n540) );
  NOR2_X1 U575 ( .A1(G900), .A2(n489), .ZN(n490) );
  NAND2_X1 U576 ( .A1(G953), .A2(n490), .ZN(n491) );
  NAND2_X1 U577 ( .A1(n492), .A2(n491), .ZN(n538) );
  NOR2_X1 U578 ( .A1(n505), .A2(n504), .ZN(n493) );
  NAND2_X1 U579 ( .A1(n538), .A2(n493), .ZN(n494) );
  XNOR2_X1 U580 ( .A(KEYINPUT72), .B(n494), .ZN(n514) );
  INV_X1 U581 ( .A(n514), .ZN(n495) );
  NAND2_X1 U582 ( .A1(n636), .A2(n495), .ZN(n496) );
  NOR2_X1 U583 ( .A1(n553), .A2(n496), .ZN(n497) );
  XNOR2_X1 U584 ( .A(n497), .B(KEYINPUT106), .ZN(n498) );
  NAND2_X1 U585 ( .A1(n498), .A2(n668), .ZN(n524) );
  NOR2_X1 U586 ( .A1(n679), .A2(n524), .ZN(n499) );
  XOR2_X1 U587 ( .A(n499), .B(KEYINPUT43), .Z(n501) );
  NAND2_X1 U588 ( .A1(n501), .A2(n500), .ZN(n549) );
  XNOR2_X1 U589 ( .A(n549), .B(G140), .ZN(G42) );
  INV_X1 U590 ( .A(n576), .ZN(n512) );
  NAND2_X1 U591 ( .A1(n668), .A2(n512), .ZN(n503) );
  XNOR2_X1 U592 ( .A(n503), .B(n502), .ZN(n507) );
  INV_X1 U593 ( .A(n504), .ZN(n681) );
  NAND2_X1 U594 ( .A1(n505), .A2(n681), .ZN(n506) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(n506), .Z(n678) );
  NAND2_X1 U596 ( .A1(n507), .A2(n575), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n538), .A2(n520), .ZN(n508) );
  NOR2_X1 U598 ( .A1(n536), .A2(n508), .ZN(n510) );
  NOR2_X1 U599 ( .A1(n500), .A2(n560), .ZN(n509) );
  NAND2_X1 U600 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U601 ( .A(KEYINPUT108), .B(n511), .ZN(n742) );
  BUF_X1 U602 ( .A(n512), .Z(n513) );
  NOR2_X1 U603 ( .A1(n514), .A2(n576), .ZN(n515) );
  XNOR2_X1 U604 ( .A(KEYINPUT28), .B(n515), .ZN(n517) );
  NAND2_X1 U605 ( .A1(n517), .A2(n516), .ZN(n533) );
  INV_X1 U606 ( .A(n518), .ZN(n519) );
  NOR2_X1 U607 ( .A1(n533), .A2(n519), .ZN(n648) );
  NOR2_X1 U608 ( .A1(n520), .A2(n560), .ZN(n521) );
  XOR2_X1 U609 ( .A(n521), .B(KEYINPUT103), .Z(n645) );
  INV_X1 U610 ( .A(n645), .ZN(n653) );
  NAND2_X1 U611 ( .A1(n540), .A2(n653), .ZN(n579) );
  INV_X1 U612 ( .A(n579), .ZN(n673) );
  NOR2_X1 U613 ( .A1(KEYINPUT69), .A2(n673), .ZN(n522) );
  NAND2_X1 U614 ( .A1(n648), .A2(n522), .ZN(n523) );
  XNOR2_X1 U615 ( .A(KEYINPUT47), .B(n523), .ZN(n530) );
  XNOR2_X1 U616 ( .A(KEYINPUT36), .B(KEYINPUT109), .ZN(n525) );
  XNOR2_X1 U617 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U618 ( .A(n656), .B(KEYINPUT82), .ZN(n529) );
  AND2_X1 U619 ( .A1(n742), .A2(n531), .ZN(n544) );
  XOR2_X1 U620 ( .A(KEYINPUT38), .B(n500), .Z(n535) );
  INV_X1 U621 ( .A(n535), .ZN(n669) );
  NAND2_X1 U622 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U623 ( .A1(n672), .A2(n671), .ZN(n532) );
  XNOR2_X1 U624 ( .A(n532), .B(KEYINPUT41), .ZN(n698) );
  NOR2_X1 U625 ( .A1(n698), .A2(n533), .ZN(n534) );
  XNOR2_X1 U626 ( .A(n534), .B(KEYINPUT42), .ZN(n745) );
  NOR2_X1 U627 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U628 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U629 ( .A(KEYINPUT39), .B(n539), .Z(n547) );
  XNOR2_X1 U630 ( .A(KEYINPUT40), .B(n541), .ZN(n744) );
  NOR2_X1 U631 ( .A1(n745), .A2(n744), .ZN(n542) );
  XNOR2_X1 U632 ( .A(n542), .B(KEYINPUT46), .ZN(n543) );
  NAND2_X1 U633 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U634 ( .A(n546), .B(n545), .ZN(n551) );
  INV_X1 U635 ( .A(n547), .ZN(n548) );
  NAND2_X1 U636 ( .A1(n548), .A2(n645), .ZN(n659) );
  AND2_X1 U637 ( .A1(n659), .A2(n549), .ZN(n550) );
  NAND2_X1 U638 ( .A1(n551), .A2(n550), .ZN(n727) );
  INV_X1 U639 ( .A(n553), .ZN(n554) );
  NAND2_X1 U640 ( .A1(n573), .A2(n554), .ZN(n556) );
  INV_X1 U641 ( .A(KEYINPUT33), .ZN(n555) );
  XNOR2_X1 U642 ( .A(n558), .B(KEYINPUT34), .ZN(n562) );
  NOR2_X1 U643 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U644 ( .A1(n562), .A2(n561), .ZN(n564) );
  INV_X1 U645 ( .A(KEYINPUT35), .ZN(n563) );
  INV_X1 U646 ( .A(KEYINPUT104), .ZN(n566) );
  INV_X1 U647 ( .A(KEYINPUT66), .ZN(n568) );
  XNOR2_X1 U648 ( .A(n569), .B(n568), .ZN(n571) );
  NAND2_X1 U649 ( .A1(n573), .A2(n513), .ZN(n687) );
  NOR2_X1 U650 ( .A1(n687), .A2(n578), .ZN(n574) );
  XNOR2_X1 U651 ( .A(n574), .B(KEYINPUT31), .ZN(n652) );
  NAND2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n639) );
  NAND2_X1 U654 ( .A1(n652), .A2(n639), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n582) );
  INV_X1 U656 ( .A(KEYINPUT64), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT45), .ZN(n584) );
  NOR2_X2 U658 ( .A1(n727), .A2(n719), .ZN(n660) );
  XNOR2_X1 U659 ( .A(n660), .B(KEYINPUT79), .ZN(n593) );
  NAND2_X1 U660 ( .A1(KEYINPUT2), .A2(KEYINPUT80), .ZN(n591) );
  INV_X1 U661 ( .A(KEYINPUT80), .ZN(n586) );
  NAND2_X1 U662 ( .A1(KEYINPUT2), .A2(n586), .ZN(n588) );
  INV_X1 U663 ( .A(KEYINPUT79), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n594) );
  AND2_X1 U666 ( .A1(n591), .A2(n594), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n600) );
  INV_X1 U668 ( .A(n594), .ZN(n596) );
  OR2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n660), .A2(KEYINPUT2), .ZN(n597) );
  AND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n599) );
  AND2_X2 U672 ( .A1(n600), .A2(n599), .ZN(n624) );
  NAND2_X1 U673 ( .A1(n624), .A2(G472), .ZN(n604) );
  XNOR2_X1 U674 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n606) );
  INV_X1 U677 ( .A(G952), .ZN(n605) );
  NOR2_X1 U678 ( .A1(n606), .A2(n714), .ZN(n609) );
  XNOR2_X1 U679 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT86), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n609), .B(n608), .ZN(G57) );
  NAND2_X1 U682 ( .A1(n624), .A2(G210), .ZN(n614) );
  XNOR2_X1 U683 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n611) );
  XNOR2_X1 U684 ( .A(n611), .B(KEYINPUT55), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n614), .B(n613), .ZN(n615) );
  NOR2_X1 U686 ( .A1(n615), .A2(n714), .ZN(n617) );
  XOR2_X1 U687 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(G51) );
  INV_X1 U689 ( .A(n624), .ZN(n618) );
  INV_X1 U690 ( .A(n618), .ZN(n709) );
  NAND2_X1 U691 ( .A1(n709), .A2(G469), .ZN(n622) );
  XOR2_X1 U692 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n619) );
  XNOR2_X1 U693 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X1 U695 ( .A1(n623), .A2(n714), .ZN(G54) );
  NAND2_X1 U696 ( .A1(n624), .A2(G475), .ZN(n628) );
  XOR2_X1 U697 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n625) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X1 U699 ( .A1(n629), .A2(n714), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U701 ( .A(n631), .B(KEYINPUT127), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n633), .B(n632), .ZN(G24) );
  XOR2_X1 U703 ( .A(G110), .B(KEYINPUT115), .Z(n635) );
  XNOR2_X1 U704 ( .A(n634), .B(n635), .ZN(G12) );
  NOR2_X1 U705 ( .A1(n639), .A2(n650), .ZN(n637) );
  XOR2_X1 U706 ( .A(KEYINPUT112), .B(n637), .Z(n638) );
  XNOR2_X1 U707 ( .A(G104), .B(n638), .ZN(G6) );
  NOR2_X1 U708 ( .A1(n639), .A2(n653), .ZN(n644) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n641) );
  XNOR2_X1 U710 ( .A(G107), .B(KEYINPUT113), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U712 ( .A(KEYINPUT26), .B(n642), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n644), .B(n643), .ZN(G9) );
  XOR2_X1 U714 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n645), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G30) );
  NAND2_X1 U717 ( .A1(n648), .A2(n636), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(G146), .ZN(G48) );
  NOR2_X1 U719 ( .A1(n650), .A2(n652), .ZN(n651) );
  XOR2_X1 U720 ( .A(G113), .B(n651), .Z(G15) );
  NOR2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U722 ( .A(G116), .B(KEYINPUT117), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(G18) );
  XNOR2_X1 U724 ( .A(n656), .B(KEYINPUT118), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT37), .ZN(n658) );
  XNOR2_X1 U726 ( .A(G125), .B(n658), .ZN(G27) );
  XNOR2_X1 U727 ( .A(G134), .B(n659), .ZN(G36) );
  BUF_X1 U728 ( .A(n660), .Z(n661) );
  INV_X1 U729 ( .A(n661), .ZN(n663) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n662) );
  NAND2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n667) );
  INV_X1 U732 ( .A(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n664), .A2(KEYINPUT78), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n661), .A2(n665), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n702) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n693) );
  OR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U742 ( .A(n680), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U744 ( .A(KEYINPUT49), .B(n683), .Z(n684) );
  NOR2_X1 U745 ( .A1(n513), .A2(n684), .ZN(n685) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n688) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U748 ( .A(KEYINPUT51), .B(n689), .ZN(n690) );
  NOR2_X1 U749 ( .A1(n698), .A2(n690), .ZN(n691) );
  XOR2_X1 U750 ( .A(KEYINPUT119), .B(n691), .Z(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n694), .B(KEYINPUT52), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n697), .B(KEYINPUT120), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n698), .A2(n676), .ZN(n699) );
  NOR2_X1 U756 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U757 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U758 ( .A1(n703), .A2(G953), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n704), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U760 ( .A1(n709), .A2(G478), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n705), .B(KEYINPUT122), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U763 ( .A1(n714), .A2(n708), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n709), .A2(G217), .ZN(n712) );
  XOR2_X1 U765 ( .A(n710), .B(KEYINPUT123), .Z(n711) );
  XNOR2_X1 U766 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(G66) );
  XOR2_X1 U768 ( .A(n715), .B(n716), .Z(n718) );
  NAND2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n726) );
  OR2_X1 U770 ( .A1(n719), .A2(G953), .ZN(n724) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n720), .B(KEYINPUT124), .ZN(n721) );
  XNOR2_X1 U773 ( .A(KEYINPUT61), .B(n721), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n722), .A2(G898), .ZN(n723) );
  AND2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n726), .B(n725), .ZN(G69) );
  BUF_X1 U777 ( .A(n727), .Z(n728) );
  XOR2_X1 U778 ( .A(KEYINPUT126), .B(n728), .Z(n734) );
  XNOR2_X1 U779 ( .A(n729), .B(KEYINPUT125), .ZN(n732) );
  INV_X1 U780 ( .A(n730), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(n737) );
  INV_X1 U782 ( .A(n737), .ZN(n733) );
  XOR2_X1 U783 ( .A(n734), .B(n733), .Z(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n741) );
  XOR2_X1 U785 ( .A(G227), .B(n737), .Z(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U789 ( .A(G143), .B(n742), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n743), .B(KEYINPUT116), .ZN(G45) );
  XOR2_X1 U791 ( .A(G131), .B(n744), .Z(G33) );
  XOR2_X1 U792 ( .A(G137), .B(n745), .Z(G39) );
endmodule

