//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT78), .ZN(new_n204));
  OR2_X1    g003(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n204), .B(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT79), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(G155gat), .B2(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT84), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT85), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n215), .B(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n214), .B(new_n218), .C1(new_n220), .C2(new_n217), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n215), .A2(new_n217), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT84), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(new_n214), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT86), .B(KEYINPUT3), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(G228gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n212), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT3), .B1(new_n232), .B2(new_n228), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n230), .B(new_n231), .C1(new_n225), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n225), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n228), .B1(new_n211), .B2(new_n203), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n202), .B1(new_n209), .B2(new_n210), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n226), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n229), .A2(new_n212), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n234), .B1(new_n231), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G78gat), .B(G106gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT31), .B(G50gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(G22gat), .ZN(new_n244));
  INV_X1    g043(.A(G22gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT88), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n240), .B(new_n247), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n250));
  INV_X1    g049(.A(G113gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G120gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT71), .B(G120gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(new_n251), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n255));
  XNOR2_X1  g054(.A(G127gat), .B(G134gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n251), .A2(G120gat), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT1), .B1(new_n260), .B2(new_n252), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n261), .A2(new_n256), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n254), .A2(KEYINPUT72), .A3(new_n255), .A4(new_n256), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OR3_X1    g063(.A1(new_n235), .A2(new_n250), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n227), .B(new_n264), .C1(new_n266), .C2(new_n225), .ZN(new_n267));
  NAND2_X1  g066(.A1(G225gat), .A2(G233gat), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n225), .A2(new_n262), .A3(new_n259), .A4(new_n263), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n250), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n265), .A2(new_n267), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n235), .A2(new_n264), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n272), .B2(new_n269), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT87), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT5), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n225), .B(new_n264), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n276), .A2(KEYINPUT87), .A3(new_n268), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT89), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT89), .B1(new_n278), .B2(new_n280), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G57gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G85gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  NOR3_X1   g085(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n265), .A2(new_n267), .A3(new_n270), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(G225gat), .A3(G233gat), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n289), .A2(KEYINPUT39), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n276), .A2(new_n268), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(KEYINPUT39), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n293), .A2(KEYINPUT40), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(KEYINPUT40), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n287), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT28), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT68), .B(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT27), .ZN(new_n301));
  OR2_X1    g100(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n302));
  AOI21_X1  g101(.A(G190gat), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n299), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  INV_X1    g114(.A(G176gat), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n318));
  OAI211_X1 g117(.A(KEYINPUT23), .B(new_n315), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G183gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n298), .ZN(new_n326));
  NAND4_X1  g125(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n322), .A2(new_n324), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n307), .A2(KEYINPUT23), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n319), .A2(new_n328), .A3(new_n311), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(G183gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n298), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n320), .A2(KEYINPUT67), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n339), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n324), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n310), .B1(KEYINPUT23), .B2(new_n307), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n329), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n307), .A2(KEYINPUT23), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT66), .B1(new_n346), .B2(new_n310), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n342), .A2(new_n345), .A3(KEYINPUT25), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n314), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT81), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT69), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n333), .A2(new_n348), .A3(KEYINPUT69), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT80), .B1(new_n361), .B2(new_n314), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n333), .A2(new_n348), .A3(KEYINPUT69), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT69), .B1(new_n333), .B2(new_n348), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT80), .B(new_n314), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n228), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n357), .B1(new_n367), .B2(new_n351), .ZN(new_n368));
  INV_X1    g167(.A(new_n213), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT82), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n352), .B1(new_n362), .B2(new_n366), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n314), .B2(new_n349), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT83), .B1(new_n372), .B2(new_n352), .ZN(new_n373));
  OR3_X1    g172(.A1(new_n372), .A2(KEYINPUT83), .A3(new_n352), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n232), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n314), .B1(new_n363), .B2(new_n364), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n379), .B2(new_n365), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n354), .B(new_n356), .C1(new_n380), .C2(new_n352), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n213), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n370), .A2(new_n376), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385));
  INV_X1    g184(.A(G64gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G92gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  OR3_X1    g188(.A1(new_n384), .A2(KEYINPUT30), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(new_n389), .ZN(new_n391));
  INV_X1    g190(.A(new_n389), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n370), .A2(new_n376), .A3(new_n383), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(KEYINPUT30), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n296), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT37), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n384), .A2(new_n396), .ZN(new_n397));
  OAI221_X1 g196(.A(KEYINPUT37), .B1(new_n381), .B2(new_n213), .C1(new_n375), .C2(new_n232), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT38), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n389), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n278), .A2(new_n280), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n402), .A2(new_n403), .A3(new_n286), .ZN(new_n404));
  OR3_X1    g203(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT6), .B1(new_n402), .B2(new_n286), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n370), .A2(new_n376), .A3(new_n383), .A4(KEYINPUT37), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n392), .B1(new_n397), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n393), .B1(new_n410), .B2(new_n400), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n249), .B(new_n395), .C1(new_n408), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n264), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n361), .A2(new_n314), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G227gat), .ZN(new_n416));
  INV_X1    g215(.A(G233gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n377), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n264), .B(new_n413), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n415), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT75), .B(G71gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G99gat), .ZN(new_n423));
  XOR2_X1   g222(.A(G15gat), .B(G43gat), .Z(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT33), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(KEYINPUT32), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(KEYINPUT74), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(KEYINPUT32), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n425), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT74), .B1(new_n421), .B2(new_n428), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT34), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n415), .B1(new_n419), .B2(new_n420), .ZN(new_n436));
  INV_X1    g235(.A(new_n418), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n435), .A3(new_n437), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n433), .A2(new_n434), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n432), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n442), .A2(new_n430), .A3(new_n425), .A4(new_n429), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n434), .A3(new_n440), .ZN(new_n444));
  INV_X1    g243(.A(new_n440), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT76), .B1(new_n445), .B2(new_n438), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n443), .A2(new_n444), .A3(new_n446), .A4(new_n427), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT36), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n441), .A2(KEYINPUT36), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n394), .A2(new_n390), .ZN(new_n453));
  INV_X1    g252(.A(new_n402), .ZN(new_n454));
  INV_X1    g253(.A(new_n286), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n404), .B1(new_n456), .B2(new_n406), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n452), .B1(new_n459), .B2(new_n248), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n248), .B1(new_n441), .B2(new_n447), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  INV_X1    g263(.A(new_n404), .ZN(new_n465));
  INV_X1    g264(.A(new_n406), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n287), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n453), .A2(new_n464), .A3(new_n467), .A4(new_n461), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n412), .A2(new_n460), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G78gat), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n470), .A2(KEYINPUT98), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT99), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT97), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(G57gat), .B2(new_n386), .ZN(new_n476));
  INV_X1    g275(.A(G57gat), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n477), .A2(KEYINPUT97), .A3(G64gat), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n476), .A2(new_n478), .B1(G57gat), .B2(new_n386), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(KEYINPUT98), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n471), .A2(new_n474), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n470), .ZN(new_n482));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(new_n472), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT21), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(new_n207), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n487), .B(new_n489), .Z(new_n490));
  XNOR2_X1  g289(.A(G127gat), .B(G155gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494));
  INV_X1    g293(.A(G1gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT16), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G8gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT94), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n496), .B(new_n498), .C1(new_n495), .C2(new_n494), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n497), .A2(KEYINPUT94), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n486), .B2(new_n485), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(G183gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(G183gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G231gat), .A2(G233gat), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n493), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n513), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n492), .A3(new_n511), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G134gat), .B(G162gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(KEYINPUT103), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G29gat), .ZN(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT14), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G29gat), .A2(G36gat), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G50gat), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT15), .B1(new_n531), .B2(G43gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(G43gat), .B2(new_n531), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n530), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT92), .B(G43gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT93), .A3(new_n531), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G43gat), .B2(new_n531), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT93), .B1(new_n536), .B2(new_n531), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n535), .B(new_n528), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n542));
  NAND2_X1  g341(.A1(G85gat), .A2(G92gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT104), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n543), .B(KEYINPUT104), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(G85gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(KEYINPUT8), .A2(new_n550), .B1(new_n551), .B2(new_n388), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G99gat), .B(G106gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n559), .A2(new_n541), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT41), .ZN(new_n564));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n564), .ZN(new_n567));
  NAND3_X1  g366(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n561), .A2(new_n567), .A3(new_n568), .A4(new_n562), .ZN(new_n569));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT102), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(new_n566), .B2(new_n569), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n521), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(new_n520), .A3(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n518), .A2(new_n579), .ZN(new_n580));
  OR3_X1    g379(.A1(new_n541), .A2(new_n501), .A3(KEYINPUT95), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT95), .B1(new_n541), .B2(new_n501), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n542), .A2(new_n501), .A3(new_n560), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT96), .ZN(new_n587));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT18), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n588), .A3(new_n584), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n541), .A2(new_n501), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n588), .B(KEYINPUT13), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n590), .A2(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT96), .B1(new_n590), .B2(new_n591), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n589), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G169gat), .B(G197gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n589), .A2(new_n596), .A3(new_n597), .A4(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT106), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT105), .ZN(new_n611));
  INV_X1    g410(.A(new_n485), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n557), .A2(new_n612), .A3(new_n558), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n553), .A2(new_n555), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n485), .B1(new_n614), .B2(new_n556), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n611), .B1(new_n616), .B2(KEYINPUT10), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT10), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n613), .A2(new_n615), .A3(KEYINPUT105), .A4(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n610), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n610), .A3(new_n622), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n316), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(G204gat), .Z(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n621), .A2(new_n622), .ZN(new_n633));
  INV_X1    g432(.A(new_n631), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n626), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n609), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n469), .A2(new_n580), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n457), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  INV_X1    g440(.A(new_n453), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n639), .B(new_n642), .C1(KEYINPUT16), .C2(G8gat), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n645));
  OR3_X1    g444(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT42), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n497), .B1(new_n639), .B2(new_n642), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n644), .B2(KEYINPUT42), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n645), .B1(new_n644), .B2(KEYINPUT42), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(G1325gat));
  AOI21_X1  g449(.A(G15gat), .B1(new_n639), .B2(new_n448), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n452), .A2(G15gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT108), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n639), .B2(new_n653), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n248), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n412), .A2(new_n460), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n463), .A2(new_n468), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n579), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n517), .A3(new_n637), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n661), .A2(G29gat), .A3(new_n458), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT45), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n517), .B(KEYINPUT109), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n637), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT110), .Z(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(KEYINPUT111), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n667), .A2(KEYINPUT111), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n660), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n668), .B1(new_n469), .B2(new_n579), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n666), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674), .B2(new_n458), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n663), .A2(new_n675), .ZN(G1328gat));
  NOR3_X1   g475(.A1(new_n661), .A2(G36gat), .A3(new_n453), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT46), .ZN(new_n678));
  OAI21_X1  g477(.A(G36gat), .B1(new_n674), .B2(new_n453), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1329gat));
  NAND2_X1  g479(.A1(new_n673), .A2(new_n452), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n536), .ZN(new_n682));
  OR2_X1    g481(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n683));
  INV_X1    g482(.A(new_n448), .ZN(new_n684));
  OR3_X1    g483(.A1(new_n661), .A2(new_n536), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1330gat));
  NOR3_X1   g487(.A1(new_n661), .A2(G50gat), .A3(new_n249), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n248), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(G50gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(KEYINPUT113), .A2(KEYINPUT48), .ZN(new_n692));
  OR2_X1    g491(.A1(KEYINPUT113), .A2(KEYINPUT48), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(G1331gat));
  NOR2_X1   g495(.A1(new_n580), .A2(new_n608), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n457), .B1(new_n394), .B2(new_n390), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n451), .B(new_n450), .C1(new_n698), .C2(new_n249), .ZN(new_n699));
  INV_X1    g498(.A(new_n393), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n397), .A2(new_n409), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n389), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n702), .B2(KEYINPUT38), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT38), .B1(new_n397), .B2(new_n398), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n467), .B1(new_n704), .B2(new_n389), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n248), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n699), .B1(new_n706), .B2(new_n395), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n463), .A2(new_n468), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n636), .B(new_n697), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(KEYINPUT114), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(KEYINPUT114), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n458), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n477), .ZN(G1332gat));
  NAND2_X1  g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n710), .A2(new_n642), .A3(new_n711), .A4(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT115), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(KEYINPUT115), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(G1333gat));
  INV_X1    g521(.A(new_n712), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(G71gat), .A3(new_n452), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n712), .A2(new_n684), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(G71gat), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT50), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n724), .B(new_n728), .C1(G71gat), .C2(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1334gat));
  NAND2_X1  g529(.A1(new_n723), .A2(new_n248), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  INV_X1    g531(.A(new_n579), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n518), .A2(new_n608), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n733), .B(new_n734), .C1(new_n707), .C2(new_n708), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT51), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n660), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n736), .A2(new_n636), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n457), .ZN(new_n740));
  INV_X1    g539(.A(new_n734), .ZN(new_n741));
  INV_X1    g540(.A(new_n636), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n671), .B2(new_n672), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(G85gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n740), .B1(new_n457), .B2(new_n746), .ZN(G1336gat));
  NOR2_X1   g546(.A1(new_n453), .A2(G92gat), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n736), .A2(new_n636), .A3(new_n738), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT118), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n453), .B(new_n744), .C1(new_n671), .C2(new_n672), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n388), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n749), .B2(KEYINPUT118), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT119), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AND4_X1   g554(.A1(new_n636), .A2(new_n736), .A3(new_n738), .A4(new_n748), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT52), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT119), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n671), .A2(new_n672), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n642), .A3(new_n743), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n758), .A2(new_n759), .A3(new_n762), .A4(new_n750), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT116), .B1(new_n751), .B2(new_n388), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT117), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n761), .A2(new_n767), .A3(G92gat), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n749), .A2(KEYINPUT117), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n765), .A2(new_n766), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n764), .A2(new_n771), .ZN(G1337gat));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n739), .A2(new_n773), .A3(new_n448), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n745), .A2(new_n452), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n773), .ZN(G1338gat));
  NAND2_X1  g575(.A1(new_n739), .A2(new_n248), .ZN(new_n777));
  INV_X1    g576(.A(G106gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n745), .A2(G106gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n249), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n779), .B(KEYINPUT53), .C1(new_n249), .C2(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1339gat));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n621), .A2(new_n610), .A3(new_n622), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n623), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n617), .A2(new_n625), .A3(new_n619), .A4(new_n620), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n633), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n631), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n631), .A4(new_n790), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n793), .A2(new_n608), .A3(new_n635), .A4(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n593), .B2(new_n595), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n585), .A2(G229gat), .A3(G233gat), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n583), .A2(KEYINPUT120), .A3(new_n592), .A4(new_n594), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n603), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n607), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n636), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n733), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n794), .A2(new_n635), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n802), .B1(new_n792), .B2(new_n791), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n733), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n664), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n697), .A2(new_n742), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n461), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n812), .A2(KEYINPUT121), .A3(new_n457), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT121), .B1(new_n812), .B2(new_n457), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n453), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n251), .A3(new_n608), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(new_n457), .A3(new_n453), .ZN(new_n818));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n609), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1340gat));
  OAI21_X1  g619(.A(G120gat), .B1(new_n818), .B2(new_n742), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n742), .A2(new_n253), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n815), .B2(new_n822), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n816), .B2(new_n518), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n818), .A2(new_n664), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(G127gat), .B2(new_n825), .ZN(G1342gat));
  NAND2_X1  g625(.A1(new_n816), .A2(new_n733), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n827), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n818), .B2(new_n579), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT56), .B1(new_n827), .B2(G134gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n453), .A2(new_n457), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n452), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n249), .B1(new_n809), .B2(new_n810), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n806), .A2(new_n807), .A3(new_n733), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n791), .A2(new_n792), .B1(new_n606), .B2(new_n607), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n806), .A2(new_n839), .B1(new_n636), .B2(new_n803), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n840), .B2(new_n733), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n841), .A2(new_n517), .B1(new_n742), .B2(new_n697), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT57), .B1(new_n842), .B2(new_n249), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n608), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(G141gat), .ZN(new_n845));
  INV_X1    g644(.A(new_n835), .ZN(new_n846));
  NOR4_X1   g645(.A1(new_n846), .A2(G141gat), .A3(new_n609), .A4(new_n834), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n845), .A2(KEYINPUT58), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n837), .A2(KEYINPUT122), .A3(new_n843), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT122), .B1(new_n837), .B2(new_n843), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n608), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n847), .B1(new_n851), .B2(G141gat), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT123), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n848), .B(new_n856), .C1(new_n852), .C2(new_n853), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1344gat));
  OAI21_X1  g657(.A(new_n636), .B1(new_n849), .B2(new_n850), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(G148gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT124), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n859), .A2(new_n863), .A3(new_n860), .A4(G148gat), .ZN(new_n864));
  INV_X1    g663(.A(G148gat), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n842), .A2(KEYINPUT57), .A3(new_n249), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n846), .A2(KEYINPUT57), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n742), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n869), .B2(new_n833), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n862), .B(new_n864), .C1(new_n860), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n846), .A2(new_n834), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n865), .A3(new_n636), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1345gat));
  AOI21_X1  g673(.A(G155gat), .B1(new_n872), .B2(new_n518), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n849), .A2(new_n850), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n664), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n872), .B2(new_n733), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n876), .A2(new_n579), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n453), .A2(new_n457), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n812), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n609), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(new_n315), .ZN(G1348gat));
  INV_X1    g684(.A(new_n883), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n636), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G176gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n317), .A2(new_n318), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(G1349gat));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n518), .A3(new_n297), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n300), .B1(new_n883), .B2(new_n664), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(KEYINPUT125), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n298), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n883), .B2(new_n579), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n886), .A2(new_n733), .B1(new_n897), .B2(new_n298), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n898), .ZN(G1351gat));
  NOR3_X1   g700(.A1(new_n452), .A2(new_n457), .A3(new_n453), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n846), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(G197gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n608), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n868), .A2(new_n609), .A3(new_n903), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n905), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n869), .A2(new_n902), .ZN(new_n909));
  XNOR2_X1  g708(.A(KEYINPUT126), .B(G204gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR4_X1   g710(.A1(new_n846), .A2(new_n742), .A3(new_n903), .A4(new_n910), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT62), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1353gat));
  NAND3_X1  g713(.A1(new_n904), .A2(new_n207), .A3(new_n518), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n866), .A2(new_n867), .A3(new_n518), .A4(new_n902), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n916), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT63), .B1(new_n916), .B2(G211gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT127), .ZN(G1354gat));
  AOI21_X1  g719(.A(G218gat), .B1(new_n904), .B2(new_n733), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n868), .A2(new_n903), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n579), .A2(new_n208), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1355gat));
endmodule


