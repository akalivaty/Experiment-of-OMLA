//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G43gat), .ZN(new_n205));
  INV_X1    g004(.A(G43gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(KEYINPUT90), .ZN(new_n214));
  OAI21_X1  g013(.A(G29gat), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT89), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n213), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT14), .A3(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(KEYINPUT14), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n210), .A2(new_n215), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT15), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT15), .B1(new_n205), .B2(new_n207), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n213), .A2(KEYINPUT90), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n211), .A2(G36gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n217), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n230), .A2(new_n223), .A3(new_n220), .A4(new_n221), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(G1gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT16), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G1gat), .B2(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G8gat), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n236), .B(new_n239), .C1(G1gat), .C2(new_n233), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n231), .A3(KEYINPUT17), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT91), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT91), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n225), .A2(new_n231), .A3(new_n245), .A4(KEYINPUT17), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT17), .B1(new_n225), .B2(new_n231), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(new_n241), .ZN(new_n249));
  AOI211_X1 g048(.A(new_n203), .B(new_n242), .C1(new_n247), .C2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT93), .B1(new_n232), .B2(new_n241), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n241), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n202), .B(KEYINPUT13), .Z(new_n254));
  AOI22_X1  g053(.A1(new_n250), .A2(KEYINPUT18), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT11), .B(G169gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT12), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n250), .B2(KEYINPUT18), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n261), .B(KEYINPUT88), .Z(new_n264));
  NAND2_X1  g063(.A1(new_n253), .A2(new_n254), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n242), .B1(new_n247), .B2(new_n249), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT18), .A3(new_n202), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT18), .B1(new_n266), .B2(new_n202), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n265), .B(new_n267), .C1(new_n268), .C2(KEYINPUT92), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT92), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n250), .A2(new_n270), .A3(KEYINPUT18), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n264), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT94), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n250), .B2(KEYINPUT18), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n266), .A2(new_n202), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT18), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT92), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n255), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(KEYINPUT94), .A3(new_n264), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n263), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G85gat), .A2(G92gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT98), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT97), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n284), .B(KEYINPUT7), .C1(KEYINPUT97), .C2(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(G99gat), .A2(G106gat), .ZN(new_n286));
  INV_X1    g085(.A(G85gat), .ZN(new_n287));
  INV_X1    g086(.A(G92gat), .ZN(new_n288));
  AOI22_X1  g087(.A1(KEYINPUT8), .A2(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n285), .B(new_n289), .C1(KEYINPUT7), .C2(new_n284), .ZN(new_n290));
  XOR2_X1   g089(.A(G99gat), .B(G106gat), .Z(new_n291));
  OR2_X1    g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n291), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(new_n248), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n247), .ZN(new_n297));
  AND2_X1   g096(.A1(G232gat), .A2(G233gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n295), .A2(new_n232), .B1(KEYINPUT41), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G190gat), .B(G218gat), .Z(new_n301));
  AND2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n300), .A2(new_n301), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n298), .A2(KEYINPUT41), .ZN(new_n304));
  XNOR2_X1  g103(.A(G134gat), .B(G162gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OR3_X1    g106(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n302), .B2(new_n303), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G71gat), .A2(G78gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(G71gat), .A2(G78gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G57gat), .B(G64gat), .Z(new_n314));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(KEYINPUT9), .B2(new_n311), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT99), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n290), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n294), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n292), .A2(new_n318), .A3(new_n293), .A4(new_n320), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n295), .A2(KEYINPUT10), .A3(new_n318), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G230gat), .ZN(new_n328));
  INV_X1    g127(.A(G233gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n322), .B2(new_n324), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n333), .A2(KEYINPUT100), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(KEYINPUT100), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G120gat), .B(G148gat), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT101), .ZN(new_n338));
  XNOR2_X1  g137(.A(G176gat), .B(G204gat), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n338), .B(new_n339), .Z(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n332), .A2(new_n334), .A3(new_n340), .A4(new_n335), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n318), .A2(KEYINPUT21), .ZN(new_n346));
  XNOR2_X1  g145(.A(G127gat), .B(G155gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n346), .B(new_n347), .Z(new_n348));
  AOI21_X1  g147(.A(new_n241), .B1(new_n318), .B2(KEYINPUT21), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  NAND2_X1  g150(.A1(G231gat), .A2(G233gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT96), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G183gat), .B(G211gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n350), .A2(new_n351), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n357), .B1(new_n350), .B2(new_n351), .ZN(new_n359));
  OR2_X1    g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n310), .A2(new_n345), .A3(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n361), .B(KEYINPUT102), .Z(new_n362));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT35), .ZN(new_n364));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n366));
  INV_X1    g165(.A(G211gat), .ZN(new_n367));
  INV_X1    g166(.A(G218gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  XOR2_X1   g169(.A(G211gat), .B(G218gat), .Z(new_n371));
  OAI21_X1  g170(.A(KEYINPUT78), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT78), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(KEYINPUT77), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n371), .B1(new_n370), .B2(KEYINPUT77), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n373), .A2(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT3), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G141gat), .B(G148gat), .Z(new_n381));
  INV_X1    g180(.A(G155gat), .ZN(new_n382));
  INV_X1    g181(.A(G162gat), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT2), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G155gat), .B(G162gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(new_n386), .A3(new_n384), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT82), .B1(new_n380), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n395), .A3(new_n389), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n379), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n398), .B2(new_n378), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n370), .A2(KEYINPUT77), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n371), .A3(new_n375), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n365), .A2(new_n369), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT78), .ZN(new_n405));
  INV_X1    g204(.A(new_n371), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n372), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT29), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n401), .B(new_n390), .C1(new_n409), .C2(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n400), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT83), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n400), .A2(new_n392), .A3(new_n413), .A4(new_n410), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n398), .A2(new_n378), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n407), .A2(KEYINPUT80), .A3(new_n372), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n370), .A2(new_n371), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT80), .B1(new_n407), .B2(new_n372), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n379), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n391), .B1(new_n422), .B2(new_n395), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n417), .B1(new_n423), .B2(KEYINPUT81), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425));
  AOI211_X1 g224(.A(new_n425), .B(new_n391), .C1(new_n422), .C2(new_n395), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n393), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G22gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n415), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT84), .ZN(new_n430));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT31), .B(G50gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n427), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G22gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n429), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n430), .A2(new_n436), .A3(new_n429), .A4(new_n433), .ZN(new_n439));
  XOR2_X1   g238(.A(G127gat), .B(G134gat), .Z(new_n440));
  XNOR2_X1  g239(.A(G113gat), .B(G120gat), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(KEYINPUT1), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n440), .A2(KEYINPUT1), .ZN(new_n444));
  INV_X1    g243(.A(G113gat), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n445), .A2(G120gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT71), .B(G120gat), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(G113gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT72), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n449), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n443), .B(new_n444), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n448), .B(new_n449), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n443), .B1(new_n454), .B2(new_n444), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n442), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(G183gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT27), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT27), .ZN(new_n460));
  AOI21_X1  g259(.A(G190gat), .B1(new_n460), .B2(G183gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n457), .A3(KEYINPUT27), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT28), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n459), .A2(new_n461), .A3(new_n463), .A4(KEYINPUT69), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n460), .A2(G183gat), .ZN(new_n470));
  INV_X1    g269(.A(G190gat), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n458), .A2(new_n470), .A3(KEYINPUT28), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(G169gat), .A2(G176gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT26), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT70), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G169gat), .A2(G176gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n474), .A2(KEYINPUT70), .A3(new_n475), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n474), .A2(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n474), .A2(KEYINPUT66), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n475), .A3(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n480), .A2(new_n483), .B1(G183gat), .B2(G190gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT25), .ZN(new_n485));
  NOR2_X1   g284(.A1(G183gat), .A2(G190gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT65), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n457), .A2(KEYINPUT24), .ZN(new_n489));
  NAND2_X1  g288(.A1(G183gat), .A2(G190gat), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n489), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n474), .B1(KEYINPUT23), .B2(new_n477), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n474), .A2(KEYINPUT23), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n485), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT23), .A3(new_n482), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n493), .A2(new_n485), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n486), .B(KEYINPUT67), .Z(new_n499));
  OAI211_X1 g298(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n491), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n473), .A2(new_n484), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n456), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT64), .ZN(new_n504));
  INV_X1    g303(.A(new_n442), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n444), .B1(new_n450), .B2(new_n451), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n507), .B2(new_n452), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n473), .A2(new_n484), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n496), .A2(new_n500), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT32), .ZN(new_n514));
  XOR2_X1   g313(.A(G15gat), .B(G43gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT75), .ZN(new_n516));
  XNOR2_X1  g315(.A(G71gat), .B(G99gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT74), .B1(new_n513), .B2(new_n519), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n514), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT34), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n502), .A2(new_n512), .ZN(new_n525));
  INV_X1    g324(.A(new_n504), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI211_X1 g326(.A(KEYINPUT34), .B(new_n504), .C1(new_n502), .C2(new_n512), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n514), .B1(KEYINPUT33), .B2(new_n518), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n523), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n534));
  INV_X1    g333(.A(new_n522), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n520), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n533), .B1(new_n536), .B2(new_n530), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n438), .A2(new_n439), .A3(new_n532), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n511), .A2(G226gat), .A3(G233gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(G226gat), .A2(G233gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n501), .B2(KEYINPUT29), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n378), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n541), .A3(new_n378), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G8gat), .B(G36gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(G64gat), .B(G92gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n544), .A2(new_n549), .A3(new_n545), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT30), .A3(new_n552), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n546), .A2(KEYINPUT30), .A3(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n508), .A2(new_n556), .A3(new_n391), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n442), .B(new_n391), .C1(new_n453), .C2(new_n455), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n396), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n508), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n557), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT5), .ZN(new_n564));
  NAND2_X1  g363(.A1(G225gat), .A2(G233gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G1gat), .B(G29gat), .Z(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G57gat), .B(G85gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n565), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n558), .B(KEYINPUT4), .C1(new_n508), .C2(new_n561), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n557), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n508), .A2(new_n391), .ZN(new_n576));
  AOI211_X1 g375(.A(new_n505), .B(new_n390), .C1(new_n507), .C2(new_n452), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT5), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n566), .B(new_n572), .C1(new_n575), .C2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n565), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(KEYINPUT5), .A3(new_n578), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n572), .B1(new_n584), .B2(new_n566), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n579), .A2(new_n575), .ZN(new_n587));
  AOI211_X1 g386(.A(KEYINPUT5), .B(new_n573), .C1(new_n574), .C2(new_n557), .ZN(new_n588));
  OAI211_X1 g387(.A(KEYINPUT6), .B(new_n571), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n555), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n364), .B1(new_n538), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n433), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n429), .B2(KEYINPUT84), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n437), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n537), .A2(new_n532), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n555), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n571), .B1(new_n587), .B2(new_n588), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(new_n581), .A3(new_n580), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n598), .B1(new_n600), .B2(new_n589), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n595), .A2(new_n597), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n592), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT76), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT36), .B1(new_n596), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607));
  AOI211_X1 g406(.A(KEYINPUT76), .B(new_n607), .C1(new_n537), .C2(new_n532), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n574), .A2(new_n573), .A3(new_n557), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n610), .A2(KEYINPUT39), .ZN(new_n611));
  OR3_X1    g410(.A1(new_n576), .A2(new_n577), .A3(new_n573), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT39), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n572), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n611), .A2(KEYINPUT40), .A3(new_n613), .A4(new_n572), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n598), .A2(new_n599), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT86), .ZN(new_n619));
  INV_X1    g418(.A(new_n545), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n378), .B1(new_n539), .B2(new_n541), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT37), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n550), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT85), .B1(new_n546), .B2(KEYINPUT37), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT85), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT37), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n544), .A2(new_n625), .A3(new_n626), .A4(new_n545), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n619), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n627), .ZN(new_n631));
  INV_X1    g430(.A(new_n623), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(KEYINPUT86), .A3(KEYINPUT38), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n632), .A3(new_n629), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n600), .A2(new_n589), .A3(new_n552), .A4(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n595), .B(new_n618), .C1(new_n635), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n438), .A2(new_n439), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n591), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n609), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  AOI211_X1 g440(.A(new_n281), .B(new_n362), .C1(new_n604), .C2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n586), .A2(new_n590), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n598), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n239), .B1(new_n642), .B2(new_n598), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n647), .B1(new_n653), .B2(new_n648), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n651), .B1(new_n652), .B2(new_n654), .ZN(G1325gat));
  INV_X1    g454(.A(G15gat), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n642), .A2(new_n656), .A3(new_n597), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n596), .A2(new_n605), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n607), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n596), .A2(new_n605), .A3(KEYINPUT36), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n642), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n662), .B2(new_n656), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n642), .A2(new_n639), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT104), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT43), .B(G22gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  INV_X1    g466(.A(new_n310), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n609), .A2(new_n638), .A3(new_n640), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n592), .A2(new_n603), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT44), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n310), .B1(new_n604), .B2(new_n641), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT105), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n640), .A2(KEYINPUT106), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n591), .A2(new_n678), .A3(new_n639), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n677), .A2(new_n609), .A3(new_n638), .A4(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n310), .B1(new_n680), .B2(new_n604), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n675), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n673), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n281), .A2(new_n360), .A3(new_n344), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n643), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n674), .A2(new_n684), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n217), .A3(new_n643), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(G1328gat));
  NAND4_X1  g490(.A1(new_n688), .A2(new_n598), .A3(new_n227), .A4(new_n228), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT107), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  OAI22_X1  g495(.A1(new_n685), .A2(new_n555), .B1(new_n212), .B2(new_n214), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(G1329gat));
  OAI21_X1  g497(.A(G43gat), .B1(new_n685), .B2(new_n609), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n688), .A2(new_n206), .A3(new_n597), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1330gat));
  AND3_X1   g502(.A1(new_n688), .A2(new_n204), .A3(new_n639), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n683), .A2(new_n639), .A3(new_n684), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(G50gat), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n705), .B2(G50gat), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI221_X4 g509(.A(new_n704), .B1(new_n707), .B2(KEYINPUT48), .C1(new_n705), .C2(G50gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(G1331gat));
  NAND3_X1  g511(.A1(new_n281), .A2(new_n360), .A3(new_n310), .ZN(new_n713));
  AOI211_X1 g512(.A(new_n345), .B(new_n713), .C1(new_n680), .C2(new_n604), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n643), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT109), .B(G57gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1332gat));
  AOI21_X1  g516(.A(new_n555), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT110), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n720), .B(new_n721), .Z(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n714), .A2(new_n723), .A3(new_n597), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n714), .A2(new_n661), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n639), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT111), .B(G78gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1335gat));
  INV_X1    g529(.A(new_n360), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n281), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n681), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT51), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n681), .A2(KEYINPUT51), .A3(new_n733), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT114), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n736), .A2(KEYINPUT114), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n643), .A2(new_n287), .A3(new_n344), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT115), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n733), .A2(new_n344), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n683), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT113), .B1(new_n745), .B2(new_n686), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G85gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n745), .A2(KEYINPUT113), .A3(new_n686), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n742), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  NOR3_X1   g548(.A1(new_n345), .A2(new_n555), .A3(G92gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n683), .A2(new_n598), .A3(new_n744), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n753), .A2(new_n756), .A3(G92gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n753), .B2(G92gat), .ZN(new_n758));
  INV_X1    g557(.A(new_n750), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n735), .B2(new_n736), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n755), .B1(new_n761), .B2(new_n752), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n596), .A2(G99gat), .A3(new_n345), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n739), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G99gat), .B1(new_n745), .B2(new_n609), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1338gat));
  NOR3_X1   g565(.A1(new_n595), .A2(G106gat), .A3(new_n345), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n739), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n683), .A2(new_n639), .A3(new_n744), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n767), .B(KEYINPUT117), .Z(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n735), .B2(new_n736), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n769), .B2(G106gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(G1339gat));
  NOR2_X1   g576(.A1(new_n713), .A2(new_n344), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n325), .A2(new_n330), .A3(new_n326), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n332), .A2(new_n779), .A3(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n330), .B1(new_n325), .B2(new_n326), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n340), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n780), .A2(KEYINPUT55), .A3(new_n783), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n786), .A2(new_n343), .A3(new_n787), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n253), .A2(new_n254), .B1(new_n266), .B2(new_n202), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n263), .B1(new_n260), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n668), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n263), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n279), .A2(KEYINPUT94), .A3(new_n264), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT94), .B1(new_n279), .B2(new_n264), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n795), .A2(new_n788), .B1(new_n344), .B2(new_n790), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n796), .B2(new_n668), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n778), .B1(new_n797), .B2(new_n731), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n639), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(new_n643), .A3(new_n555), .A4(new_n597), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n445), .A3(new_n281), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n713), .A2(new_n344), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n789), .A2(new_n260), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n792), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n343), .A3(new_n787), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n804), .A2(new_n805), .A3(new_n310), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n344), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n281), .B2(new_n805), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n808), .B2(new_n310), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n802), .B1(new_n809), .B2(new_n360), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n643), .A3(new_n595), .A4(new_n597), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n598), .ZN(new_n812));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n795), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n801), .A2(new_n813), .ZN(G1340gat));
  OAI21_X1  g613(.A(G120gat), .B1(new_n800), .B2(new_n345), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n447), .A3(new_n344), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1341gat));
  OAI21_X1  g616(.A(G127gat), .B1(new_n800), .B2(new_n731), .ZN(new_n818));
  INV_X1    g617(.A(G127gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n812), .A2(new_n819), .A3(new_n360), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1342gat));
  NAND2_X1  g620(.A1(new_n668), .A2(new_n555), .ZN(new_n822));
  OR3_X1    g621(.A1(new_n811), .A2(G134gat), .A3(new_n822), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n824));
  OAI21_X1  g623(.A(G134gat), .B1(new_n800), .B2(new_n310), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n661), .A2(new_n595), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n810), .A2(new_n829), .A3(new_n643), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT120), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n281), .A2(G141gat), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n810), .A2(new_n829), .A3(new_n833), .A4(new_n643), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n831), .A2(new_n555), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n609), .A2(new_n643), .A3(new_n555), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n837), .B1(new_n798), .B2(new_n595), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n810), .A2(KEYINPUT57), .A3(new_n639), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n281), .B(new_n836), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(G141gat), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n828), .B(new_n835), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n836), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n798), .A2(new_n837), .A3(new_n595), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n810), .B2(new_n639), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n795), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n849), .A2(KEYINPUT121), .A3(new_n828), .A4(new_n835), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  INV_X1    g651(.A(new_n832), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n830), .A2(new_n598), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n848), .B2(G141gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n828), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n841), .B1(new_n857), .B2(new_n795), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT119), .B(KEYINPUT58), .C1(new_n858), .C2(new_n854), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n851), .A2(new_n860), .A3(KEYINPUT122), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n831), .A2(new_n834), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n598), .ZN(new_n867));
  INV_X1    g666(.A(G148gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n344), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n362), .A2(new_n795), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n731), .B2(new_n797), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n837), .B1(new_n872), .B2(new_n595), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n839), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n344), .A3(new_n845), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n870), .B1(new_n875), .B2(G148gat), .ZN(new_n876));
  AOI211_X1 g675(.A(KEYINPUT59), .B(new_n868), .C1(new_n857), .C2(new_n344), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n869), .B1(new_n876), .B2(new_n877), .ZN(G1345gat));
  NAND3_X1  g677(.A1(new_n867), .A2(new_n382), .A3(new_n360), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n857), .A2(new_n360), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n382), .B2(new_n880), .ZN(G1346gat));
  NOR3_X1   g680(.A1(new_n866), .A2(G162gat), .A3(new_n822), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n383), .B1(new_n857), .B2(new_n668), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT123), .Z(G1347gat));
  NOR4_X1   g684(.A1(new_n798), .A2(new_n643), .A3(new_n555), .A4(new_n538), .ZN(new_n886));
  AOI21_X1  g685(.A(G169gat), .B1(new_n886), .B2(new_n795), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n643), .A2(new_n555), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n799), .A2(new_n597), .A3(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n795), .A2(G169gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(G1348gat));
  OAI21_X1  g693(.A(G176gat), .B1(new_n891), .B2(new_n345), .ZN(new_n895));
  INV_X1    g694(.A(G176gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n886), .A2(new_n896), .A3(new_n344), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1349gat));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(KEYINPUT60), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(KEYINPUT60), .ZN(new_n901));
  OAI21_X1  g700(.A(G183gat), .B1(new_n891), .B2(new_n731), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n458), .A3(new_n470), .A4(new_n360), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n900), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  AND4_X1   g703(.A1(new_n899), .A2(new_n902), .A3(KEYINPUT60), .A4(new_n903), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1350gat));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n471), .A3(new_n668), .ZN(new_n907));
  OAI21_X1  g706(.A(G190gat), .B1(new_n891), .B2(new_n310), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(KEYINPUT61), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(KEYINPUT61), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(G1351gat));
  NOR2_X1   g710(.A1(new_n798), .A2(new_n643), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n661), .A2(new_n555), .A3(new_n595), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n795), .ZN(new_n916));
  INV_X1    g715(.A(new_n874), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n609), .A2(new_n888), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT126), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n795), .A2(G197gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(G1352gat));
  NOR3_X1   g722(.A1(new_n914), .A2(G204gat), .A3(new_n345), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT62), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n917), .A2(new_n345), .A3(new_n920), .ZN(new_n926));
  INV_X1    g725(.A(G204gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n915), .A2(new_n367), .A3(new_n360), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n874), .A2(new_n609), .A3(new_n360), .A4(new_n888), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  NAND4_X1  g732(.A1(new_n874), .A2(G218gat), .A3(new_n668), .A4(new_n919), .ZN(new_n934));
  AOI21_X1  g733(.A(G218gat), .B1(new_n915), .B2(new_n668), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


