//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1199, new_n1200, new_n1201,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n208), .B1(G68), .B2(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n203), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NOR2_X1   g0026(.A1(G58), .A2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n223), .A2(new_n226), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n220), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  INV_X1    g0039(.A(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT64), .Z(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G169), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(G238), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G226), .A2(G1698), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(new_n220), .B2(G1698), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n260), .A2(new_n261), .B1(G33), .B2(G97), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n256), .B(new_n258), .C1(new_n262), .C2(new_n253), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n251), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT14), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT72), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  OR3_X1    g0069(.A1(new_n263), .A2(new_n268), .A3(KEYINPUT13), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT74), .B1(new_n271), .B2(G179), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT74), .ZN(new_n273));
  INV_X1    g0073(.A(G179), .ZN(new_n274));
  AOI211_X1 g0074(.A(new_n273), .B(new_n274), .C1(new_n269), .C2(new_n270), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n267), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n254), .A2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(G13), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(KEYINPUT12), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(KEYINPUT69), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n231), .B1(new_n203), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(new_n277), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT12), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n280), .B1(new_n287), .B2(G68), .ZN(new_n288));
  INV_X1    g0088(.A(G68), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n281), .A2(KEYINPUT12), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n283), .A2(G20), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n291), .A2(G77), .B1(G20), .B2(new_n289), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n214), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n284), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n297), .A2(KEYINPUT11), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT11), .B1(new_n297), .B2(new_n298), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n288), .B(new_n290), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n276), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(G190), .B2(new_n271), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n264), .B2(new_n265), .ZN(new_n305));
  XOR2_X1   g0105(.A(new_n305), .B(KEYINPUT71), .Z(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G222), .ZN(new_n310));
  INV_X1    g0110(.A(G223), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n261), .B(new_n310), .C1(new_n311), .C2(new_n309), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(new_n252), .C1(G77), .C2(new_n261), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n253), .A2(new_n255), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n258), .C1(new_n215), .C2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(new_n315), .B(KEYINPUT65), .Z(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G200), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n315), .B(KEYINPUT65), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G190), .ZN(new_n319));
  INV_X1    g0119(.A(new_n277), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n320), .A2(KEYINPUT66), .A3(new_n214), .ZN(new_n321));
  INV_X1    g0121(.A(new_n279), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT66), .B1(new_n320), .B2(new_n214), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n285), .A4(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n294), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n291), .B2(new_n329), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n324), .B1(G50), .B2(new_n322), .C1(new_n330), .C2(new_n285), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT9), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n317), .A2(new_n319), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT10), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n318), .A2(new_n274), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n331), .C1(G169), .C2(new_n318), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n286), .A2(new_n216), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n328), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n293), .ZN(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT15), .B(G87), .Z(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n285), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n282), .A2(G77), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n337), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G238), .A2(G1698), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n220), .B2(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n261), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n210), .B2(new_n261), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(KEYINPUT67), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(KEYINPUT67), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n252), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n253), .A2(G244), .A3(new_n255), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n353), .A2(new_n258), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(KEYINPUT70), .A3(new_n274), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n355), .B2(G179), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n345), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n251), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n308), .A2(new_n334), .A3(new_n336), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n261), .B2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G33), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT7), .A3(new_n230), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G68), .ZN(new_n372));
  AND2_X1   g0172(.A1(G58), .A2(G68), .ZN(new_n373));
  OAI21_X1  g0173(.A(G20), .B1(new_n373), .B2(new_n227), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT76), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n293), .A2(G159), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT76), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(G20), .C1(new_n373), .C2(new_n227), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT16), .B1(new_n372), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n285), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n367), .A2(KEYINPUT75), .A3(G33), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT75), .B1(new_n367), .B2(G33), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n366), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n364), .A3(new_n230), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n367), .A2(G33), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT75), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n283), .B2(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n367), .A2(KEYINPUT75), .A3(G33), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT7), .B1(new_n393), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(new_n394), .A3(G68), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n380), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n289), .B1(new_n365), .B2(new_n370), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n379), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT77), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n383), .A2(new_n384), .A3(new_n396), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n396), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n284), .B1(new_n399), .B2(KEYINPUT77), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT78), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n322), .B1(new_n328), .B2(new_n284), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n277), .B2(new_n328), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT79), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n401), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n311), .A2(new_n309), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n393), .B(new_n409), .C1(G226), .C2(new_n309), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n253), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n258), .B1(new_n314), .B2(new_n220), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT80), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT80), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n258), .C1(new_n314), .C2(new_n220), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n412), .A2(new_n413), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n274), .A2(new_n417), .B1(new_n418), .B2(new_n251), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n408), .A2(KEYINPUT18), .A3(new_n419), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n418), .A2(new_n304), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n401), .A2(new_n404), .A3(new_n428), .A4(new_n407), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n345), .B1(new_n355), .B2(new_n425), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n356), .A2(new_n304), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n363), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT89), .ZN(new_n437));
  INV_X1    g0237(.A(G45), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(G1), .ZN(new_n439));
  AND2_X1   g0239(.A1(KEYINPUT5), .A2(G41), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n253), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n211), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n205), .A2(new_n309), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n207), .A2(G1698), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n393), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G294), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n437), .B(new_n445), .C1(new_n450), .C2(new_n253), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n442), .A2(new_n257), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n253), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT89), .B1(new_n453), .B2(new_n444), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n304), .ZN(new_n456));
  INV_X1    g0256(.A(new_n452), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n453), .A2(new_n444), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n425), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n283), .A2(G1), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n279), .A2(new_n284), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G107), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n393), .A2(KEYINPUT22), .A3(G87), .ZN(new_n465));
  NAND2_X1  g0265(.A1(G33), .A2(G116), .ZN(new_n466));
  AOI21_X1  g0266(.A(G20), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n369), .A2(G20), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT22), .B1(new_n468), .B2(G87), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n210), .A2(G20), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n471), .B(KEYINPUT23), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n464), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NOR4_X1   g0274(.A1(new_n467), .A2(KEYINPUT24), .A3(new_n469), .A4(new_n472), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n284), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n279), .A2(new_n210), .ZN(new_n477));
  XOR2_X1   g0277(.A(new_n477), .B(KEYINPUT25), .Z(new_n478));
  NAND4_X1  g0278(.A1(new_n460), .A2(new_n463), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(new_n463), .A3(new_n478), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n455), .A2(new_n274), .B1(new_n251), .B2(new_n458), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n443), .A2(new_n240), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n207), .A2(new_n309), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n393), .B(new_n486), .C1(G264), .C2(new_n309), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n369), .A2(G303), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n452), .B(new_n485), .C1(new_n489), .C2(new_n253), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT86), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n253), .B1(new_n487), .B2(new_n488), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(new_n484), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n494), .A3(new_n452), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(G200), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n230), .C1(G33), .C2(new_n206), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G20), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n498), .A2(new_n284), .A3(KEYINPUT20), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n284), .A3(new_n500), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n506), .A2(KEYINPUT88), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(KEYINPUT88), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n281), .A2(new_n499), .ZN(new_n510));
  INV_X1    g0310(.A(new_n461), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n282), .A2(G116), .A3(new_n285), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n494), .B1(new_n493), .B2(new_n452), .ZN(new_n515));
  NOR4_X1   g0315(.A1(new_n492), .A2(new_n457), .A3(KEYINPUT86), .A4(new_n484), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n496), .B(new_n514), .C1(new_n517), .C2(new_n425), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n517), .A2(KEYINPUT21), .A3(G169), .A4(new_n513), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n490), .A2(new_n274), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n491), .A2(new_n513), .A3(new_n495), .A4(G169), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT21), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n518), .A2(new_n519), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n497), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n217), .A2(G1698), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n393), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n369), .A2(new_n205), .A3(new_n309), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n528), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT82), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n531), .A2(new_n533), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n252), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n253), .A2(new_n442), .A3(G257), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n452), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n541), .B(KEYINPUT83), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n538), .B2(new_n252), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n543), .A2(G200), .B1(new_n544), .B2(G190), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n322), .A2(G97), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n462), .A2(G97), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n371), .A2(G107), .B1(G77), .B2(new_n293), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT81), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT6), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n210), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n556), .A2(G107), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n548), .B1(new_n558), .B2(new_n230), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n546), .B(new_n547), .C1(new_n559), .C2(new_n284), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n545), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n284), .ZN(new_n562));
  INV_X1    g0362(.A(new_n546), .ZN(new_n563));
  INV_X1    g0363(.A(new_n547), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n539), .A2(new_n542), .A3(new_n274), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n527), .B(new_n532), .C1(new_n530), .C2(new_n529), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n537), .A2(new_n536), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n253), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n251), .B1(new_n569), .B2(new_n541), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n561), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n393), .A2(new_n230), .A3(G68), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G97), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n230), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT84), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n204), .A2(new_n206), .A3(new_n210), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(new_n230), .C1(new_n574), .C2(new_n575), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n291), .A2(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n575), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n573), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n341), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n284), .B1(new_n281), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G250), .B1(new_n438), .B2(G1), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n439), .A2(G274), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n252), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G238), .A2(G1698), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n217), .B2(G1698), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n393), .A2(new_n592), .B1(G33), .B2(G116), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n590), .B1(new_n593), .B2(new_n253), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n462), .A2(G87), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n586), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(G190), .B(new_n590), .C1(new_n593), .C2(new_n253), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT85), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n462), .A2(new_n341), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n586), .A2(new_n602), .B1(new_n251), .B2(new_n594), .ZN(new_n603));
  INV_X1    g0403(.A(new_n594), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n274), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n572), .A2(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n436), .A2(new_n483), .A3(new_n526), .A4(new_n608), .ZN(G372));
  NAND4_X1  g0409(.A1(new_n586), .A2(new_n595), .A3(new_n596), .A4(new_n598), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n455), .A2(new_n304), .B1(new_n425), .B2(new_n458), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n480), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT90), .B1(new_n614), .B2(new_n572), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n547), .B1(new_n559), .B2(new_n284), .ZN(new_n616));
  INV_X1    g0416(.A(new_n541), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n539), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n616), .A2(new_n563), .B1(new_n618), .B2(new_n251), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(new_n566), .B1(new_n545), .B2(new_n560), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT90), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(new_n479), .A3(new_n621), .A4(new_n612), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n482), .A2(new_n521), .A3(new_n519), .A4(new_n524), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n615), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n606), .B(KEYINPUT91), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n612), .A2(new_n627), .A3(new_n566), .A4(new_n619), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT26), .B1(new_n571), .B2(new_n607), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n436), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g0432(.A(new_n632), .B(KEYINPUT92), .Z(new_n633));
  INV_X1    g0433(.A(new_n362), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n307), .B1(new_n301), .B2(new_n276), .ZN(new_n635));
  INV_X1    g0435(.A(new_n430), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n424), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n334), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n638), .A2(new_n336), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(new_n639), .ZN(G369));
  NAND3_X1  g0440(.A1(new_n519), .A2(new_n524), .A3(new_n521), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n278), .A2(G20), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n254), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n514), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n525), .B2(new_n650), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G330), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n480), .A2(new_n648), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n480), .A2(new_n481), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n483), .A2(new_n655), .B1(new_n656), .B2(new_n648), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n641), .A2(new_n649), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n658), .A2(new_n483), .B1(new_n656), .B2(new_n649), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n224), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n578), .A2(G116), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n229), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n526), .A2(new_n483), .A3(new_n608), .A4(new_n649), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n451), .A2(new_n454), .A3(new_n604), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT93), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT93), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n451), .A2(new_n454), .A3(new_n674), .A4(new_n604), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n520), .A3(new_n544), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n675), .A2(new_n544), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(KEYINPUT30), .A3(new_n520), .A4(new_n673), .ZN(new_n680));
  AOI21_X1  g0480(.A(G179), .B1(new_n539), .B2(new_n542), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n517), .A2(new_n455), .A3(new_n594), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n671), .A2(KEYINPUT31), .B1(new_n648), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n683), .A2(KEYINPUT94), .A3(KEYINPUT31), .A4(new_n648), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(G330), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n597), .A2(new_n600), .B1(new_n603), .B2(new_n605), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n619), .A2(new_n693), .A3(new_n627), .A4(new_n566), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n571), .B2(new_n611), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n626), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT95), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n623), .A2(new_n479), .A3(new_n620), .A4(new_n612), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT95), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n626), .A2(new_n695), .A3(new_n699), .A4(new_n694), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n692), .B1(new_n701), .B2(new_n649), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n631), .A2(new_n649), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  OR4_X1    g0504(.A1(KEYINPUT96), .A2(new_n691), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n704), .A2(new_n702), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT96), .B1(new_n706), .B2(new_n691), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n670), .B1(new_n708), .B2(G1), .ZN(G364));
  NAND2_X1  g0509(.A1(new_n642), .A2(G45), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n666), .A2(G1), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT97), .Z(new_n712));
  NOR2_X1   g0512(.A1(new_n654), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(G330), .B2(new_n652), .ZN(new_n714));
  OAI211_X1 g0514(.A(G1), .B(G13), .C1(new_n230), .C2(G169), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT98), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(KEYINPUT98), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n230), .A2(new_n425), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n274), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G322), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n304), .A2(G179), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n230), .A2(G190), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G283), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n274), .A2(new_n304), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n725), .ZN(new_n730));
  INV_X1    g0530(.A(G317), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n731), .A2(KEYINPUT33), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(KEYINPUT33), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n725), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n728), .B(new_n734), .C1(G329), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n720), .A2(new_n725), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G311), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n230), .B1(new_n735), .B2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G294), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n719), .A2(new_n729), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n261), .B1(new_n746), .B2(G326), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n738), .A2(new_n741), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n719), .A2(new_n724), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n723), .B(new_n748), .C1(G303), .C2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n721), .B(KEYINPUT99), .Z(new_n752));
  OAI21_X1  g0552(.A(new_n261), .B1(new_n752), .B2(new_n219), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n730), .A2(new_n289), .B1(new_n742), .B2(new_n206), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT100), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT32), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n737), .B2(G159), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(G50), .B2(new_n746), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n737), .A2(new_n756), .A3(G159), .ZN(new_n759));
  INV_X1    g0559(.A(new_n726), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G77), .A2(new_n740), .B1(new_n760), .B2(G107), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n755), .A2(new_n758), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n753), .B(new_n762), .C1(G87), .C2(new_n750), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n718), .B1(new_n751), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n712), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n261), .A2(G355), .A3(new_n224), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n249), .A2(new_n438), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n393), .A2(new_n664), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G45), .B2(new_n229), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n766), .B1(G116), .B2(new_n224), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n718), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n765), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n773), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n764), .B(new_n775), .C1(new_n652), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n714), .A2(new_n777), .ZN(G396));
  OAI21_X1  g0578(.A(KEYINPUT104), .B1(new_n345), .B2(new_n649), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT104), .ZN(new_n780));
  INV_X1    g0580(.A(new_n343), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n216), .B2(new_n286), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n780), .B(new_n648), .C1(new_n782), .C2(new_n344), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n779), .B(new_n783), .C1(new_n432), .C2(new_n433), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n362), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n360), .A2(new_n361), .A3(new_n649), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT105), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n648), .B1(new_n624), .B2(new_n630), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n648), .B(new_n787), .C1(new_n624), .C2(new_n630), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(new_n690), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n765), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n718), .A2(new_n771), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n745), .A2(new_n797), .B1(new_n742), .B2(new_n206), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n760), .A2(G87), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n727), .B2(new_n730), .C1(new_n800), .C2(new_n736), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n798), .B(new_n801), .C1(G116), .C2(new_n740), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n802), .B(new_n369), .C1(new_n210), .C2(new_n749), .ZN(new_n803));
  INV_X1    g0603(.A(new_n721), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G294), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n730), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G137), .A2(new_n746), .B1(new_n806), .B2(G150), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  INV_X1    g0608(.A(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n739), .C1(new_n752), .C2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n749), .A2(new_n214), .B1(new_n726), .B2(new_n289), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT101), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n812), .A2(KEYINPUT101), .B1(G58), .B2(new_n743), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n393), .B1(new_n816), .B2(new_n736), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT102), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n805), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n718), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n712), .B1(G77), .B2(new_n796), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT103), .ZN(new_n822));
  INV_X1    g0622(.A(new_n787), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n772), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n794), .A2(new_n824), .ZN(G384));
  INV_X1    g0625(.A(KEYINPUT35), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n230), .B(new_n231), .C1(new_n558), .C2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n827), .B(G116), .C1(new_n826), .C2(new_n558), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  OAI21_X1  g0629(.A(G77), .B1(new_n219), .B2(new_n289), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n229), .A2(new_n830), .B1(G50), .B2(new_n289), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(G1), .A3(new_n278), .ZN(new_n832));
  XOR2_X1   g0632(.A(KEYINPUT110), .B(KEYINPUT38), .Z(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n646), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n408), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n431), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n420), .A2(new_n836), .A3(new_n429), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n834), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT108), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n395), .A2(KEYINPUT107), .A3(new_n380), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n397), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT107), .B1(new_n395), .B2(new_n380), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n843), .B(new_n284), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n396), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n395), .A2(new_n380), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT107), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(new_n397), .A3(new_n844), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n843), .B1(new_n852), .B2(new_n284), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n407), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n835), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT109), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(KEYINPUT109), .A3(new_n835), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n401), .A2(new_n404), .A3(new_n407), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n854), .A2(new_n419), .B1(new_n859), .B2(new_n428), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n842), .B1(new_n861), .B2(KEYINPUT37), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n430), .A2(new_n424), .B1(new_n857), .B2(new_n858), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n841), .B1(new_n864), .B2(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n671), .A2(KEYINPUT31), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n683), .A2(new_n648), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n685), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n301), .A2(new_n648), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n302), .A2(new_n307), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n276), .A2(new_n301), .A3(new_n648), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n787), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT40), .B1(new_n865), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT109), .B1(new_n854), .B2(new_n835), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n854), .A2(KEYINPUT109), .A3(new_n835), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n431), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n876), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n880), .B2(new_n860), .ZN(new_n881));
  OAI211_X1 g0681(.A(KEYINPUT38), .B(new_n878), .C1(new_n881), .C2(new_n842), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n862), .B2(new_n863), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(new_n873), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n868), .B2(new_n685), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n875), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n436), .A2(new_n869), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(G330), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n862), .A2(new_n883), .A3(new_n863), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n894), .B1(new_n895), .B2(new_n841), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n302), .A2(new_n648), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT39), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  INV_X1    g0700(.A(new_n786), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n789), .B2(new_n823), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n871), .A2(new_n872), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(KEYINPUT106), .B(new_n903), .C1(new_n791), .C2(new_n901), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n885), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n424), .A2(new_n835), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n899), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n436), .B1(new_n704), .B2(new_n702), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n639), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n893), .A2(new_n913), .B1(new_n254), .B2(new_n642), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT111), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n893), .A2(new_n913), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n829), .B(new_n832), .C1(new_n915), .C2(new_n916), .ZN(G367));
  NAND2_X1  g0717(.A1(new_n586), .A2(new_n596), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n625), .A2(new_n918), .A3(new_n648), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n648), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n612), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n765), .B1(new_n923), .B2(new_n773), .ZN(new_n924));
  INV_X1    g0724(.A(new_n768), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n774), .B1(new_n224), .B2(new_n585), .C1(new_n241), .C2(new_n925), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G283), .A2(new_n740), .B1(new_n737), .B2(G317), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n749), .A2(new_n499), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n927), .B1(KEYINPUT46), .B2(new_n928), .C1(new_n752), .C2(new_n797), .ZN(new_n929));
  INV_X1    g0729(.A(G294), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n730), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n928), .A2(KEYINPUT46), .ZN(new_n932));
  AOI22_X1  g0732(.A1(G311), .A2(new_n746), .B1(new_n760), .B2(G97), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n933), .B(new_n387), .C1(new_n210), .C2(new_n742), .ZN(new_n934));
  NOR4_X1   g0734(.A1(new_n929), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n726), .A2(new_n216), .ZN(new_n936));
  INV_X1    g0736(.A(G137), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n749), .A2(new_n219), .B1(new_n736), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT113), .Z(new_n939));
  OAI22_X1  g0739(.A1(new_n721), .A2(new_n326), .B1(new_n742), .B2(new_n289), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT112), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n940), .A2(new_n941), .B1(G159), .B2(new_n806), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n746), .A2(G143), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n939), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n936), .B(new_n945), .C1(G50), .C2(new_n740), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n935), .B1(new_n946), .B2(new_n261), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT47), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n924), .B(new_n926), .C1(new_n820), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n710), .A2(G1), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n620), .B1(new_n560), .B2(new_n649), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n619), .A2(new_n566), .A3(new_n648), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n662), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT45), .Z(new_n955));
  NOR2_X1   g0755(.A1(new_n662), .A2(new_n953), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n654), .B2(new_n660), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n658), .A2(new_n483), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n653), .A2(new_n659), .A3(new_n657), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n661), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n708), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n665), .B(KEYINPUT41), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n950), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n953), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(new_n960), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT42), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n571), .B1(new_n951), .B2(new_n482), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n649), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n968), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n661), .A2(new_n966), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n949), .B1(new_n965), .B2(new_n975), .ZN(G387));
  INV_X1    g0776(.A(new_n962), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n665), .B1(new_n708), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n962), .B1(new_n705), .B2(new_n707), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n657), .A2(new_n773), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n750), .A2(G294), .B1(new_n743), .B2(G283), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G311), .A2(new_n806), .B1(new_n740), .B2(G303), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n722), .B2(new_n745), .C1(new_n752), .C2(new_n731), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT48), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT115), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT49), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n737), .A2(G326), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n393), .B1(new_n760), .B2(G116), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G159), .A2(new_n746), .B1(new_n740), .B2(G68), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n750), .A2(G77), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n743), .A2(new_n341), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n737), .A2(G150), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n387), .B1(G50), .B2(new_n804), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n329), .A2(new_n806), .B1(new_n760), .B2(G97), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n820), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n925), .B1(new_n237), .B2(G45), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n339), .A2(new_n214), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1005), .A2(new_n1006), .A3(new_n438), .A4(new_n667), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n289), .A2(new_n216), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n261), .A2(new_n224), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(G107), .B2(new_n224), .C1(new_n667), .C2(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(KEYINPUT114), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(KEYINPUT114), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1012), .A2(new_n774), .A3(new_n1013), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n1002), .A2(new_n765), .A3(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n981), .A2(new_n1015), .B1(new_n977), .B2(new_n950), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n980), .A2(new_n1016), .ZN(G393));
  OAI22_X1  g0817(.A1(new_n745), .A2(new_n731), .B1(new_n721), .B2(new_n800), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT52), .Z(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G303), .B2(new_n806), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n210), .B2(new_n726), .C1(new_n499), .C2(new_n742), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n749), .A2(new_n727), .B1(new_n736), .B2(new_n722), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT116), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n369), .C1(new_n930), .C2(new_n739), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n749), .A2(new_n289), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n799), .B(new_n393), .C1(new_n216), .C2(new_n742), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G143), .B2(new_n737), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n806), .A2(G50), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n745), .A2(new_n326), .B1(new_n721), .B2(new_n808), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT51), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n339), .A2(new_n740), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1021), .A2(new_n1024), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n765), .B1(new_n1033), .B2(new_n718), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n953), .B2(new_n776), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n245), .A2(new_n768), .B1(G97), .B2(new_n664), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n774), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n958), .B(new_n661), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n950), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n959), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n979), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n979), .B2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1039), .B1(new_n1042), .B2(new_n666), .ZN(G390));
  INV_X1    g0843(.A(KEYINPUT117), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n896), .A2(new_n898), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n897), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n902), .B2(new_n904), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n838), .A2(new_n840), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n833), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n882), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n701), .A2(new_n649), .A3(new_n785), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n786), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n897), .B1(new_n1052), .B2(new_n903), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1045), .A2(new_n1047), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(G330), .B(new_n823), .C1(new_n684), .C2(new_n689), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(new_n904), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1044), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n882), .A2(new_n884), .A3(KEYINPUT39), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT39), .B1(new_n882), .B2(new_n1049), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1047), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1053), .A2(new_n1050), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1060), .A2(new_n1044), .A3(new_n1061), .A4(new_n1056), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1065));
  INV_X1    g0865(.A(G330), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n874), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n950), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT119), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n721), .A2(new_n816), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n742), .A2(new_n808), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n750), .A2(G150), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT53), .ZN(new_n1074));
  INV_X1    g0874(.A(G128), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n745), .A2(new_n1075), .B1(new_n726), .B2(new_n214), .ZN(new_n1076));
  INV_X1    g0876(.A(G125), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n261), .B1(new_n736), .B2(new_n1077), .C1(new_n937), .C2(new_n730), .ZN(new_n1078));
  OR4_X1    g0878(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(KEYINPUT54), .B(G143), .Z(new_n1080));
  AOI211_X1 g0880(.A(new_n1071), .B(new_n1079), .C1(new_n740), .C2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n726), .A2(new_n289), .B1(new_n736), .B2(new_n930), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1082), .A2(KEYINPUT118), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n261), .B1(new_n804), .B2(G116), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n204), .B2(new_n749), .C1(new_n210), .C2(new_n730), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1082), .A2(KEYINPUT118), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n739), .A2(new_n206), .B1(new_n742), .B2(new_n216), .ZN(new_n1087));
  OR4_X1    g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G283), .B2(new_n746), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n718), .B1(new_n1081), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n712), .C1(new_n329), .C2(new_n796), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1045), .A2(new_n771), .B1(new_n1070), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n1070), .B2(new_n1091), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n911), .B(new_n639), .C1(new_n891), .C2(new_n1066), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n869), .A2(G330), .A3(new_n788), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n904), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1096), .A2(new_n1056), .A3(new_n786), .A4(new_n1051), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n888), .A2(G330), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1055), .A2(new_n904), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n786), .B1(new_n703), .B2(new_n787), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1094), .B1(new_n1097), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1060), .A2(new_n1061), .A3(new_n1056), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1106), .A2(new_n1068), .A3(new_n1062), .A4(new_n1103), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n665), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1069), .B(new_n1093), .C1(new_n1104), .C2(new_n1108), .ZN(G378));
  INV_X1    g0909(.A(KEYINPUT57), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1094), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n334), .A2(new_n336), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT55), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n331), .A2(new_n835), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1066), .B1(new_n875), .B2(new_n889), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1120), .A2(new_n910), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n910), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n886), .B1(new_n1050), .B2(new_n888), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n685), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n873), .B(new_n886), .C1(new_n684), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n882), .B2(new_n884), .ZN(new_n1127));
  OAI21_X1  g0927(.A(G330), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1128), .A2(new_n909), .A3(new_n899), .A4(new_n907), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1120), .A2(new_n910), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(new_n1118), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1110), .B1(new_n1112), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1129), .A2(new_n1130), .A3(new_n1118), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1118), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1134), .A2(new_n1135), .A3(new_n1110), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n665), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(G41), .B1(new_n746), .B2(G116), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n740), .A2(new_n341), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1140), .A2(new_n387), .A3(new_n995), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n760), .A2(G58), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n289), .B2(new_n742), .C1(new_n727), .C2(new_n736), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G107), .C2(new_n804), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n206), .B2(new_n730), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT58), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n391), .A2(new_n392), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n1148), .B2(G33), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n739), .A2(new_n937), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n745), .A2(new_n1077), .B1(new_n742), .B2(new_n326), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT120), .Z(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(new_n750), .C2(new_n1080), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n1075), .B2(new_n721), .C1(new_n816), .C2(new_n730), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G33), .B1(new_n737), .B2(G124), .ZN(new_n1156));
  INV_X1    g0956(.A(G41), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n808), .C2(new_n726), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT121), .Z(new_n1159));
  OAI221_X1 g0959(.A(new_n1147), .B1(G50), .B2(new_n1149), .C1(new_n1155), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n765), .B1(new_n1160), .B2(new_n718), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1118), .B2(new_n772), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n796), .A2(G50), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n950), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1139), .A2(new_n1166), .ZN(G375));
  INV_X1    g0967(.A(new_n1103), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1097), .A2(new_n1102), .A3(new_n1094), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n964), .B(KEYINPUT123), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1143), .B1(new_n816), .B2(new_n745), .C1(new_n808), .C2(new_n749), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n752), .A2(new_n937), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G50), .C2(new_n743), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n387), .B1(G150), .B2(new_n740), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n1075), .C2(new_n736), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n806), .B2(new_n1080), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n721), .A2(new_n727), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n216), .A2(new_n726), .B1(new_n739), .B2(new_n210), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n996), .B1(new_n930), .B2(new_n745), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G303), .C2(new_n737), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n369), .C1(new_n206), .C2(new_n749), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1178), .B(new_n1182), .C1(G116), .C2(new_n806), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n718), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n712), .C1(G68), .C2(new_n796), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n904), .B2(new_n771), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n950), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1171), .A2(new_n1188), .ZN(G381));
  NOR2_X1   g0989(.A1(G375), .A2(G378), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G393), .A2(G396), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(G387), .A2(G390), .ZN(new_n1193));
  INV_X1    g0993(.A(G384), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1192), .A2(G381), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT124), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(G407));
  NAND2_X1  g0998(.A1(new_n647), .A2(G213), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT125), .Z(new_n1200));
  NAND2_X1  g1000(.A1(new_n1190), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(G407), .A2(G213), .A3(new_n1201), .ZN(G409));
  AND2_X1   g1002(.A1(G393), .A2(G396), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(new_n1191), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1193), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(G387), .A2(G390), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(KEYINPUT127), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT127), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1206), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n1193), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1204), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1210), .A2(new_n1204), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT60), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n666), .B1(new_n1169), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n1168), .C1(new_n1214), .C2(new_n1169), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1188), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1217), .A2(new_n1194), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1194), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1200), .A2(G2897), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(G2897), .A3(new_n1200), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1165), .A2(new_n1137), .A3(new_n1170), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G378), .B1(new_n1226), .B2(new_n1166), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1123), .A2(KEYINPUT57), .A3(new_n1131), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n665), .B1(new_n1112), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1165), .B2(new_n1137), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G378), .B(new_n1166), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT126), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT126), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1139), .A2(new_n1233), .A3(G378), .A4(new_n1166), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1227), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1223), .B(new_n1225), .C1(new_n1235), .C2(new_n1200), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1235), .A2(new_n1200), .A3(new_n1224), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1227), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n950), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1132), .A2(new_n1241), .B1(new_n1163), .B2(new_n1162), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n666), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(new_n1133), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1233), .B1(new_n1244), .B2(G378), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1231), .A2(KEYINPUT126), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1240), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1200), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1238), .A3(new_n1248), .A4(new_n1221), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1213), .B1(new_n1239), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1247), .A2(new_n1248), .A3(new_n1221), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1237), .B2(KEYINPUT63), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1252), .A2(new_n1260), .ZN(G405));
  NAND2_X1  g1061(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1244), .A2(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(new_n1221), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(new_n1213), .ZN(G402));
endmodule


