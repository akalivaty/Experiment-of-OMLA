

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G651), .A2(n575), .ZN(n669) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n783) );
  AND2_X1 U555 ( .A1(n547), .A2(G2105), .ZN(n995) );
  NOR2_X1 U556 ( .A1(n770), .A2(n769), .ZN(n771) );
  AND2_X1 U557 ( .A1(n528), .A2(n522), .ZN(n762) );
  NAND2_X2 U558 ( .A1(n783), .A2(n701), .ZN(n744) );
  AND2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n996) );
  AND2_X1 U560 ( .A1(n526), .A2(n532), .ZN(n525) );
  NAND2_X1 U561 ( .A1(n525), .A2(n524), .ZN(n523) );
  XNOR2_X1 U562 ( .A(n718), .B(KEYINPUT26), .ZN(n524) );
  INV_X1 U563 ( .A(n744), .ZN(n723) );
  INV_X1 U564 ( .A(KEYINPUT31), .ZN(n711) );
  NAND2_X1 U565 ( .A1(n752), .A2(G8), .ZN(n529) );
  NAND2_X1 U566 ( .A1(n700), .A2(n699), .ZN(n782) );
  NAND2_X1 U567 ( .A1(n554), .A2(n547), .ZN(n527) );
  XNOR2_X1 U568 ( .A(n529), .B(n753), .ZN(n819) );
  OR2_X1 U569 ( .A1(n761), .A2(n911), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n720), .A2(n523), .ZN(n721) );
  INV_X1 U571 ( .A(n962), .ZN(n526) );
  XNOR2_X2 U572 ( .A(n527), .B(KEYINPUT17), .ZN(n999) );
  NAND2_X1 U573 ( .A1(n819), .A2(n759), .ZN(n528) );
  NAND2_X1 U574 ( .A1(n530), .A2(G286), .ZN(n743) );
  NAND2_X1 U575 ( .A1(n530), .A2(n755), .ZN(n756) );
  NAND2_X1 U576 ( .A1(n741), .A2(n742), .ZN(n530) );
  INV_X1 U577 ( .A(n782), .ZN(n701) );
  NOR2_X1 U578 ( .A1(n764), .A2(KEYINPUT33), .ZN(n766) );
  XNOR2_X1 U579 ( .A(n766), .B(n765), .ZN(n770) );
  NOR2_X1 U580 ( .A1(n754), .A2(n702), .ZN(n531) );
  OR2_X1 U581 ( .A1(n723), .A2(n719), .ZN(n532) );
  AND2_X1 U582 ( .A1(n553), .A2(n552), .ZN(n533) );
  INV_X1 U583 ( .A(G8), .ZN(n702) );
  OR2_X1 U584 ( .A1(n963), .A2(n717), .ZN(n722) );
  INV_X1 U585 ( .A(KEYINPUT29), .ZN(n736) );
  XNOR2_X1 U586 ( .A(n737), .B(n736), .ZN(n740) );
  INV_X1 U587 ( .A(KEYINPUT99), .ZN(n765) );
  XNOR2_X1 U588 ( .A(KEYINPUT15), .B(n609), .ZN(n914) );
  XNOR2_X1 U589 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U590 ( .A(G1348), .B(G2427), .ZN(n543) );
  XOR2_X1 U591 ( .A(G2451), .B(G2430), .Z(n535) );
  INV_X1 U592 ( .A(G1341), .ZN(n719) );
  XOR2_X1 U593 ( .A(n719), .B(G2443), .Z(n534) );
  XNOR2_X1 U594 ( .A(n535), .B(n534), .ZN(n539) );
  XOR2_X1 U595 ( .A(G2438), .B(G2435), .Z(n537) );
  XNOR2_X1 U596 ( .A(KEYINPUT101), .B(G2454), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U598 ( .A(n539), .B(n538), .Z(n541) );
  XNOR2_X1 U599 ( .A(G2446), .B(KEYINPUT102), .ZN(n540) );
  XNOR2_X1 U600 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n543), .B(n542), .ZN(n544) );
  AND2_X1 U602 ( .A1(n544), .A2(G14), .ZN(G401) );
  NAND2_X1 U603 ( .A1(n999), .A2(G137), .ZN(n700) );
  INV_X1 U604 ( .A(G2105), .ZN(n554) );
  AND2_X1 U605 ( .A1(G101), .A2(n554), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G2104), .A2(n545), .ZN(n546) );
  XNOR2_X1 U607 ( .A(KEYINPUT23), .B(n546), .ZN(n551) );
  INV_X1 U608 ( .A(G2104), .ZN(n547) );
  NAND2_X1 U609 ( .A1(G125), .A2(n995), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G113), .A2(n996), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n698) );
  AND2_X1 U613 ( .A1(n700), .A2(n698), .ZN(G160) );
  AND2_X1 U614 ( .A1(n999), .A2(G138), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G126), .A2(n995), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G114), .A2(n996), .ZN(n552) );
  AND2_X1 U617 ( .A1(G2104), .A2(n554), .ZN(n1001) );
  NAND2_X1 U618 ( .A1(G102), .A2(n1001), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n533), .A2(n555), .ZN(n556) );
  NOR2_X1 U620 ( .A1(n557), .A2(n556), .ZN(G164) );
  NAND2_X1 U621 ( .A1(G123), .A2(n995), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(KEYINPUT18), .ZN(n565) );
  NAND2_X1 U623 ( .A1(G99), .A2(n1001), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G111), .A2(n996), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G135), .A2(n999), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT73), .B(n561), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT74), .B(n566), .ZN(n1020) );
  XNOR2_X1 U631 ( .A(n1020), .B(G2096), .ZN(n567) );
  OR2_X1 U632 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  INV_X1 U635 ( .A(G120), .ZN(G236) );
  INV_X1 U636 ( .A(G69), .ZN(G235) );
  INV_X1 U637 ( .A(G108), .ZN(G238) );
  NOR2_X1 U638 ( .A1(G651), .A2(G543), .ZN(n660) );
  NAND2_X1 U639 ( .A1(n660), .A2(G89), .ZN(n568) );
  XNOR2_X1 U640 ( .A(n568), .B(KEYINPUT4), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT0), .B(G543), .Z(n575) );
  INV_X1 U642 ( .A(G651), .ZN(n572) );
  NOR2_X1 U643 ( .A1(n575), .A2(n572), .ZN(n665) );
  NAND2_X1 U644 ( .A1(G76), .A2(n665), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U646 ( .A(KEYINPUT5), .B(n571), .ZN(n581) );
  NOR2_X1 U647 ( .A1(G543), .A2(n572), .ZN(n574) );
  XNOR2_X1 U648 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n573) );
  XNOR2_X1 U649 ( .A(n574), .B(n573), .ZN(n661) );
  NAND2_X1 U650 ( .A1(G63), .A2(n661), .ZN(n577) );
  NAND2_X1 U651 ( .A1(G51), .A2(n669), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n579) );
  XOR2_X1 U653 ( .A(KEYINPUT70), .B(KEYINPUT6), .Z(n578) );
  XNOR2_X1 U654 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U656 ( .A(KEYINPUT7), .B(n582), .ZN(G168) );
  NAND2_X1 U657 ( .A1(G94), .A2(G452), .ZN(n583) );
  XOR2_X1 U658 ( .A(KEYINPUT68), .B(n583), .Z(G173) );
  NAND2_X1 U659 ( .A1(G7), .A2(G661), .ZN(n584) );
  XOR2_X1 U660 ( .A(n584), .B(KEYINPUT10), .Z(n1032) );
  NAND2_X1 U661 ( .A1(n1032), .A2(G567), .ZN(n585) );
  XOR2_X1 U662 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U663 ( .A1(G56), .A2(n661), .ZN(n586) );
  XOR2_X1 U664 ( .A(KEYINPUT14), .B(n586), .Z(n592) );
  NAND2_X1 U665 ( .A1(n660), .A2(G81), .ZN(n587) );
  XNOR2_X1 U666 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U667 ( .A1(G68), .A2(n665), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U669 ( .A(KEYINPUT13), .B(n590), .Z(n591) );
  NOR2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n669), .A2(G43), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n962) );
  INV_X1 U673 ( .A(G860), .ZN(n631) );
  OR2_X1 U674 ( .A1(n962), .A2(n631), .ZN(G153) );
  NAND2_X1 U675 ( .A1(G64), .A2(n661), .ZN(n596) );
  NAND2_X1 U676 ( .A1(G52), .A2(n669), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n601) );
  NAND2_X1 U678 ( .A1(G90), .A2(n660), .ZN(n598) );
  NAND2_X1 U679 ( .A1(G77), .A2(n665), .ZN(n597) );
  NAND2_X1 U680 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U681 ( .A(KEYINPUT9), .B(n599), .Z(n600) );
  NOR2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U683 ( .A(KEYINPUT67), .B(n602), .ZN(G301) );
  NAND2_X1 U684 ( .A1(G868), .A2(G301), .ZN(n611) );
  NAND2_X1 U685 ( .A1(G92), .A2(n660), .ZN(n604) );
  NAND2_X1 U686 ( .A1(G66), .A2(n661), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G79), .A2(n665), .ZN(n606) );
  NAND2_X1 U689 ( .A1(G54), .A2(n669), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n609) );
  INV_X1 U692 ( .A(G868), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n914), .A2(n624), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n611), .A2(n610), .ZN(G284) );
  NAND2_X1 U695 ( .A1(G78), .A2(n665), .ZN(n613) );
  NAND2_X1 U696 ( .A1(G65), .A2(n661), .ZN(n612) );
  NAND2_X1 U697 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G91), .A2(n660), .ZN(n614) );
  XNOR2_X1 U699 ( .A(KEYINPUT69), .B(n614), .ZN(n615) );
  NOR2_X1 U700 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n669), .A2(G53), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(G299) );
  XOR2_X1 U703 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U704 ( .A1(G868), .A2(G299), .ZN(n620) );
  NOR2_X1 U705 ( .A1(G286), .A2(n624), .ZN(n619) );
  NOR2_X1 U706 ( .A1(n620), .A2(n619), .ZN(G297) );
  NAND2_X1 U707 ( .A1(n631), .A2(G559), .ZN(n621) );
  INV_X1 U708 ( .A(n914), .ZN(n963) );
  NAND2_X1 U709 ( .A1(n621), .A2(n963), .ZN(n622) );
  XNOR2_X1 U710 ( .A(n622), .B(KEYINPUT16), .ZN(n623) );
  XOR2_X1 U711 ( .A(KEYINPUT71), .B(n623), .Z(G148) );
  NOR2_X1 U712 ( .A1(n914), .A2(n624), .ZN(n625) );
  XOR2_X1 U713 ( .A(KEYINPUT72), .B(n625), .Z(n626) );
  NOR2_X1 U714 ( .A1(G559), .A2(n626), .ZN(n628) );
  NOR2_X1 U715 ( .A1(G868), .A2(n962), .ZN(n627) );
  NOR2_X1 U716 ( .A1(n628), .A2(n627), .ZN(G282) );
  XNOR2_X1 U717 ( .A(n962), .B(KEYINPUT75), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n963), .A2(G559), .ZN(n629) );
  XNOR2_X1 U719 ( .A(n630), .B(n629), .ZN(n677) );
  NAND2_X1 U720 ( .A1(n631), .A2(n677), .ZN(n638) );
  NAND2_X1 U721 ( .A1(G67), .A2(n661), .ZN(n633) );
  NAND2_X1 U722 ( .A1(G55), .A2(n669), .ZN(n632) );
  NAND2_X1 U723 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U724 ( .A1(G93), .A2(n660), .ZN(n635) );
  NAND2_X1 U725 ( .A1(G80), .A2(n665), .ZN(n634) );
  NAND2_X1 U726 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U727 ( .A1(n637), .A2(n636), .ZN(n679) );
  XOR2_X1 U728 ( .A(n638), .B(n679), .Z(G145) );
  NAND2_X1 U729 ( .A1(G49), .A2(n669), .ZN(n640) );
  NAND2_X1 U730 ( .A1(G87), .A2(n575), .ZN(n639) );
  NAND2_X1 U731 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U732 ( .A1(n661), .A2(n641), .ZN(n643) );
  NAND2_X1 U733 ( .A1(G651), .A2(G74), .ZN(n642) );
  NAND2_X1 U734 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G85), .A2(n660), .ZN(n645) );
  NAND2_X1 U736 ( .A1(G72), .A2(n665), .ZN(n644) );
  NAND2_X1 U737 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U738 ( .A(KEYINPUT64), .B(n646), .ZN(n650) );
  NAND2_X1 U739 ( .A1(G60), .A2(n661), .ZN(n648) );
  NAND2_X1 U740 ( .A1(G47), .A2(n669), .ZN(n647) );
  NAND2_X1 U741 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U742 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U743 ( .A(KEYINPUT66), .B(n651), .Z(G290) );
  NAND2_X1 U744 ( .A1(n669), .A2(G50), .ZN(n653) );
  NAND2_X1 U745 ( .A1(n661), .A2(G62), .ZN(n652) );
  NAND2_X1 U746 ( .A1(n653), .A2(n652), .ZN(n658) );
  NAND2_X1 U747 ( .A1(G88), .A2(n660), .ZN(n655) );
  NAND2_X1 U748 ( .A1(G75), .A2(n665), .ZN(n654) );
  NAND2_X1 U749 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U750 ( .A(KEYINPUT77), .B(n656), .Z(n657) );
  NOR2_X1 U751 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U752 ( .A(KEYINPUT78), .B(n659), .ZN(G166) );
  INV_X1 U753 ( .A(G166), .ZN(G303) );
  NAND2_X1 U754 ( .A1(G86), .A2(n660), .ZN(n663) );
  NAND2_X1 U755 ( .A1(G61), .A2(n661), .ZN(n662) );
  NAND2_X1 U756 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U757 ( .A(KEYINPUT76), .B(n664), .ZN(n668) );
  NAND2_X1 U758 ( .A1(n665), .A2(G73), .ZN(n666) );
  XOR2_X1 U759 ( .A(KEYINPUT2), .B(n666), .Z(n667) );
  NOR2_X1 U760 ( .A1(n668), .A2(n667), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n669), .A2(G48), .ZN(n670) );
  NAND2_X1 U762 ( .A1(n671), .A2(n670), .ZN(G305) );
  XOR2_X1 U763 ( .A(n679), .B(KEYINPUT19), .Z(n672) );
  XNOR2_X1 U764 ( .A(G288), .B(n672), .ZN(n673) );
  XOR2_X1 U765 ( .A(G299), .B(n673), .Z(n676) );
  XOR2_X1 U766 ( .A(G290), .B(G303), .Z(n674) );
  XNOR2_X1 U767 ( .A(n674), .B(G305), .ZN(n675) );
  XNOR2_X1 U768 ( .A(n676), .B(n675), .ZN(n966) );
  XNOR2_X1 U769 ( .A(n677), .B(n966), .ZN(n678) );
  NAND2_X1 U770 ( .A1(n678), .A2(G868), .ZN(n681) );
  OR2_X1 U771 ( .A1(G868), .A2(n679), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n681), .A2(n680), .ZN(G295) );
  XOR2_X1 U773 ( .A(KEYINPUT79), .B(KEYINPUT21), .Z(n685) );
  NAND2_X1 U774 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U775 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U776 ( .A1(n683), .A2(G2090), .ZN(n684) );
  XNOR2_X1 U777 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U778 ( .A1(G2072), .A2(n686), .ZN(G158) );
  NOR2_X1 U779 ( .A1(G235), .A2(G236), .ZN(n687) );
  XOR2_X1 U780 ( .A(KEYINPUT80), .B(n687), .Z(n688) );
  NOR2_X1 U781 ( .A1(G238), .A2(n688), .ZN(n689) );
  NAND2_X1 U782 ( .A1(G57), .A2(n689), .ZN(n960) );
  NAND2_X1 U783 ( .A1(G567), .A2(n960), .ZN(n690) );
  XNOR2_X1 U784 ( .A(n690), .B(KEYINPUT81), .ZN(n695) );
  NOR2_X1 U785 ( .A1(G220), .A2(G219), .ZN(n691) );
  XNOR2_X1 U786 ( .A(KEYINPUT22), .B(n691), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n692), .A2(G96), .ZN(n693) );
  OR2_X1 U788 ( .A1(G218), .A2(n693), .ZN(n961) );
  AND2_X1 U789 ( .A1(G2106), .A2(n961), .ZN(n694) );
  NOR2_X1 U790 ( .A1(n695), .A2(n694), .ZN(G319) );
  INV_X1 U791 ( .A(G319), .ZN(n1024) );
  NAND2_X1 U792 ( .A1(G661), .A2(G483), .ZN(n696) );
  NOR2_X1 U793 ( .A1(n1024), .A2(n696), .ZN(n839) );
  NAND2_X1 U794 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U795 ( .A(G301), .ZN(G171) );
  AND2_X1 U796 ( .A1(n698), .A2(G40), .ZN(n699) );
  NAND2_X1 U797 ( .A1(G8), .A2(n744), .ZN(n827) );
  NOR2_X1 U798 ( .A1(G1966), .A2(n827), .ZN(n757) );
  INV_X1 U799 ( .A(n757), .ZN(n703) );
  NOR2_X1 U800 ( .A1(G2084), .A2(n744), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n703), .A2(n531), .ZN(n704) );
  XNOR2_X1 U802 ( .A(n704), .B(KEYINPUT30), .ZN(n705) );
  NOR2_X1 U803 ( .A1(G168), .A2(n705), .ZN(n706) );
  XNOR2_X1 U804 ( .A(n706), .B(KEYINPUT92), .ZN(n710) );
  XOR2_X1 U805 ( .A(G1961), .B(KEYINPUT86), .Z(n935) );
  NAND2_X1 U806 ( .A1(n935), .A2(n744), .ZN(n708) );
  XNOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .ZN(n885) );
  NAND2_X1 U808 ( .A1(n723), .A2(n885), .ZN(n707) );
  NAND2_X1 U809 ( .A1(n708), .A2(n707), .ZN(n738) );
  NOR2_X1 U810 ( .A1(n738), .A2(G171), .ZN(n709) );
  NOR2_X1 U811 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U812 ( .A(n712), .B(n711), .ZN(n742) );
  NAND2_X1 U813 ( .A1(n723), .A2(G2067), .ZN(n713) );
  XNOR2_X1 U814 ( .A(KEYINPUT91), .B(n713), .ZN(n716) );
  NAND2_X1 U815 ( .A1(G1348), .A2(n744), .ZN(n714) );
  XOR2_X1 U816 ( .A(KEYINPUT90), .B(n714), .Z(n715) );
  NOR2_X1 U817 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U818 ( .A1(n963), .A2(n717), .ZN(n720) );
  XOR2_X1 U819 ( .A(G1996), .B(KEYINPUT89), .Z(n886) );
  NAND2_X1 U820 ( .A1(n723), .A2(n886), .ZN(n718) );
  NAND2_X1 U821 ( .A1(n722), .A2(n721), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n723), .A2(G2072), .ZN(n724) );
  XNOR2_X1 U823 ( .A(KEYINPUT27), .B(n724), .ZN(n727) );
  NAND2_X1 U824 ( .A1(G1956), .A2(n744), .ZN(n725) );
  XNOR2_X1 U825 ( .A(KEYINPUT87), .B(n725), .ZN(n726) );
  NOR2_X1 U826 ( .A1(n727), .A2(n726), .ZN(n731) );
  INV_X1 U827 ( .A(G299), .ZN(n730) );
  NAND2_X1 U828 ( .A1(n731), .A2(n730), .ZN(n728) );
  NAND2_X1 U829 ( .A1(n729), .A2(n728), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n731), .A2(n730), .ZN(n733) );
  XOR2_X1 U831 ( .A(KEYINPUT28), .B(KEYINPUT88), .Z(n732) );
  XNOR2_X1 U832 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U833 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U834 ( .A1(n738), .A2(G171), .ZN(n739) );
  NAND2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U836 ( .A(n743), .B(KEYINPUT94), .ZN(n750) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n744), .ZN(n745) );
  XNOR2_X1 U838 ( .A(KEYINPUT95), .B(n745), .ZN(n748) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n827), .ZN(n746) );
  NOR2_X1 U840 ( .A1(G166), .A2(n746), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U843 ( .A(n751), .B(KEYINPUT96), .ZN(n752) );
  XOR2_X1 U844 ( .A(KEYINPUT32), .B(KEYINPUT97), .Z(n753) );
  NAND2_X1 U845 ( .A1(G8), .A2(n754), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U847 ( .A(KEYINPUT93), .B(n758), .ZN(n820) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n917) );
  AND2_X1 U849 ( .A1(n820), .A2(n917), .ZN(n759) );
  INV_X1 U850 ( .A(n917), .ZN(n761) );
  NOR2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G303), .A2(G1971), .ZN(n760) );
  NOR2_X1 U853 ( .A1(n767), .A2(n760), .ZN(n911) );
  XNOR2_X1 U854 ( .A(n762), .B(KEYINPUT98), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n827), .A2(n763), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n767), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U857 ( .A1(n827), .A2(n768), .ZN(n769) );
  XNOR2_X1 U858 ( .A(n771), .B(KEYINPUT100), .ZN(n808) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n906) );
  NAND2_X1 U860 ( .A1(G104), .A2(n1001), .ZN(n773) );
  NAND2_X1 U861 ( .A1(G140), .A2(n999), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U863 ( .A(KEYINPUT34), .B(n774), .ZN(n780) );
  NAND2_X1 U864 ( .A1(n996), .A2(G116), .ZN(n775) );
  XOR2_X1 U865 ( .A(KEYINPUT83), .B(n775), .Z(n777) );
  NAND2_X1 U866 ( .A1(n995), .A2(G128), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U868 ( .A(KEYINPUT35), .B(n778), .Z(n779) );
  NOR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U870 ( .A(KEYINPUT36), .B(n781), .ZN(n1007) );
  XNOR2_X1 U871 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NOR2_X1 U872 ( .A1(n1007), .A2(n815), .ZN(n871) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n818) );
  NAND2_X1 U874 ( .A1(n871), .A2(n818), .ZN(n813) );
  INV_X1 U875 ( .A(n813), .ZN(n805) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n912) );
  NAND2_X1 U877 ( .A1(n912), .A2(n818), .ZN(n784) );
  XNOR2_X1 U878 ( .A(n784), .B(KEYINPUT82), .ZN(n803) );
  NAND2_X1 U879 ( .A1(G129), .A2(n995), .ZN(n786) );
  NAND2_X1 U880 ( .A1(G117), .A2(n996), .ZN(n785) );
  NAND2_X1 U881 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n1001), .A2(G105), .ZN(n787) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n999), .A2(G141), .ZN(n790) );
  NAND2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n1010) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n1010), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G107), .A2(n996), .ZN(n792) );
  XNOR2_X1 U889 ( .A(n792), .B(KEYINPUT84), .ZN(n799) );
  NAND2_X1 U890 ( .A1(G95), .A2(n1001), .ZN(n794) );
  NAND2_X1 U891 ( .A1(G119), .A2(n995), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U893 ( .A1(G131), .A2(n999), .ZN(n795) );
  XNOR2_X1 U894 ( .A(KEYINPUT85), .B(n795), .ZN(n796) );
  NOR2_X1 U895 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n1009) );
  NAND2_X1 U897 ( .A1(G1991), .A2(n1009), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n865) );
  NAND2_X1 U899 ( .A1(n865), .A2(n818), .ZN(n802) );
  NAND2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n831) );
  INV_X1 U902 ( .A(n831), .ZN(n806) );
  AND2_X1 U903 ( .A1(n906), .A2(n806), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n835) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n1010), .ZN(n862) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n1009), .ZN(n867) );
  NOR2_X1 U908 ( .A1(n809), .A2(n867), .ZN(n810) );
  NOR2_X1 U909 ( .A1(n865), .A2(n810), .ZN(n811) );
  NOR2_X1 U910 ( .A1(n862), .A2(n811), .ZN(n812) );
  XNOR2_X1 U911 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n1007), .A2(n815), .ZN(n875) );
  NAND2_X1 U914 ( .A1(n816), .A2(n875), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n833) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n823) );
  NOR2_X1 U917 ( .A1(G2090), .A2(G303), .ZN(n821) );
  NAND2_X1 U918 ( .A1(G8), .A2(n821), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  AND2_X1 U920 ( .A1(n824), .A2(n827), .ZN(n829) );
  NOR2_X1 U921 ( .A1(G1981), .A2(G305), .ZN(n825) );
  XOR2_X1 U922 ( .A(n825), .B(KEYINPUT24), .Z(n826) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  OR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  AND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U928 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n1032), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U931 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(G188) );
  NAND2_X1 U935 ( .A1(G124), .A2(n995), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n840), .B(KEYINPUT110), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G100), .A2(n1001), .ZN(n842) );
  NAND2_X1 U939 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U940 ( .A1(G136), .A2(n999), .ZN(n845) );
  NAND2_X1 U941 ( .A1(G112), .A2(n996), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G162) );
  NAND2_X1 U944 ( .A1(G103), .A2(n1001), .ZN(n849) );
  NAND2_X1 U945 ( .A1(G139), .A2(n999), .ZN(n848) );
  NAND2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n855) );
  NAND2_X1 U947 ( .A1(n996), .A2(G115), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT112), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G127), .A2(n995), .ZN(n851) );
  NAND2_X1 U950 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT47), .B(n853), .Z(n854) );
  NOR2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n1019) );
  XNOR2_X1 U953 ( .A(n1019), .B(G2072), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n856), .B(KEYINPUT120), .ZN(n859) );
  XOR2_X1 U955 ( .A(G164), .B(G2078), .Z(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT121), .B(n857), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT50), .B(n860), .ZN(n878) );
  XOR2_X1 U959 ( .A(G2090), .B(G162), .Z(n861) );
  NOR2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n863), .B(KEYINPUT51), .ZN(n864) );
  NOR2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n873) );
  XNOR2_X1 U963 ( .A(G160), .B(G2084), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n866), .A2(n1020), .ZN(n868) );
  NOR2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U966 ( .A(KEYINPUT118), .B(n869), .Z(n870) );
  NOR2_X1 U967 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U969 ( .A(n874), .B(KEYINPUT119), .ZN(n876) );
  NAND2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U971 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U972 ( .A(KEYINPUT52), .B(n879), .Z(n880) );
  NOR2_X1 U973 ( .A1(KEYINPUT55), .A2(n880), .ZN(n881) );
  XOR2_X1 U974 ( .A(KEYINPUT122), .B(n881), .Z(n882) );
  NAND2_X1 U975 ( .A1(G29), .A2(n882), .ZN(n958) );
  XNOR2_X1 U976 ( .A(G2072), .B(G33), .ZN(n884) );
  XNOR2_X1 U977 ( .A(G2067), .B(G26), .ZN(n883) );
  NOR2_X1 U978 ( .A1(n884), .A2(n883), .ZN(n890) );
  XOR2_X1 U979 ( .A(n885), .B(G27), .Z(n888) );
  XNOR2_X1 U980 ( .A(G32), .B(n886), .ZN(n887) );
  NOR2_X1 U981 ( .A1(n888), .A2(n887), .ZN(n889) );
  NAND2_X1 U982 ( .A1(n890), .A2(n889), .ZN(n895) );
  XNOR2_X1 U983 ( .A(G1991), .B(KEYINPUT123), .ZN(n891) );
  XNOR2_X1 U984 ( .A(n891), .B(G25), .ZN(n892) );
  NAND2_X1 U985 ( .A1(G28), .A2(n892), .ZN(n893) );
  XNOR2_X1 U986 ( .A(KEYINPUT124), .B(n893), .ZN(n894) );
  NOR2_X1 U987 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U988 ( .A(KEYINPUT53), .B(n896), .Z(n899) );
  XOR2_X1 U989 ( .A(G34), .B(KEYINPUT54), .Z(n897) );
  XNOR2_X1 U990 ( .A(G2084), .B(n897), .ZN(n898) );
  NAND2_X1 U991 ( .A1(n899), .A2(n898), .ZN(n901) );
  XNOR2_X1 U992 ( .A(G35), .B(G2090), .ZN(n900) );
  NOR2_X1 U993 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U994 ( .A(KEYINPUT55), .B(n902), .Z(n903) );
  NOR2_X1 U995 ( .A1(G29), .A2(n903), .ZN(n904) );
  XNOR2_X1 U996 ( .A(KEYINPUT125), .B(n904), .ZN(n905) );
  NAND2_X1 U997 ( .A1(n905), .A2(G11), .ZN(n956) );
  INV_X1 U998 ( .A(G16), .ZN(n952) );
  XOR2_X1 U999 ( .A(n952), .B(KEYINPUT56), .Z(n928) );
  XNOR2_X1 U1000 ( .A(G168), .B(G1966), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n908), .B(KEYINPUT57), .ZN(n926) );
  XOR2_X1 U1003 ( .A(G1341), .B(n962), .Z(n910) );
  NAND2_X1 U1004 ( .A1(G1971), .A2(G303), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n924) );
  INV_X1 U1006 ( .A(n911), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(n922) );
  XOR2_X1 U1008 ( .A(n914), .B(G1348), .Z(n916) );
  XOR2_X1 U1009 ( .A(G301), .B(G1961), .Z(n915) );
  NAND2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n920) );
  XOR2_X1 U1011 ( .A(G299), .B(G1956), .Z(n918) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1015 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1016 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1017 ( .A1(n928), .A2(n927), .ZN(n954) );
  XNOR2_X1 U1018 ( .A(G1971), .B(G22), .ZN(n930) );
  XNOR2_X1 U1019 ( .A(G24), .B(G1986), .ZN(n929) );
  NOR2_X1 U1020 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1021 ( .A(G1976), .B(G23), .Z(n931) );
  NAND2_X1 U1022 ( .A1(n932), .A2(n931), .ZN(n934) );
  XOR2_X1 U1023 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n933) );
  XNOR2_X1 U1024 ( .A(n934), .B(n933), .ZN(n939) );
  XOR2_X1 U1025 ( .A(n935), .B(G5), .Z(n937) );
  XNOR2_X1 U1026 ( .A(G21), .B(G1966), .ZN(n936) );
  NOR2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1028 ( .A1(n939), .A2(n938), .ZN(n949) );
  XOR2_X1 U1029 ( .A(G19), .B(G1341), .Z(n943) );
  XNOR2_X1 U1030 ( .A(G1956), .B(G20), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(G1981), .B(G6), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1034 ( .A(KEYINPUT59), .B(G1348), .Z(n944) );
  XNOR2_X1 U1035 ( .A(G4), .B(n944), .ZN(n945) );
  NOR2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1037 ( .A(KEYINPUT60), .B(n947), .Z(n948) );
  NOR2_X1 U1038 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1039 ( .A(KEYINPUT61), .B(n950), .ZN(n951) );
  NAND2_X1 U1040 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1041 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1042 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1043 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1044 ( .A(KEYINPUT62), .B(n959), .Z(G311) );
  XNOR2_X1 U1045 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1046 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1047 ( .A1(n961), .A2(n960), .ZN(G325) );
  INV_X1 U1048 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1049 ( .A(n962), .B(KEYINPUT114), .ZN(n965) );
  XOR2_X1 U1050 ( .A(G301), .B(n963), .Z(n964) );
  XNOR2_X1 U1051 ( .A(n965), .B(n964), .ZN(n968) );
  XNOR2_X1 U1052 ( .A(G286), .B(n966), .ZN(n967) );
  XNOR2_X1 U1053 ( .A(n968), .B(n967), .ZN(n969) );
  NOR2_X1 U1054 ( .A1(G37), .A2(n969), .ZN(n970) );
  XOR2_X1 U1055 ( .A(KEYINPUT115), .B(n970), .Z(G397) );
  XNOR2_X1 U1056 ( .A(G2078), .B(G2072), .ZN(n971) );
  XNOR2_X1 U1057 ( .A(n971), .B(G2100), .ZN(n981) );
  XOR2_X1 U1058 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n973) );
  XNOR2_X1 U1059 ( .A(G2678), .B(KEYINPUT105), .ZN(n972) );
  XNOR2_X1 U1060 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1061 ( .A(KEYINPUT103), .B(G2096), .Z(n975) );
  XNOR2_X1 U1062 ( .A(G2090), .B(KEYINPUT43), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(n975), .B(n974), .ZN(n976) );
  XOR2_X1 U1064 ( .A(n977), .B(n976), .Z(n979) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G2084), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(n979), .B(n978), .ZN(n980) );
  XNOR2_X1 U1067 ( .A(n981), .B(n980), .ZN(G227) );
  XOR2_X1 U1068 ( .A(G1986), .B(G1976), .Z(n983) );
  XNOR2_X1 U1069 ( .A(G1961), .B(G1996), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(n983), .B(n982), .ZN(n984) );
  XOR2_X1 U1071 ( .A(n984), .B(KEYINPUT109), .Z(n986) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G1981), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(n986), .B(n985), .ZN(n994) );
  XOR2_X1 U1074 ( .A(KEYINPUT106), .B(G1991), .Z(n988) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G1956), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(n988), .B(n987), .ZN(n992) );
  XOR2_X1 U1077 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT107), .B(G2474), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n990), .B(n989), .ZN(n991) );
  XOR2_X1 U1080 ( .A(n992), .B(n991), .Z(n993) );
  XNOR2_X1 U1081 ( .A(n994), .B(n993), .ZN(G229) );
  NAND2_X1 U1082 ( .A1(G130), .A2(n995), .ZN(n998) );
  NAND2_X1 U1083 ( .A1(G118), .A2(n996), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n1006) );
  NAND2_X1 U1085 ( .A1(n999), .A2(G142), .ZN(n1000) );
  XOR2_X1 U1086 ( .A(KEYINPUT111), .B(n1000), .Z(n1003) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(G106), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1089 ( .A(n1004), .B(KEYINPUT45), .Z(n1005) );
  NOR2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(n1008), .B(n1007), .ZN(n1013) );
  XNOR2_X1 U1092 ( .A(G162), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XOR2_X1 U1094 ( .A(n1013), .B(n1012), .Z(n1018) );
  XOR2_X1 U1095 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1015) );
  XNOR2_X1 U1096 ( .A(G164), .B(KEYINPUT113), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(n1015), .B(n1014), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(G160), .B(n1016), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(n1018), .B(n1017), .ZN(n1022) );
  XNOR2_X1 U1100 ( .A(n1020), .B(n1019), .ZN(n1021) );
  XNOR2_X1 U1101 ( .A(n1022), .B(n1021), .ZN(n1023) );
  NOR2_X1 U1102 ( .A1(G37), .A2(n1023), .ZN(G395) );
  NOR2_X1 U1103 ( .A1(G401), .A2(n1024), .ZN(n1029) );
  NOR2_X1 U1104 ( .A1(G227), .A2(G229), .ZN(n1026) );
  XNOR2_X1 U1105 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n1025) );
  XNOR2_X1 U1106 ( .A(n1026), .B(n1025), .ZN(n1027) );
  NOR2_X1 U1107 ( .A1(G397), .A2(n1027), .ZN(n1028) );
  NAND2_X1 U1108 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1109 ( .A1(n1030), .A2(G395), .ZN(n1031) );
  XOR2_X1 U1110 ( .A(n1031), .B(KEYINPUT117), .Z(G308) );
  INV_X1 U1111 ( .A(G308), .ZN(G225) );
  INV_X1 U1112 ( .A(G57), .ZN(G237) );
  INV_X1 U1113 ( .A(n1032), .ZN(G223) );
endmodule

