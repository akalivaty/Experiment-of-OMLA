//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT77), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(G148gat), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n210), .A2(new_n212), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G155gat), .B(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n207), .A2(G148gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n218), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT86), .ZN(new_n227));
  XNOR2_X1  g026(.A(G211gat), .B(G218gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G211gat), .A2(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT74), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT22), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n232), .B1(new_n231), .B2(new_n233), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n227), .B(new_n229), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n229), .B1(new_n235), .B2(new_n236), .ZN(new_n238));
  INV_X1    g037(.A(new_n236), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n239), .A2(new_n228), .A3(new_n230), .A4(new_n234), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n226), .B(new_n237), .C1(new_n241), .C2(new_n227), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n225), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n213), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(new_n214), .ZN(new_n246));
  XNOR2_X1  g045(.A(G141gat), .B(G148gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n212), .ZN(new_n250));
  AND2_X1   g049(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n250), .B1(new_n253), .B2(G148gat), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n245), .B1(new_n215), .B2(new_n214), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n249), .B(new_n243), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n241), .B1(new_n226), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G228gat), .ZN(new_n258));
  INV_X1    g057(.A(G233gat), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n244), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n257), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n258), .A2(new_n259), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT3), .B1(new_n241), .B2(new_n226), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n261), .B(new_n262), .C1(new_n225), .C2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n205), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n204), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n238), .A2(KEYINPUT86), .A3(new_n240), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n237), .A2(new_n226), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n243), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n249), .B1(new_n254), .B2(new_n255), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n257), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n264), .B1(new_n272), .B2(new_n262), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G22gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n260), .A2(new_n205), .A3(new_n264), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT87), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n275), .A3(new_n204), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT88), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT88), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n274), .A2(new_n275), .A3(new_n280), .A4(new_n204), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G134gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G127gat), .ZN(new_n284));
  INV_X1    g083(.A(G127gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G134gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(KEYINPUT1), .ZN(new_n289));
  INV_X1    g088(.A(G120gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G113gat), .ZN(new_n291));
  INV_X1    g090(.A(G113gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G120gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT4), .B1(new_n271), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n289), .A2(new_n297), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n225), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT3), .B1(new_n217), .B2(new_n224), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n256), .A3(new_n298), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n225), .A2(new_n300), .A3(KEYINPUT81), .A4(new_n301), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT5), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n304), .A2(new_n306), .A3(new_n307), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT82), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n306), .A2(new_n307), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n304), .A4(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n302), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n308), .A4(new_n306), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n271), .A2(new_n298), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n210), .A2(new_n212), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n216), .A2(new_n213), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(new_n249), .B1(new_n297), .B2(new_n289), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n309), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n298), .B1(new_n217), .B2(new_n224), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n323), .A2(new_n297), .A3(new_n289), .A4(new_n249), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n308), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n319), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n308), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n318), .B1(new_n335), .B2(new_n317), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n312), .B(new_n316), .C1(new_n333), .C2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G1gat), .B(G29gat), .Z(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n337), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT85), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n337), .A2(KEYINPUT85), .A3(new_n343), .A4(new_n345), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n299), .A2(new_n302), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT78), .B1(new_n351), .B2(new_n334), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(new_n319), .A3(new_n326), .A4(new_n332), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n353), .A2(new_n342), .A3(new_n312), .A4(new_n316), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n344), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT84), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n343), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(KEYINPUT84), .A3(new_n344), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n241), .ZN(new_n362));
  INV_X1    g161(.A(G226gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(new_n259), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365));
  INV_X1    g164(.A(G169gat), .ZN(new_n366));
  INV_X1    g165(.A(G176gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(KEYINPUT66), .B2(KEYINPUT23), .ZN(new_n370));
  AND2_X1   g169(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n367), .A2(KEYINPUT23), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT24), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT24), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(G183gat), .A3(G190gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT64), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n372), .B(new_n376), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n382), .A2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n365), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT67), .B(new_n365), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n379), .A2(new_n381), .ZN(new_n390));
  XOR2_X1   g189(.A(KEYINPUT68), .B(G190gat), .Z(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(G183gat), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n365), .B1(new_n373), .B2(new_n366), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n372), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n388), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT27), .B(G183gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT69), .B1(new_n397), .B2(new_n391), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT28), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT26), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n378), .B1(new_n368), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT26), .B1(new_n366), .B2(new_n367), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n369), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n398), .B2(new_n399), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n364), .B1(new_n408), .B2(new_n226), .ZN(new_n409));
  INV_X1    g208(.A(new_n394), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n386), .B2(new_n387), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n411), .B2(new_n389), .ZN(new_n412));
  INV_X1    g211(.A(new_n364), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n362), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n412), .B2(KEYINPUT29), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n408), .A2(new_n364), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n241), .ZN(new_n418));
  XOR2_X1   g217(.A(G8gat), .B(G36gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT75), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n422), .ZN(new_n426));
  INV_X1    g225(.A(new_n418), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n241), .B1(new_n416), .B2(new_n417), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n415), .A2(KEYINPUT30), .A3(new_n418), .A4(new_n422), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n282), .B1(new_n361), .B2(new_n432), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n298), .B(new_n406), .C1(new_n411), .C2(new_n389), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n300), .B1(new_n395), .B2(new_n407), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT70), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT70), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT34), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n434), .A2(new_n435), .ZN(new_n441));
  INV_X1    g240(.A(new_n437), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(KEYINPUT34), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT71), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n442), .A2(KEYINPUT34), .ZN(new_n446));
  NOR4_X1   g245(.A1(new_n434), .A2(new_n435), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n442), .B1(new_n434), .B2(new_n435), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT32), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G15gat), .B(G43gat), .Z(new_n454));
  XNOR2_X1  g253(.A(G71gat), .B(G99gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n456), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n450), .B(KEYINPUT32), .C1(new_n452), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n449), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n440), .A2(new_n448), .A3(new_n457), .A4(new_n459), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(KEYINPUT73), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT73), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n461), .A2(KEYINPUT36), .A3(new_n462), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n433), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n470));
  INV_X1    g269(.A(new_n304), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n309), .B1(new_n471), .B2(new_n313), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n328), .A2(new_n329), .A3(new_n308), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT39), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(new_n309), .C1(new_n471), .C2(new_n313), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(new_n477), .A3(new_n342), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n476), .B2(new_n342), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n474), .B(KEYINPUT40), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n358), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n342), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT89), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n476), .A2(new_n477), .A3(new_n342), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT40), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n470), .B1(new_n431), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n241), .B1(new_n412), .B2(new_n413), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n409), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n426), .B1(new_n491), .B2(new_n428), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n489), .B1(new_n415), .B2(new_n418), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT91), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(KEYINPUT38), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n348), .A2(new_n349), .A3(new_n423), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n312), .A2(new_n316), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n342), .B1(new_n500), .B2(new_n353), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT90), .B1(new_n355), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n358), .A2(new_n503), .A3(new_n344), .A4(new_n354), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n422), .A2(KEYINPUT38), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n491), .B2(new_n428), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(new_n493), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n499), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n488), .B1(new_n498), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT92), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n488), .B(new_n512), .C1(new_n498), .C2(new_n509), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n469), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n463), .A2(new_n465), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n505), .A2(new_n350), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n470), .A2(new_n431), .A3(KEYINPUT35), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n361), .A2(new_n432), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n461), .A2(new_n462), .A3(new_n282), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT35), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n514), .A2(KEYINPUT93), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT93), .B1(new_n514), .B2(new_n522), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT14), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G29gat), .A2(G36gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT94), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(KEYINPUT15), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(KEYINPUT96), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n537), .A2(new_n533), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n536), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(G1gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(G1gat), .B2(new_n548), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G8gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(KEYINPUT17), .B(new_n536), .C1(new_n541), .C2(new_n544), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n545), .A2(new_n552), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT97), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n545), .B(new_n552), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n556), .B(KEYINPUT13), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n560), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G197gat), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT11), .B(G169gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT12), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n562), .A2(new_n572), .A3(new_n565), .A4(new_n566), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G57gat), .B(G64gat), .Z(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  INV_X1    g377(.A(G71gat), .ZN(new_n579));
  INV_X1    g378(.A(G78gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n285), .ZN(new_n589));
  INV_X1    g388(.A(new_n583), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n582), .B(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n552), .B1(KEYINPUT21), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n588), .B(G127gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  INV_X1    g396(.A(G155gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT98), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n599), .B(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n593), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n593), .B2(new_n596), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT99), .ZN(new_n608));
  XNOR2_X1  g407(.A(G190gat), .B(G218gat), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n608), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G99gat), .B(G106gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n616), .A2(new_n624), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n547), .A2(new_n554), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n545), .A2(new_n628), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n609), .A2(new_n610), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n630), .B2(new_n633), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n613), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n630), .A2(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n631), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n612), .A3(new_n634), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G230gat), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n259), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n584), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n591), .A2(new_n625), .A3(new_n623), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n650), .B2(new_n643), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  OR2_X1    g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n647), .A2(new_n648), .ZN(new_n656));
  INV_X1    g455(.A(new_n643), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n650), .A2(new_n643), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n605), .A2(new_n641), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n525), .A2(new_n576), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n361), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(G1gat), .Z(G1324gat));
  OAI21_X1  g466(.A(G8gat), .B1(new_n665), .B2(new_n432), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT102), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n665), .A2(new_n432), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  NOR4_X1   g474(.A1(new_n665), .A2(KEYINPUT42), .A3(new_n432), .A4(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n669), .B(new_n670), .C1(new_n674), .C2(new_n676), .ZN(G1325gat));
  NAND2_X1  g476(.A1(new_n467), .A2(new_n468), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n665), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n515), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n665), .B2(new_n681), .ZN(G1326gat));
  NOR2_X1   g481(.A1(new_n665), .A2(new_n282), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT43), .B(G22gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1327gat));
  INV_X1    g484(.A(new_n605), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n662), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n641), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n525), .A2(new_n576), .A3(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(G29gat), .A3(new_n361), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n641), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n523), .B2(new_n524), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n514), .A2(new_n522), .ZN(new_n695));
  INV_X1    g494(.A(new_n641), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n692), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n361), .ZN(new_n700));
  INV_X1    g499(.A(new_n576), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n687), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G29gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n691), .A2(new_n704), .A3(new_n705), .ZN(G1328gat));
  NOR3_X1   g505(.A1(new_n689), .A2(G36gat), .A3(new_n432), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n699), .A2(new_n431), .A3(new_n702), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G36gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n708), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(G1329gat));
  INV_X1    g512(.A(new_n678), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n699), .A2(G43gat), .A3(new_n714), .A4(new_n702), .ZN(new_n715));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n689), .B2(new_n680), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  NAND4_X1  g522(.A1(new_n699), .A2(G50gat), .A3(new_n470), .A4(new_n702), .ZN(new_n724));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n689), .B2(new_n282), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT48), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n724), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1331gat));
  NOR4_X1   g530(.A1(new_n686), .A2(new_n576), .A3(new_n696), .A4(new_n662), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n695), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n361), .ZN(new_n734));
  XNOR2_X1  g533(.A(KEYINPUT104), .B(G57gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1332gat));
  XNOR2_X1  g535(.A(new_n733), .B(KEYINPUT105), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n431), .B(KEYINPUT106), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n737), .B2(new_n678), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n695), .A2(new_n515), .A3(new_n732), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n579), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1334gat));
  NOR2_X1   g550(.A1(new_n737), .A2(new_n282), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n580), .ZN(G1335gat));
  NOR3_X1   g552(.A1(new_n605), .A2(new_n576), .A3(new_n662), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n699), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n361), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n605), .A2(new_n576), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n695), .A2(new_n696), .A3(new_n757), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n758), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n758), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n700), .A2(new_n618), .A3(new_n661), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n756), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  NAND2_X1  g567(.A1(new_n758), .A2(KEYINPUT109), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n762), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n758), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n738), .A2(G92gat), .A3(new_n662), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT110), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n770), .A2(new_n775), .A3(new_n771), .A4(new_n772), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n694), .A2(new_n431), .A3(new_n698), .A4(new_n754), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G92gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT52), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(new_n765), .B2(new_n772), .ZN(new_n781));
  OAI21_X1  g580(.A(G92gat), .B1(new_n755), .B2(new_n738), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n755), .B2(new_n678), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n680), .A2(G99gat), .A3(new_n662), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT111), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n766), .B2(new_n787), .ZN(G1338gat));
  NOR3_X1   g587(.A1(new_n282), .A2(new_n662), .A3(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n765), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n694), .A2(new_n470), .A3(new_n698), .A4(new_n754), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT112), .B1(new_n792), .B2(G106gat), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n770), .A2(new_n771), .A3(new_n789), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n798), .B2(new_n791), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n663), .A2(new_n576), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n647), .A2(new_n648), .A3(new_n643), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n654), .B1(new_n649), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n576), .A2(new_n660), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n563), .A2(new_n564), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n571), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n575), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n661), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n641), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n807), .A2(new_n660), .A3(new_n808), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n818), .A2(new_n641), .A3(new_n819), .A4(new_n813), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n696), .A3(new_n814), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n819), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n817), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n800), .B1(new_n825), .B2(new_n686), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n361), .A3(new_n520), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n738), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n576), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n738), .A2(new_n700), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n826), .A2(new_n470), .A3(new_n680), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n701), .A2(new_n292), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(G1340gat));
  AOI21_X1  g633(.A(G120gat), .B1(new_n829), .B2(new_n661), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n662), .A2(new_n290), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n832), .B2(new_n836), .ZN(G1341gat));
  NAND3_X1  g636(.A1(new_n829), .A2(new_n285), .A3(new_n605), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n832), .A2(new_n605), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n285), .B2(new_n839), .ZN(G1342gat));
  NAND2_X1  g639(.A1(new_n432), .A2(new_n696), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(G134gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT114), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT114), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT115), .Z(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n844), .B2(new_n846), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n283), .B1(new_n832), .B2(new_n696), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(new_n854), .ZN(G1343gat));
  NOR2_X1   g654(.A1(new_n826), .A2(new_n282), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n826), .B2(new_n282), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n714), .A2(new_n831), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n858), .A2(new_n861), .A3(new_n576), .A4(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n253), .ZN(new_n864));
  INV_X1    g663(.A(new_n826), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n865), .A2(new_n700), .A3(new_n470), .A4(new_n678), .ZN(new_n866));
  INV_X1    g665(.A(new_n738), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n701), .A2(G141gat), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n863), .A2(new_n864), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n872), .B(new_n873), .Z(G1344gat));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n858), .A2(new_n861), .A3(new_n661), .A4(new_n862), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(G148gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n818), .A2(new_n641), .A3(new_n813), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT113), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n820), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n605), .B1(new_n881), .B2(new_n817), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n470), .B(new_n860), .C1(new_n882), .C2(new_n800), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n696), .B1(new_n809), .B2(new_n815), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n686), .B1(new_n885), .B2(new_n879), .ZN(new_n886));
  INV_X1    g685(.A(new_n800), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n282), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n884), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n822), .A2(new_n576), .B1(new_n814), .B2(new_n661), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n823), .B1(new_n890), .B2(new_n696), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n800), .B1(new_n891), .B2(new_n686), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT119), .B(new_n857), .C1(new_n892), .C2(new_n282), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n883), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n714), .A2(new_n662), .A3(new_n831), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(KEYINPUT120), .A3(new_n895), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(G148gat), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n878), .B1(new_n900), .B2(KEYINPUT59), .ZN(new_n901));
  NOR4_X1   g700(.A1(new_n866), .A2(G148gat), .A3(new_n662), .A4(new_n867), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n875), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(G148gat), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT120), .B1(new_n894), .B2(new_n895), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT59), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n878), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n902), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n903), .A2(new_n910), .ZN(G1345gat));
  NAND3_X1  g710(.A1(new_n868), .A2(new_n598), .A3(new_n605), .ZN(new_n912));
  INV_X1    g711(.A(new_n858), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n861), .A2(new_n862), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n686), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n598), .ZN(G1346gat));
  OR3_X1    g715(.A1(new_n866), .A2(G162gat), .A3(new_n841), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n913), .A2(new_n914), .A3(new_n641), .ZN(new_n918));
  INV_X1    g717(.A(G162gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(G1347gat));
  NOR3_X1   g719(.A1(new_n826), .A2(new_n470), .A3(new_n680), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n361), .A2(new_n431), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT122), .Z(new_n923));
  AND2_X1   g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n366), .B1(new_n924), .B2(new_n576), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT123), .ZN(new_n926));
  NOR4_X1   g725(.A1(new_n826), .A2(new_n700), .A3(new_n520), .A4(new_n738), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(new_n576), .A3(new_n374), .A4(new_n375), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1348gat));
  INV_X1    g728(.A(new_n924), .ZN(new_n930));
  OAI21_X1  g729(.A(G176gat), .B1(new_n930), .B2(new_n662), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n367), .A3(new_n661), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n930), .B2(new_n686), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n686), .A2(new_n397), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n927), .A2(new_n935), .B1(new_n936), .B2(KEYINPUT60), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(KEYINPUT60), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n938), .B(new_n939), .Z(G1350gat));
  NOR2_X1   g739(.A1(new_n641), .A2(new_n391), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n927), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(G190gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n943), .B1(new_n924), .B2(new_n696), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n945), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NOR3_X1   g750(.A1(new_n826), .A2(new_n700), .A3(new_n738), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n470), .A3(new_n678), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n576), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n923), .A2(new_n678), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT126), .Z(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n894), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n576), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n661), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G204gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n953), .A2(G204gat), .A3(new_n662), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1353gat));
  NAND2_X1  g764(.A1(new_n958), .A2(new_n605), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G211gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT63), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n969), .A3(G211gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n953), .A2(G211gat), .A3(new_n686), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT127), .Z(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n954), .A2(new_n974), .A3(new_n696), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n958), .A2(new_n696), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n974), .ZN(G1355gat));
endmodule


