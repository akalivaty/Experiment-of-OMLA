//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n203), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n202), .C2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n206), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n206), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n218), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n217), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT66), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  NOR2_X1   g0046(.A1(new_n213), .A2(KEYINPUT8), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  MUX2_X1   g0048(.A(new_n247), .B(new_n248), .S(KEYINPUT67), .Z(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n221), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n250), .B2(G20), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n252), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  MUX2_X1   g0056(.A(G223), .B(G226), .S(G1698), .Z(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT71), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT71), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n261), .A3(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n257), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G87), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT75), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G190), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(G232), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n267), .A2(KEYINPUT75), .A3(new_n268), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n271), .A2(new_n272), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(G200), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n285));
  INV_X1    g0085(.A(G68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n258), .A2(G33), .ZN(new_n287));
  AOI21_X1  g0087(.A(G20), .B1(new_n264), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT73), .B1(new_n288), .B2(KEYINPUT7), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT73), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT7), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n290), .B(new_n291), .C1(new_n292), .C2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT71), .B(KEYINPUT3), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n287), .B1(new_n295), .B2(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n291), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n286), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(G58), .B(G68), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n300), .A2(G20), .B1(G159), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n285), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(G20), .B1(new_n262), .B2(new_n264), .ZN(new_n305));
  OAI21_X1  g0105(.A(G68), .B1(new_n305), .B2(new_n291), .ZN(new_n306));
  AOI211_X1 g0106(.A(KEYINPUT7), .B(G20), .C1(new_n262), .C2(new_n264), .ZN(new_n307));
  OAI211_X1 g0107(.A(KEYINPUT16), .B(new_n302), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n304), .A2(KEYINPUT74), .A3(new_n254), .A4(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n308), .A2(new_n254), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT74), .B1(new_n311), .B2(new_n304), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n256), .B(new_n284), .C1(new_n310), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT17), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n256), .B1(new_n310), .B2(new_n312), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT18), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n271), .A2(new_n318), .A3(new_n278), .A4(new_n279), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT76), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n281), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n320), .B1(new_n319), .B2(new_n322), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n316), .A2(new_n317), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n256), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT74), .ZN(new_n329));
  INV_X1    g0129(.A(new_n285), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n264), .A2(new_n287), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n222), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n290), .B1(new_n332), .B2(new_n291), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n288), .A2(KEYINPUT73), .A3(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n298), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G68), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n330), .B1(new_n336), .B2(new_n302), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n308), .A2(new_n254), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n329), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n328), .B1(new_n339), .B2(new_n309), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n319), .A2(new_n322), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT76), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n323), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT18), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(KEYINPUT17), .A3(new_n284), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n315), .A2(new_n327), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n277), .A2(G238), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n268), .A2(new_n273), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n276), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n268), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n214), .A2(G1698), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n292), .B(new_n353), .C1(G226), .C2(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT13), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n355), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n268), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n275), .B1(G238), .B2(new_n277), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n321), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n357), .A2(new_n362), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n363), .A2(new_n364), .B1(new_n365), .B2(new_n318), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n363), .A2(new_n364), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT70), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT70), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n363), .A2(new_n369), .A3(new_n364), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n366), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n251), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n286), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT12), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n263), .A2(G20), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(G77), .B1(G20), .B2(new_n286), .ZN(new_n376));
  INV_X1    g0176(.A(G50), .ZN(new_n377));
  INV_X1    g0177(.A(new_n301), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n380));
  INV_X1    g0180(.A(new_n255), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n374), .B(new_n380), .C1(new_n286), .C2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT11), .B1(new_n379), .B2(new_n254), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n371), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n365), .B2(new_n272), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n282), .B1(new_n357), .B2(new_n362), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n372), .A2(new_n377), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n381), .B2(new_n377), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n377), .A2(new_n213), .A3(new_n286), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(G20), .B1(G150), .B2(new_n301), .ZN(new_n393));
  INV_X1    g0193(.A(new_n375), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n249), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(new_n254), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G222), .A2(G1698), .ZN(new_n397));
  INV_X1    g0197(.A(G1698), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(G223), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n292), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(new_n268), .C1(G77), .C2(new_n292), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n277), .A2(G226), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n350), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(G179), .ZN(new_n404));
  AOI211_X1 g0204(.A(new_n396), .B(new_n404), .C1(new_n321), .C2(new_n403), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n396), .A2(KEYINPUT9), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT69), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(G200), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n408), .B1(new_n272), .B2(new_n403), .C1(new_n396), .C2(KEYINPUT9), .ZN(new_n409));
  OR3_X1    g0209(.A1(new_n407), .A2(KEYINPUT10), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT10), .B1(new_n407), .B2(new_n409), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n405), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n268), .A2(new_n276), .A3(new_n209), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n292), .A2(G232), .A3(new_n398), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n292), .A2(G238), .A3(G1698), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(new_n203), .C2(new_n292), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n275), .B(new_n413), .C1(new_n416), .C2(new_n268), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT68), .A3(G190), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT15), .B(G87), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n419), .A2(new_n394), .B1(new_n222), .B2(new_n208), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n248), .A2(new_n378), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n254), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n251), .A2(G77), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n255), .B2(G77), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n418), .B(new_n426), .C1(new_n282), .C2(new_n417), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT68), .B1(new_n417), .B2(G190), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n417), .A2(new_n318), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n425), .C1(G169), .C2(new_n417), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n347), .A2(new_n389), .A3(new_n412), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G45), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G1), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(G250), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n273), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n352), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n264), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n295), .B2(G33), .ZN(new_n440));
  NOR2_X1   g0240(.A1(G238), .A2(G1698), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n209), .B2(G1698), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n440), .A2(new_n442), .B1(G33), .B2(G116), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n318), .B(new_n438), .C1(new_n443), .C2(new_n352), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n262), .A3(new_n264), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G116), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n352), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n438), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n321), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n449), .A3(KEYINPUT80), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n447), .A2(new_n448), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT80), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n318), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NOR4_X1   g0254(.A1(KEYINPUT81), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G87), .A2(G97), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n203), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT19), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n222), .B1(new_n355), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n262), .A2(new_n264), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n222), .A2(G68), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n459), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n222), .A2(G33), .A3(G97), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n460), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT82), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n254), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n419), .A2(new_n372), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n250), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n251), .A2(new_n471), .A3(new_n221), .A4(new_n253), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n419), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT83), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n469), .A2(new_n478), .A3(new_n470), .A4(new_n475), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n454), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(G200), .B1(new_n447), .B2(new_n448), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n438), .B1(new_n443), .B2(new_n352), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n272), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n473), .A2(G87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n469), .A2(new_n484), .A3(new_n470), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT84), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n480), .A2(KEYINPUT84), .A3(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT86), .B1(new_n222), .B2(G107), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT23), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT23), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT86), .B(new_n495), .C1(new_n222), .C2(G107), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n494), .A2(new_n496), .B1(G116), .B2(new_n375), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n222), .A2(G87), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT22), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n262), .A2(new_n500), .A3(new_n264), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n331), .B2(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT24), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n497), .A2(new_n501), .A3(new_n505), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n254), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT25), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n251), .B2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n251), .A2(new_n509), .A3(G107), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n511), .A2(new_n512), .B1(new_n203), .B2(new_n472), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G250), .A2(G1698), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n215), .B2(G1698), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n262), .A3(new_n264), .ZN(new_n517));
  XOR2_X1   g0317(.A(KEYINPUT87), .B(G294), .Z(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G33), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n352), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G41), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n435), .A2(KEYINPUT78), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G41), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n250), .B(G45), .C1(new_n525), .C2(KEYINPUT5), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(KEYINPUT5), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n349), .A2(new_n524), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT78), .B1(new_n435), .B2(new_n523), .ZN(new_n532));
  OAI211_X1 g0332(.A(G264), .B(new_n352), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n521), .A2(G190), .A3(new_n530), .A4(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n440), .A2(new_n516), .B1(G33), .B2(new_n518), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n530), .B(new_n533), .C1(new_n535), .C2(new_n352), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n508), .A2(new_n514), .A3(new_n534), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n321), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n521), .A2(new_n318), .A3(new_n530), .A4(new_n533), .ZN(new_n540));
  INV_X1    g0340(.A(new_n254), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n504), .B2(new_n506), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n540), .C1(new_n542), .C2(new_n513), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G270), .B(new_n352), .C1(new_n531), .C2(new_n532), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n292), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G257), .A2(G1698), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n210), .B2(G1698), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n548), .B1(new_n440), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n546), .B(new_n530), .C1(new_n551), .C2(new_n352), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n251), .A2(new_n471), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT85), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n541), .A4(G116), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT85), .B1(new_n472), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G283), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n559), .B(new_n222), .C1(G33), .C2(new_n202), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n556), .A2(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n254), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n560), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n372), .A2(new_n556), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n558), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n552), .A2(new_n568), .A3(KEYINPUT21), .A4(G169), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n552), .A2(new_n568), .A3(G169), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n552), .A2(G200), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n550), .A2(new_n262), .A3(new_n264), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n547), .B2(new_n292), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n268), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(G190), .A3(new_n546), .A4(new_n530), .ZN(new_n577));
  INV_X1    g0377(.A(new_n568), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n552), .A2(new_n318), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n568), .ZN(new_n581));
  AND4_X1   g0381(.A1(new_n569), .A2(new_n572), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n203), .B1(new_n294), .B2(new_n298), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G97), .A2(G107), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT6), .B1(new_n204), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n203), .A2(KEYINPUT6), .A3(G97), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n587), .A2(new_n222), .B1(new_n208), .B2(new_n378), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n254), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n372), .A2(new_n202), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT77), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(G97), .B2(new_n473), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(new_n352), .C1(new_n531), .C2(new_n532), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n594), .A2(new_n530), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n209), .A2(G1698), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT4), .B1(new_n440), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n209), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n292), .A2(new_n398), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n601), .A3(new_n559), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n268), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n595), .A2(new_n603), .A3(new_n318), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(new_n603), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n321), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT79), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n595), .A2(new_n603), .A3(new_n608), .A4(new_n318), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n593), .A2(new_n605), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n598), .A2(new_n601), .A3(new_n559), .ZN(new_n611));
  INV_X1    g0411(.A(new_n596), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n599), .B1(new_n463), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n352), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n594), .A2(new_n530), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G190), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(G200), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n589), .A4(new_n592), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n545), .A2(new_n582), .A3(new_n610), .A4(new_n619), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n433), .A2(new_n492), .A3(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n385), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n388), .B2(new_n431), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n623), .A2(new_n315), .A3(new_n345), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n327), .A2(new_n344), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n410), .A2(new_n411), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n405), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n542), .A2(new_n513), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n537), .A2(new_n534), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n486), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n543), .A2(new_n569), .A3(new_n572), .A4(new_n581), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(new_n610), .A4(new_n619), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n476), .A2(new_n444), .A3(new_n449), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n610), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n490), .A2(KEYINPUT26), .A3(new_n491), .A4(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n487), .A2(new_n635), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(new_n610), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n636), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n629), .B1(new_n433), .B2(new_n642), .ZN(G369));
  NAND3_X1  g0443(.A1(new_n250), .A2(new_n222), .A3(G13), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G343), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT88), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n543), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n649), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n538), .B1(new_n630), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n543), .ZN(new_n653));
  INV_X1    g0453(.A(new_n650), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT89), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n572), .A2(new_n581), .A3(new_n569), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n651), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n650), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n651), .A2(new_n578), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n658), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n572), .A2(new_n579), .A3(new_n581), .A4(new_n569), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n660), .A2(new_n667), .ZN(G399));
  NAND2_X1  g0468(.A1(new_n459), .A2(new_n556), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n225), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(G1), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n220), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT29), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT91), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n638), .A2(new_n641), .ZN(new_n680));
  INV_X1    g0480(.A(new_n636), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n679), .B1(new_n682), .B2(new_n651), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n642), .A2(KEYINPUT91), .A3(new_n649), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n678), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT92), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT92), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n687), .B(new_n678), .C1(new_n683), .C2(new_n684), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n480), .A2(KEYINPUT84), .A3(new_n487), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT84), .B1(new_n480), .B2(new_n487), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n639), .A3(new_n637), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT26), .B1(new_n640), .B2(new_n610), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n634), .A2(new_n693), .A3(new_n635), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n649), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n686), .A2(new_n688), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n552), .A2(new_n482), .A3(new_n318), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT90), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n606), .A4(new_n536), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  INV_X1    g0502(.A(new_n533), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n520), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(new_n603), .A3(new_n451), .A4(new_n595), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n576), .A2(G179), .A3(new_n546), .A4(new_n530), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n482), .A2(new_n703), .A3(new_n520), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n580), .A3(KEYINPUT30), .A4(new_n616), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n536), .B1(new_n614), .B2(new_n615), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n552), .A2(new_n482), .A3(new_n318), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT90), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n701), .A2(new_n707), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT31), .B1(new_n713), .B2(new_n649), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n707), .B(new_n709), .C1(new_n711), .C2(new_n710), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n649), .A2(KEYINPUT31), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n610), .A2(new_n619), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(new_n663), .A3(new_n544), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n691), .A2(new_n719), .A3(new_n651), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n698), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n697), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n677), .B1(new_n724), .B2(G1), .ZN(G364));
  INV_X1    g0525(.A(new_n665), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n222), .A2(G13), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n250), .B1(new_n727), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n672), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(G330), .B2(new_n664), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n671), .A2(new_n331), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G355), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G116), .B2(new_n225), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n440), .A2(new_n671), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n434), .B2(new_n220), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n240), .A2(G45), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(G1), .B(G13), .C1(new_n222), .C2(G169), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT93), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n730), .B1(new_n740), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n222), .A2(G179), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n272), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n203), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n222), .A2(new_n318), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n755), .A2(new_n282), .A3(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n272), .A2(new_n282), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n757), .A2(new_n286), .B1(new_n759), .B2(new_n377), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n753), .B(new_n760), .C1(G77), .C2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n755), .A2(new_n272), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n292), .B1(new_n766), .B2(new_n213), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n272), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n222), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(G97), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n758), .A2(new_n751), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT94), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G87), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n751), .A2(new_n761), .ZN(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n764), .A2(new_n771), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  NOR2_X1   g0583(.A1(new_n757), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G311), .B2(new_n763), .ZN(new_n785));
  INV_X1    g0585(.A(new_n752), .ZN(new_n786));
  INV_X1    g0586(.A(new_n778), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n786), .A2(G283), .B1(new_n787), .B2(G329), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT96), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n770), .A2(new_n518), .ZN(new_n790));
  INV_X1    g0590(.A(new_n759), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n765), .A2(G322), .B1(new_n791), .B2(G326), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n785), .A2(new_n789), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n331), .B1(new_n775), .B2(new_n547), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n782), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n750), .B1(new_n796), .B2(new_n744), .ZN(new_n797));
  INV_X1    g0597(.A(new_n747), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n664), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n732), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  INV_X1    g0601(.A(new_n730), .ZN(new_n802));
  INV_X1    g0602(.A(new_n744), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n746), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT97), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n802), .B1(new_n806), .B2(new_n208), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n765), .A2(G143), .B1(new_n791), .B2(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G150), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n809), .B2(new_n757), .C1(new_n779), .C2(new_n762), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n786), .A2(G68), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n440), .C1(new_n813), .C2(new_n778), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G58), .B2(new_n770), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n811), .B(new_n815), .C1(new_n377), .C2(new_n775), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n786), .A2(G87), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G311), .B2(new_n787), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT98), .Z(new_n819));
  OAI221_X1 g0619(.A(new_n331), .B1(new_n762), .B2(new_n556), .C1(new_n769), .C2(new_n202), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n757), .A2(new_n821), .B1(new_n759), .B2(new_n547), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G294), .C2(new_n765), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n819), .B(new_n823), .C1(new_n203), .C2(new_n775), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n431), .A2(new_n649), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n429), .B1(new_n426), .B2(new_n651), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(new_n431), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n807), .B1(new_n803), .B2(new_n825), .C1(new_n828), .C2(new_n746), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n682), .A2(new_n432), .A3(new_n651), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n683), .A2(new_n684), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n828), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n832), .A2(KEYINPUT99), .A3(new_n722), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n833), .B(new_n802), .C1(new_n722), .C2(new_n832), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT99), .B1(new_n832), .B2(new_n722), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n829), .B1(new_n834), .B2(new_n835), .ZN(G384));
  INV_X1    g0636(.A(new_n587), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(KEYINPUT35), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n838), .A2(G116), .A3(new_n223), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n220), .B(G77), .C1(new_n213), .C2(new_n286), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n377), .A2(G68), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n250), .B(G13), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n433), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n686), .A2(new_n847), .A3(new_n688), .A4(new_n696), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n848), .A2(new_n629), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT103), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT7), .B1(new_n440), .B2(G20), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n305), .A2(new_n291), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n852), .A2(new_n853), .A3(G68), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n330), .B1(new_n854), .B2(new_n302), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n256), .B1(new_n338), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n647), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(KEYINPUT102), .A3(new_n647), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n346), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n342), .A2(new_n323), .A3(new_n856), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n313), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n864), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n316), .A2(new_n326), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n316), .A2(new_n647), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n868), .A4(new_n313), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n862), .A2(new_n870), .A3(KEYINPUT38), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n313), .B1(new_n343), .B2(new_n340), .ZN(new_n872));
  INV_X1    g0672(.A(new_n647), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n340), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n346), .A2(new_n874), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n851), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n862), .A2(new_n870), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n862), .A2(new_n870), .A3(KEYINPUT38), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n622), .A2(new_n649), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n879), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n625), .A2(new_n647), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n883), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n651), .A2(KEYINPUT101), .A3(new_n384), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT101), .ZN(new_n890));
  INV_X1    g0690(.A(new_n384), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n649), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n385), .B2(new_n388), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n893), .B1(new_n387), .B2(new_n386), .C1(new_n371), .C2(new_n384), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n826), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n830), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n887), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n886), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n850), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n828), .A2(new_n895), .A3(new_n896), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT105), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n492), .A2(new_n620), .A3(new_n649), .ZN(new_n905));
  INV_X1    g0705(.A(new_n714), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n904), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n714), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n720), .A2(new_n911), .A3(KEYINPUT105), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n903), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n862), .B2(new_n870), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n871), .B2(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n917), .B(new_n903), .C1(new_n909), .C2(new_n912), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n876), .A2(new_n877), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n881), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n883), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n915), .A2(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n909), .A2(new_n912), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n922), .A2(new_n847), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n847), .B2(new_n923), .ZN(new_n925));
  OR3_X1    g0725(.A1(new_n924), .A2(new_n925), .A3(new_n698), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n902), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n250), .B2(new_n727), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n902), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n846), .B1(new_n928), .B2(new_n929), .ZN(G367));
  NAND2_X1  g0730(.A1(new_n637), .A2(new_n649), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n593), .A2(new_n649), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n610), .A2(new_n619), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n666), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n936));
  INV_X1    g0736(.A(new_n543), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n619), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n649), .B1(new_n938), .B2(new_n610), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n657), .A2(new_n659), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n934), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n939), .B1(new_n942), .B2(KEYINPUT42), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(KEYINPUT42), .B2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n649), .A2(new_n485), .ZN(new_n945));
  MUX2_X1   g0745(.A(new_n635), .B(new_n640), .S(new_n945), .Z(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT106), .Z(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n944), .B2(new_n949), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n936), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  INV_X1    g0753(.A(new_n936), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n672), .B(KEYINPUT41), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n657), .A2(new_n659), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n941), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(new_n665), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n724), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT108), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n724), .A2(KEYINPUT108), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n660), .A2(new_n934), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT45), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n660), .A2(new_n968), .A3(new_n934), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n660), .B2(new_n934), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n967), .A2(new_n971), .A3(new_n667), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n667), .B1(new_n967), .B2(new_n971), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n963), .A2(new_n964), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n957), .B1(new_n975), .B2(new_n724), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n952), .B(new_n956), .C1(new_n976), .C2(new_n729), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n748), .B1(new_n225), .B2(new_n419), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n737), .A2(new_n236), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n730), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n757), .A2(new_n779), .B1(new_n762), .B2(new_n377), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G137), .B2(new_n787), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n791), .A2(G143), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n766), .B2(new_n809), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n752), .A2(new_n208), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n984), .A2(new_n331), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n770), .A2(G68), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n776), .A2(G58), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n982), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n752), .A2(new_n202), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n766), .A2(new_n547), .B1(new_n778), .B2(new_n991), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(G311), .C2(new_n791), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n770), .A2(G107), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n756), .A2(new_n518), .B1(G283), .B2(new_n763), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n993), .A2(new_n463), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n775), .A2(new_n556), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n989), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT47), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n803), .B1(new_n999), .B2(new_n1000), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n980), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n947), .B2(new_n798), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n977), .A2(new_n1004), .ZN(G387));
  NAND2_X1  g0805(.A1(new_n656), .A2(new_n747), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n248), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g0808(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT109), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1008), .B(new_n1009), .C1(new_n1010), .C2(new_n669), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n670), .A2(KEYINPUT109), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n736), .B1(new_n233), .B2(new_n434), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n669), .A2(new_n733), .B1(new_n203), .B2(new_n671), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(KEYINPUT110), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n748), .ZN(new_n1016));
  AOI21_X1  g0816(.A(KEYINPUT110), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n730), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n766), .A2(new_n991), .B1(new_n762), .B2(new_n547), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT112), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(KEYINPUT112), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n756), .A2(G311), .B1(new_n791), .B2(G322), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n776), .A2(new_n518), .B1(G283), .B2(new_n770), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n786), .A2(G116), .B1(new_n787), .B2(G326), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1030), .A2(new_n463), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G159), .A2(new_n791), .B1(new_n763), .B2(G68), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n809), .B2(new_n778), .C1(new_n249), .C2(new_n757), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n775), .A2(new_n208), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n440), .B1(new_n202), .B2(new_n752), .C1(new_n766), .C2(new_n377), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n769), .A2(new_n419), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT111), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1033), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1018), .B1(new_n1041), .B2(new_n744), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n960), .A2(new_n729), .B1(new_n1006), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n961), .A2(new_n672), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n724), .A2(new_n960), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(G393));
  NOR2_X1   g0846(.A1(new_n245), .A2(new_n737), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n748), .B1(new_n202), .B2(new_n225), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n730), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n765), .A2(G311), .B1(new_n791), .B2(G317), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n787), .A2(G322), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n757), .B2(new_n547), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G294), .B2(new_n763), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n776), .A2(G283), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n292), .B(new_n753), .C1(G116), .C2(new_n770), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n765), .A2(G159), .B1(new_n791), .B2(G150), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT51), .Z(new_n1060));
  AOI211_X1 g0860(.A(new_n463), .B(new_n817), .C1(G143), .C2(new_n787), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n286), .C2(new_n775), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n770), .A2(G77), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n248), .B2(new_n762), .C1(new_n757), .C2(new_n377), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT113), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1058), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1049), .B1(new_n1066), .B2(new_n744), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n934), .B2(new_n798), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n974), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n728), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n673), .B1(new_n1069), .B2(new_n961), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n975), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  AOI21_X1  g0873(.A(new_n698), .B1(new_n909), .B2(new_n912), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n847), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n895), .A2(new_n896), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n721), .B2(new_n828), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n828), .A2(new_n895), .A3(new_n896), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1077), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n642), .A2(new_n649), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n826), .B1(new_n1080), .B2(new_n432), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1076), .B1(new_n1074), .B2(new_n828), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n827), .A2(new_n431), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n826), .B1(new_n695), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n721), .A2(new_n1076), .A3(new_n828), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1079), .A2(new_n1081), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n849), .A2(new_n1075), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n885), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1081), .B2(new_n897), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT39), .B1(new_n920), .B2(new_n883), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n871), .A2(new_n914), .A3(new_n851), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n885), .B1(new_n920), .B2(new_n883), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n695), .A2(new_n1084), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1076), .B1(new_n1096), .B2(new_n826), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1098), .A3(new_n1086), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1099), .B1(new_n1101), .B2(KEYINPUT115), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1100), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n830), .A2(new_n898), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1076), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n879), .A2(new_n884), .B1(new_n1105), .B2(new_n1090), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1107));
  OAI211_X1 g0907(.A(KEYINPUT115), .B(new_n1103), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1089), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1110));
  AND4_X1   g0910(.A1(new_n629), .A2(new_n1088), .A3(new_n848), .A4(new_n1075), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT115), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n879), .A2(new_n884), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1113), .A2(new_n1091), .B1(new_n1097), .B2(new_n1095), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1114), .B2(new_n1100), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1111), .A2(new_n1108), .A3(new_n1099), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1110), .A2(new_n672), .A3(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1115), .A2(new_n1108), .A3(new_n729), .A4(new_n1099), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1113), .A2(new_n745), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n756), .A2(G137), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT54), .B(G143), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1120), .B1(new_n762), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1122), .A2(KEYINPUT116), .B1(G159), .B2(new_n770), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(KEYINPUT116), .B2(new_n1122), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT117), .Z(new_n1125));
  NAND2_X1  g0925(.A1(new_n776), .A2(G150), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n765), .A2(G132), .B1(new_n791), .B2(G128), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n331), .B1(new_n787), .B2(G125), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n377), .C2(new_n752), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G107), .A2(new_n756), .B1(new_n765), .B2(G116), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n777), .B(new_n1132), .C1(new_n202), .C2(new_n762), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n791), .A2(G283), .B1(new_n787), .B2(G294), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1134), .A2(new_n331), .A3(new_n1063), .A4(new_n812), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT118), .Z(new_n1137));
  OAI21_X1  g0937(.A(new_n744), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n802), .B1(new_n806), .B2(new_n249), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1119), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1118), .A2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1117), .A2(KEYINPUT119), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT119), .B1(new_n1117), .B2(new_n1141), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(G378));
  NOR2_X1   g0944(.A1(new_n396), .A2(new_n873), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT55), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n412), .B(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1148));
  XOR2_X1   g0948(.A(new_n1147), .B(new_n1148), .Z(new_n1149));
  OAI211_X1 g0949(.A(new_n913), .B(KEYINPUT40), .C1(new_n871), .C2(new_n878), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n720), .A2(new_n911), .A3(KEYINPUT105), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT105), .B1(new_n720), .B2(new_n911), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1078), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n883), .B2(new_n882), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n916), .ZN(new_n1155));
  OAI211_X1 g0955(.A(G330), .B(new_n1150), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n886), .A3(new_n900), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n901), .A2(G330), .A3(new_n922), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1149), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1149), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n729), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n730), .B1(new_n804), .B2(G50), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n377), .B1(G33), .B2(G41), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n463), .B2(new_n525), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1036), .A2(G41), .A3(new_n440), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n756), .A2(G97), .B1(new_n474), .B2(new_n763), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT120), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n778), .A2(new_n821), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n556), .A2(new_n759), .B1(new_n752), .B2(new_n213), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(G107), .C2(new_n765), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1166), .A2(new_n987), .A3(new_n1168), .A4(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT58), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1165), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1121), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n776), .A2(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(KEYINPUT121), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G125), .A2(new_n791), .B1(new_n763), .B2(G137), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n765), .A2(G128), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n813), .C2(new_n757), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G150), .B2(new_n770), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1177), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n786), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1174), .B1(new_n1173), .B2(new_n1172), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1163), .B1(new_n1189), .B2(new_n744), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1149), .B2(new_n746), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1162), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n849), .A2(new_n1075), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1116), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1160), .A2(KEYINPUT57), .A3(new_n1161), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n672), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1116), .A2(new_n1195), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1157), .A2(new_n1158), .A3(new_n1149), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(new_n1159), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1193), .B1(new_n1198), .B2(new_n1202), .ZN(G375));
  INV_X1    g1003(.A(new_n1088), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1194), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n957), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1089), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n765), .A2(G137), .B1(G128), .B2(new_n787), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n813), .B2(new_n759), .C1(new_n757), .C2(new_n1121), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G159), .B2(new_n776), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n213), .A2(new_n752), .B1(new_n762), .B2(new_n809), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n463), .B(new_n1211), .C1(G50), .C2(new_n770), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n556), .A2(new_n757), .B1(new_n766), .B2(new_n821), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1213), .A2(new_n1038), .A3(new_n985), .A4(new_n292), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G294), .A2(new_n791), .B1(new_n763), .B2(G107), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n547), .B2(new_n778), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G97), .B2(new_n776), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1210), .A2(new_n1212), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n730), .B1(new_n805), .B2(G68), .C1(new_n1218), .C2(new_n803), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n897), .B2(new_n745), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1088), .B2(new_n729), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1207), .A2(new_n1221), .ZN(G381));
  NAND3_X1  g1022(.A1(new_n977), .A2(new_n1004), .A3(new_n1072), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1200), .A2(new_n1159), .A3(new_n1226), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n673), .B1(new_n1228), .B2(new_n1199), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1192), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1117), .A2(new_n1141), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1224), .A2(new_n1230), .A3(new_n1232), .A4(new_n1233), .ZN(G407));
  OR3_X1    g1034(.A1(G375), .A2(G343), .A3(new_n1231), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1200), .A2(new_n1159), .A3(new_n728), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1191), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1199), .A2(new_n1206), .A3(new_n1201), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1162), .A2(KEYINPUT123), .A3(new_n1191), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1232), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT119), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1231), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1117), .A2(KEYINPUT119), .A3(new_n1141), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1244), .B1(new_n1248), .B2(G375), .ZN(new_n1249));
  INV_X1    g1049(.A(G213), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(G343), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1194), .B2(new_n1204), .ZN(new_n1255));
  AOI211_X1 g1055(.A(KEYINPUT60), .B(new_n1088), .C1(new_n849), .C2(new_n1075), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n672), .B(new_n1089), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(KEYINPUT124), .B(new_n829), .C1(new_n834), .C2(new_n835), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1258), .A2(new_n1221), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT124), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G384), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1257), .A2(new_n1259), .A3(new_n1262), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1251), .A2(G2897), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G393), .B(new_n800), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1072), .B1(new_n977), .B2(new_n1004), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1271), .B1(new_n1224), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(G390), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1271), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1223), .A3(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1265), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1262), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1249), .A2(new_n1281), .A3(new_n1252), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1282), .A2(KEYINPUT125), .A3(KEYINPUT63), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT63), .B1(new_n1282), .B2(KEYINPUT125), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1270), .B(new_n1277), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(G378), .A2(new_n1230), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1251), .B1(new_n1286), .B2(new_n1244), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT62), .B1(new_n1287), .B2(new_n1281), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(G378), .A2(new_n1230), .B1(new_n1232), .B2(new_n1243), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1280), .A4(new_n1251), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1270), .B(KEYINPUT126), .C1(new_n1288), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1282), .A2(new_n1290), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1287), .A2(KEYINPUT62), .A3(new_n1281), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT126), .B1(new_n1297), .B2(new_n1270), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1285), .B1(new_n1294), .B2(new_n1298), .ZN(G405));
  OAI21_X1  g1099(.A(new_n1286), .B1(new_n1231), .B2(new_n1230), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(new_n1280), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  OR3_X1    g1102(.A1(new_n1301), .A2(new_n1277), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1277), .A2(new_n1302), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1293), .A2(KEYINPUT127), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n1301), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1306), .ZN(G402));
endmodule


