//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G20), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT64), .Z(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n212), .B1(new_n216), .B2(new_n217), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  NAND2_X1  g0035(.A1(new_n202), .A2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(G68), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G107), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G97), .ZN(new_n243));
  INV_X1    g0043(.A(G97), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G107), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n241), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT76), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n213), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT16), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT7), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n254), .B1(new_n259), .B2(G20), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n237), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G58), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n237), .ZN(new_n267));
  OAI21_X1  g0067(.A(G20), .B1(new_n267), .B2(new_n201), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G159), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n253), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT75), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n268), .A2(KEYINPUT16), .A3(new_n270), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n265), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT7), .B1(new_n263), .B2(new_n207), .ZN(new_n276));
  NOR4_X1   g0076(.A1(new_n261), .A2(new_n262), .A3(new_n254), .A4(G20), .ZN(new_n277));
  OAI21_X1  g0077(.A(G68), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n268), .A2(KEYINPUT16), .A3(new_n270), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT75), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n252), .B(new_n272), .C1(new_n275), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  OR3_X1    g0083(.A1(new_n266), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n252), .B1(new_n206), .B2(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G20), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n290), .B2(new_n285), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT18), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  INV_X1    g0096(.A(G226), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G1698), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n298), .B1(G223), .B2(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G87), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  AOI21_X1  g0103(.A(G1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n296), .A3(G274), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n228), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(G169), .B2(new_n309), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n293), .A2(new_n294), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n273), .B1(new_n265), .B2(new_n274), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n278), .A2(KEYINPUT75), .A3(new_n279), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n252), .ZN(new_n318));
  INV_X1    g0118(.A(new_n271), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n278), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n320), .B2(new_n253), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n291), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT18), .B1(new_n322), .B2(new_n312), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n250), .B1(new_n314), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n309), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n301), .A2(new_n308), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n281), .A2(new_n329), .A3(new_n292), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(KEYINPUT76), .A2(KEYINPUT18), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n322), .B2(new_n312), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n322), .A2(KEYINPUT17), .A3(new_n329), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G1698), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n257), .B2(new_n258), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G223), .ZN(new_n340));
  AOI21_X1  g0140(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G222), .ZN(new_n342));
  INV_X1    g0142(.A(G77), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n340), .B(new_n342), .C1(new_n343), .C2(new_n259), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT66), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n296), .B1(new_n344), .B2(KEYINPUT66), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n305), .B1(new_n297), .B2(new_n307), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(G179), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n256), .A2(G20), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n283), .A2(new_n352), .A3(new_n284), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n269), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n318), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n286), .A2(G50), .ZN(new_n356));
  INV_X1    g0156(.A(new_n290), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n202), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n348), .B1(new_n345), .B2(new_n346), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(G169), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n351), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n360), .A2(KEYINPUT9), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n360), .A2(KEYINPUT9), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n365), .B(new_n366), .C1(new_n362), .C2(new_n325), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(G190), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT10), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n350), .A2(G200), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n368), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n364), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n337), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT77), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT71), .ZN(new_n379));
  INV_X1    g0179(.A(G238), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n305), .B1(new_n380), .B2(new_n307), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n297), .A2(new_n338), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n228), .A2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n382), .B(new_n383), .C1(new_n261), .C2(new_n262), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G97), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n296), .B1(new_n386), .B2(KEYINPUT70), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT70), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n384), .A2(new_n388), .A3(new_n385), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n381), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n379), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n327), .B1(new_n390), .B2(new_n391), .ZN(new_n393));
  INV_X1    g0193(.A(new_n389), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n388), .B1(new_n384), .B2(new_n385), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n394), .A2(new_n395), .A3(new_n296), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT71), .B(KEYINPUT13), .C1(new_n396), .C2(new_n381), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT72), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n392), .A2(new_n393), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n269), .A2(G50), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT73), .ZN(new_n404));
  INV_X1    g0204(.A(new_n352), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n405), .A2(new_n343), .B1(new_n207), .B2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n252), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT11), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n289), .A2(G20), .A3(new_n237), .A4(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(KEYINPUT74), .A2(KEYINPUT12), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n412), .B(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(G68), .B2(new_n286), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT13), .B1(new_n396), .B2(new_n381), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n390), .A2(new_n391), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(G200), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n402), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n310), .B1(new_n390), .B2(new_n391), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n392), .A2(new_n422), .A3(new_n397), .ZN(new_n423));
  INV_X1    g0223(.A(G169), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n417), .B2(new_n418), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI211_X1 g0227(.A(KEYINPUT14), .B(new_n424), .C1(new_n417), .C2(new_n418), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n416), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n339), .A2(G238), .B1(new_n263), .B2(G107), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n341), .A2(G232), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n296), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G244), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n305), .B1(new_n434), .B2(new_n307), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n310), .ZN(new_n437));
  INV_X1    g0237(.A(new_n282), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n269), .B1(G20), .B2(G77), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT68), .B1(new_n440), .B2(new_n405), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n440), .A2(new_n405), .A3(KEYINPUT68), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n252), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n290), .A2(G77), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(G77), .B2(new_n286), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n424), .B1(new_n433), .B2(new_n435), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n437), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n444), .B(new_n446), .C1(new_n436), .C2(new_n325), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n451), .A2(KEYINPUT69), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n451), .A2(KEYINPUT69), .B1(G190), .B2(new_n436), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n377), .A2(new_n378), .A3(new_n430), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n430), .A2(new_n454), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT77), .B1(new_n456), .B2(new_n376), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n357), .A2(new_n244), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(new_n206), .A3(G33), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT78), .B1(new_n256), .B2(G1), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n290), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n463), .A2(new_n252), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n459), .B1(new_n464), .B2(new_n244), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT6), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n244), .A2(new_n242), .ZN(new_n467));
  NOR2_X1   g0267(.A1(G97), .A2(G107), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n466), .B2(new_n243), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G20), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n276), .B2(new_n277), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n269), .A2(G77), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n465), .B1(new_n252), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n296), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n341), .A2(KEYINPUT4), .A3(G244), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT4), .B1(new_n341), .B2(G244), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(KEYINPUT79), .ZN(new_n480));
  OAI211_X1 g0280(.A(G244), .B(new_n338), .C1(new_n261), .C2(new_n262), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT79), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n339), .B2(G250), .ZN(new_n485));
  OAI211_X1 g0285(.A(G250), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(KEYINPUT80), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n476), .B1(new_n480), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n206), .A2(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G274), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n214), .B2(new_n295), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n303), .A2(G1), .ZN(new_n498));
  INV_X1    g0298(.A(new_n493), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n491), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(G257), .A3(new_n296), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT81), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n497), .B2(new_n501), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n489), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n475), .B1(new_n424), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n486), .A2(KEYINPUT80), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n259), .A2(new_n484), .A3(G250), .A4(G1698), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n479), .A2(KEYINPUT79), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT79), .B1(new_n481), .B2(new_n482), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n296), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n497), .A2(new_n501), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n508), .B1(new_n520), .B2(new_n310), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n489), .A2(new_n310), .A3(new_n505), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n507), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT83), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n520), .A2(new_n508), .A3(new_n310), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(new_n507), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n506), .A2(G200), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n531), .B(new_n475), .C1(new_n327), .C2(new_n506), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT19), .B1(new_n352), .B2(G97), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n263), .A2(G20), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G68), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT85), .B(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n468), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n207), .B1(new_n385), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT84), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT84), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n207), .C1(new_n385), .C2(new_n538), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n537), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n318), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n357), .A2(new_n440), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G87), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n464), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n296), .A2(G274), .A3(new_n498), .ZN(new_n549));
  AND2_X1   g0349(.A1(G33), .A2(G41), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n490), .B(G250), .C1(new_n550), .C2(new_n213), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G238), .B(new_n338), .C1(new_n261), .C2(new_n262), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(new_n556), .B2(new_n476), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(G190), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n557), .A2(new_n325), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n464), .A2(new_n440), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n562), .A2(new_n544), .A3(new_n545), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n557), .A2(G169), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n310), .B2(new_n557), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n559), .A2(new_n561), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  AND4_X1   g0367(.A1(new_n525), .A2(new_n530), .A3(new_n532), .A4(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G257), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n569));
  OAI211_X1 g0369(.A(G250), .B(new_n338), .C1(new_n261), .C2(new_n262), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G294), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g0372(.A(KEYINPUT5), .B(G41), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n498), .B1(new_n214), .B2(new_n295), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n572), .A2(new_n476), .B1(new_n574), .B2(G264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n497), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(G179), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n424), .B2(new_n576), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n242), .A2(KEYINPUT23), .A3(G20), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT23), .B1(new_n242), .B2(G20), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(G20), .B2(new_n555), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n259), .A2(new_n207), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n547), .B1(KEYINPUT87), .B2(KEYINPUT22), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT88), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT87), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT88), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n259), .A2(new_n590), .A3(new_n207), .A4(new_n585), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n587), .A2(new_n591), .B1(new_n588), .B2(new_n589), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n583), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT24), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n587), .A2(new_n591), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n588), .A2(new_n589), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n592), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(new_n583), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n318), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n464), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT25), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n290), .B2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(G107), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n578), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n601), .B1(new_n600), .B2(new_n583), .ZN(new_n611));
  AOI211_X1 g0411(.A(KEYINPUT24), .B(new_n582), .C1(new_n599), .C2(new_n592), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n252), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n576), .A2(new_n325), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(G190), .B2(new_n576), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n608), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  INV_X1    g0418(.A(G116), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n357), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n464), .B2(new_n619), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n477), .B(new_n207), .C1(G33), .C2(new_n244), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT86), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(G20), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n252), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n252), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(KEYINPUT20), .B(new_n622), .C1(new_n625), .C2(new_n626), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n621), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n574), .A2(G270), .B1(new_n496), .B2(new_n494), .ZN(new_n632));
  OAI211_X1 g0432(.A(G264), .B(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n633));
  OAI211_X1 g0433(.A(G257), .B(new_n338), .C1(new_n261), .C2(new_n262), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n257), .A2(G303), .A3(new_n258), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n476), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G169), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n618), .B1(new_n631), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n629), .A2(new_n630), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n641), .B(new_n620), .C1(new_n619), .C2(new_n464), .ZN(new_n642));
  INV_X1    g0442(.A(new_n639), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(KEYINPUT21), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(G200), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n632), .A2(new_n637), .A3(G190), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n631), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n632), .A2(new_n637), .A3(G179), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  AND4_X1   g0450(.A1(new_n640), .A2(new_n644), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n458), .A2(new_n568), .A3(new_n617), .A4(new_n651), .ZN(G372));
  NAND2_X1  g0452(.A1(new_n314), .A2(new_n323), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n419), .A2(G200), .ZN(new_n654));
  INV_X1    g0454(.A(new_n416), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n399), .B2(new_n401), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n429), .B1(new_n657), .B2(new_n449), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n332), .A2(new_n335), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n653), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n370), .A2(new_n374), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n661), .A2(new_n663), .B1(new_n351), .B2(new_n363), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n458), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n557), .A2(new_n310), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n556), .A2(new_n476), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n549), .A2(KEYINPUT89), .A3(new_n551), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT89), .B1(new_n549), .B2(new_n551), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n667), .B1(new_n673), .B2(G169), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n563), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(G200), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT90), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n559), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n578), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n613), .B2(new_n608), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n640), .A2(new_n644), .A3(new_n650), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n616), .B(new_n678), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n525), .A2(new_n530), .A3(new_n532), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n563), .B2(new_n674), .ZN(new_n684));
  INV_X1    g0484(.A(new_n524), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(new_n678), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n559), .A2(new_n561), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n564), .A2(new_n566), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n525), .B2(new_n530), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n691), .B2(new_n686), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n665), .B1(new_n666), .B2(new_n693), .ZN(G369));
  NAND2_X1  g0494(.A1(new_n289), .A2(new_n207), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  XOR2_X1   g0496(.A(new_n696), .B(KEYINPUT91), .Z(new_n697));
  INV_X1    g0497(.A(G213), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n695), .B2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G343), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n603), .B2(new_n609), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n617), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT92), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n617), .A2(new_n704), .A3(KEYINPUT92), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n680), .A2(new_n703), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n651), .B1(new_n631), .B2(new_n702), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n681), .A2(new_n642), .A3(new_n703), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n681), .A2(new_n702), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n707), .A2(new_n708), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n680), .A2(new_n702), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n717), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n210), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n537), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n217), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n702), .B1(new_n684), .B2(new_n692), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n678), .A2(KEYINPUT26), .A3(new_n528), .A4(new_n507), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT95), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT95), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n685), .A2(new_n735), .A3(KEYINPUT26), .A4(new_n678), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n525), .A2(new_n530), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT26), .B1(new_n738), .B2(new_n567), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(KEYINPUT29), .B(new_n702), .C1(new_n740), .C2(new_n684), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n732), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n575), .A2(new_n557), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n489), .A2(new_n744), .A3(new_n505), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT93), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n648), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n632), .A2(new_n637), .A3(KEYINPUT93), .A4(G179), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  AND4_X1   g0550(.A1(new_n310), .A2(new_n576), .A3(new_n672), .A4(new_n638), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(KEYINPUT30), .B1(new_n506), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n745), .B2(new_n749), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n743), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT94), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g0558(.A(KEYINPUT94), .B(new_n753), .C1(new_n745), .C2(new_n749), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n702), .B1(new_n760), .B2(new_n752), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n525), .A2(new_n530), .A3(new_n532), .A4(new_n567), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n610), .A2(new_n651), .A3(new_n616), .A4(new_n702), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n756), .B1(new_n761), .B2(KEYINPUT31), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G330), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n742), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n729), .B1(new_n766), .B2(G1), .ZN(G364));
  NOR2_X1   g0567(.A1(new_n288), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n206), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n724), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n213), .B1(G20), .B2(new_n424), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n207), .A2(G179), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT98), .B(G159), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n775), .A2(new_n327), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n263), .B(new_n782), .C1(G107), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n207), .A2(new_n310), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT96), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n207), .A2(new_n310), .A3(KEYINPUT96), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n776), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(KEYINPUT97), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G77), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n786), .A2(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n327), .A2(G200), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n207), .B1(new_n799), .B2(new_n310), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n798), .A2(new_n237), .B1(new_n244), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n202), .B1(new_n803), .B2(new_n536), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n799), .B1(new_n788), .B2(new_n789), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G58), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n785), .A2(new_n795), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n259), .B1(new_n778), .B2(G329), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n783), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G322), .B2(new_n807), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n803), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G294), .ZN(new_n816));
  INV_X1    g0616(.A(G326), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n800), .B1(new_n802), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT33), .B(G317), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n815), .B(new_n818), .C1(new_n797), .C2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n813), .B(new_n820), .C1(new_n821), .C2(new_n793), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n774), .B1(new_n809), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G13), .A2(G33), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G20), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n773), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n723), .A2(new_n263), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(G355), .B1(new_n619), .B2(new_n723), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n723), .A2(new_n259), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(G45), .B2(new_n217), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n241), .A2(new_n303), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n772), .B(new_n823), .C1(new_n827), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT99), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n713), .A2(new_n714), .A3(new_n826), .ZN(new_n836));
  INV_X1    g0636(.A(new_n716), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n771), .ZN(new_n838));
  INV_X1    g0638(.A(G330), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n713), .A2(new_n839), .A3(new_n714), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n835), .A2(new_n836), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NOR2_X1   g0642(.A1(new_n703), .A2(new_n449), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n452), .A2(new_n453), .B1(new_n703), .B2(new_n447), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n845), .B2(new_n450), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n730), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n702), .B(new_n848), .C1(new_n684), .C2(new_n692), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n771), .B1(new_n850), .B2(new_n765), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n765), .B2(new_n850), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n774), .A2(new_n825), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n771), .B1(G77), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(G150), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n798), .A2(new_n855), .B1(new_n802), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n807), .B2(G143), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n793), .B2(new_n779), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT102), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n860), .A2(KEYINPUT34), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(KEYINPUT34), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n259), .B1(new_n777), .B2(new_n863), .C1(new_n237), .C2(new_n783), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n800), .A2(new_n266), .B1(new_n803), .B2(new_n202), .ZN(new_n865));
  OR4_X1    g0665(.A1(new_n861), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n794), .A2(G116), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n797), .A2(KEYINPUT100), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n797), .A2(KEYINPUT100), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n263), .B1(new_n803), .B2(new_n242), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n870), .A2(G283), .B1(KEYINPUT101), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n871), .A2(KEYINPUT101), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n800), .A2(new_n244), .B1(new_n777), .B2(new_n821), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n802), .A2(new_n814), .B1(new_n783), .B2(new_n547), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n874), .B(new_n875), .C1(new_n807), .C2(G294), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n867), .A2(new_n872), .A3(new_n873), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n866), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n854), .B1(new_n878), .B2(new_n773), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n825), .B2(new_n848), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n852), .A2(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n768), .A2(new_n206), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n732), .A2(new_n741), .A3(new_n458), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT105), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT105), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n732), .A2(new_n741), .A3(new_n885), .A4(new_n458), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n664), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n653), .A2(new_n700), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n330), .B1(new_n322), .B2(new_n312), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n322), .A2(new_n700), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n293), .A2(new_n313), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n293), .A2(new_n701), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n330), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n889), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n891), .B1(new_n324), .B2(new_n336), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n892), .A2(new_n896), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n891), .B1(new_n653), .B2(new_n659), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n899), .A2(new_n902), .A3(KEYINPUT39), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT104), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n897), .A2(new_n904), .A3(new_n898), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n897), .B2(new_n898), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n898), .A2(new_n900), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n905), .A2(new_n906), .B1(KEYINPUT38), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n903), .B1(new_n908), .B2(KEYINPUT39), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n429), .A2(new_n703), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n888), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n849), .A2(new_n844), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n703), .A2(new_n416), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n421), .A2(new_n429), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n421), .B2(new_n429), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n913), .A2(new_n908), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n887), .B(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n898), .B2(new_n900), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n897), .A2(new_n898), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT104), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n897), .A2(new_n904), .A3(new_n898), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n425), .A2(new_n426), .ZN(new_n928));
  INV_X1    g0728(.A(new_n428), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n423), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n416), .B(new_n703), .C1(new_n657), .C2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n421), .A2(new_n429), .A3(new_n914), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n846), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI211_X1 g0733(.A(KEYINPUT106), .B(new_n743), .C1(new_n760), .C2(new_n752), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT106), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n520), .A2(new_n744), .A3(new_n747), .A4(new_n748), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT94), .B1(new_n936), .B2(new_n753), .ZN(new_n937));
  INV_X1    g0737(.A(new_n759), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n752), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n743), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n762), .A2(new_n763), .B1(new_n761), .B2(KEYINPUT31), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n933), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n922), .B1(new_n927), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT40), .B1(new_n899), .B2(new_n902), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  AND4_X1   g0747(.A1(new_n610), .A2(new_n651), .A3(new_n616), .A4(new_n702), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT31), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n939), .A2(new_n703), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n568), .A2(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n939), .A2(new_n940), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n939), .A2(new_n935), .A3(new_n940), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n458), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n947), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n947), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(G330), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n882), .B1(new_n921), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n921), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(new_n216), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(G116), .C1(new_n470), .C2(KEYINPUT35), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT103), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(KEYINPUT103), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT36), .ZN(new_n969));
  OAI21_X1  g0769(.A(G77), .B1(new_n266), .B2(new_n237), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n236), .B1(new_n970), .B2(new_n217), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(G1), .A3(new_n288), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n962), .A2(new_n969), .A3(new_n972), .ZN(G367));
  INV_X1    g0773(.A(new_n766), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n702), .A2(new_n475), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n683), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n685), .A2(new_n703), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n719), .B2(new_n720), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT109), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  INV_X1    g0784(.A(new_n978), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n721), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n719), .A2(KEYINPUT45), .A3(new_n720), .A4(new_n978), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n717), .A2(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n717), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n986), .A2(new_n987), .ZN(new_n992));
  OAI211_X1 g0792(.A(KEYINPUT109), .B(new_n989), .C1(new_n981), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n719), .B1(new_n711), .B2(new_n718), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n837), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n974), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n724), .B(KEYINPUT41), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n769), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n976), .A2(KEYINPUT107), .A3(new_n977), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT107), .B1(new_n976), .B2(new_n977), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n717), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT108), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n985), .A2(new_n719), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT42), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n680), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n738), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n703), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1005), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n703), .A2(new_n548), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n678), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n703), .A2(new_n675), .A3(new_n548), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1005), .B(new_n1016), .C1(new_n1008), .C2(new_n1011), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT43), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1004), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1003), .B(new_n1021), .C1(new_n1026), .C2(new_n1023), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n999), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1017), .A2(new_n826), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n794), .A2(G283), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n803), .A2(new_n619), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n806), .A2(new_n814), .B1(new_n1031), .B2(KEYINPUT46), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(KEYINPUT46), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n870), .A2(G294), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n242), .A2(new_n800), .B1(new_n802), .B2(new_n821), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n783), .A2(new_n244), .ZN(new_n1036));
  INV_X1    g0836(.A(G317), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n263), .B1(new_n777), .B2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1030), .A2(new_n1033), .A3(new_n1034), .A4(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n783), .A2(new_n343), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n263), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT111), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n870), .B2(new_n780), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n802), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1046), .A2(G143), .B1(new_n778), .B2(G137), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n266), .B2(new_n803), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1045), .B(new_n1049), .C1(new_n202), .C2(new_n793), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n800), .A2(new_n237), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n807), .B2(G150), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT110), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1040), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT47), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n773), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n830), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n827), .B1(new_n210), .B2(new_n440), .C1(new_n1057), .C2(new_n234), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1029), .A2(new_n1056), .A3(new_n771), .A4(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1028), .A2(new_n1059), .ZN(G387));
  NAND2_X1  g0860(.A1(new_n231), .A2(G45), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT112), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n282), .A2(G50), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1064));
  XNOR2_X1  g0864(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n726), .B(new_n303), .C1(new_n237), .C2(new_n343), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1062), .B(new_n830), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n828), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(G107), .B2(new_n210), .C1(new_n726), .C2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n772), .B1(new_n1069), .B2(new_n827), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n807), .A2(G317), .B1(G322), .B2(new_n1046), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n870), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(new_n814), .B2(new_n793), .C1(new_n1072), .C2(new_n821), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT115), .Z(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n800), .A2(new_n811), .B1(new_n803), .B2(new_n816), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1079), .A2(KEYINPUT49), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n263), .B1(new_n777), .B2(new_n817), .C1(new_n619), .C2(new_n783), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT116), .Z(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1079), .B2(KEYINPUT49), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n793), .A2(new_n237), .B1(new_n285), .B2(new_n798), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT114), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n803), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(G77), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n263), .B(new_n1036), .C1(G150), .C2(new_n778), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n800), .A2(new_n440), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G159), .B2(new_n1046), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n807), .A2(G50), .ZN(new_n1091));
  AND4_X1   g0891(.A1(new_n1087), .A2(new_n1088), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1080), .A2(new_n1083), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1070), .B1(new_n1093), .B2(new_n774), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n712), .B2(new_n826), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n770), .B2(new_n996), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n996), .A2(new_n766), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(KEYINPUT117), .A3(new_n724), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n766), .B2(new_n996), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT117), .B1(new_n1097), .B2(new_n724), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(G393));
  NAND3_X1  g0901(.A1(new_n994), .A2(new_n766), .A3(new_n996), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n991), .A2(new_n993), .A3(new_n1097), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n724), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n994), .A2(new_n770), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1002), .A2(G20), .A3(new_n825), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n263), .B1(new_n778), .B2(G143), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n237), .B2(new_n803), .C1(new_n547), .C2(new_n783), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT118), .Z(new_n1109));
  INV_X1    g0909(.A(G159), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n806), .A2(new_n1110), .B1(new_n855), .B2(new_n802), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT51), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n794), .A2(new_n438), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n800), .A2(new_n343), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n870), .B2(G50), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1109), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT119), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n259), .B1(new_n778), .B2(G322), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n242), .B2(new_n783), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n800), .A2(new_n619), .B1(new_n803), .B2(new_n811), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n870), .C2(G303), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n816), .B2(new_n793), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n806), .A2(new_n821), .B1(new_n1037), .B2(new_n802), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT52), .Z(new_n1125));
  OAI21_X1  g0925(.A(new_n1118), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n773), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n827), .B1(new_n244), .B2(new_n210), .C1(new_n1057), .C2(new_n248), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n771), .A3(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1104), .B(new_n1105), .C1(new_n1106), .C2(new_n1130), .ZN(G390));
  AOI21_X1  g0931(.A(new_n839), .B1(new_n951), .B2(new_n955), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n933), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n899), .A2(new_n902), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT39), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n927), .B2(new_n1136), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n913), .A2(new_n918), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n911), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1135), .A2(new_n910), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n845), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n449), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n702), .B(new_n1144), .C1(new_n740), .C2(new_n684), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n844), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1142), .B1(new_n1146), .B2(new_n918), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1134), .B1(new_n1140), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n917), .B1(new_n849), .B2(new_n844), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n909), .B1(new_n1149), .B2(new_n910), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n764), .A2(new_n918), .A3(G330), .A4(new_n848), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n917), .B1(new_n1145), .B2(new_n844), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(new_n1151), .C1(new_n1152), .C2(new_n1142), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n769), .ZN(new_n1155));
  INV_X1    g0955(.A(G125), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n259), .B1(new_n777), .B2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n800), .A2(new_n1110), .B1(new_n783), .B2(new_n202), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(G128), .C2(new_n1046), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n863), .B2(new_n806), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n803), .A2(new_n855), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1072), .B2(new_n856), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1160), .B(new_n1163), .C1(new_n794), .C2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n803), .A2(new_n547), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1167), .B(new_n1114), .C1(G283), .C2(new_n1046), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n263), .B1(new_n777), .B2(new_n816), .C1(new_n237), .C2(new_n783), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G116), .B2(new_n807), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n1072), .C2(new_n242), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n794), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n773), .B1(new_n1166), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n285), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n771), .C1(new_n1174), .C2(new_n853), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n909), .B2(new_n824), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1155), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n458), .A2(new_n1132), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n764), .A2(G330), .A3(new_n848), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n917), .A2(new_n1179), .B1(new_n1132), .B2(new_n933), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n913), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1145), .A2(new_n1151), .A3(new_n844), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n918), .B1(new_n1132), .B2(new_n848), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1180), .A2(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n887), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1154), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1178), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n664), .B(new_n1187), .C1(new_n884), .C2(new_n886), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1188), .A2(new_n1153), .A3(new_n1148), .A4(new_n1184), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1186), .A2(new_n1189), .A3(new_n724), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1177), .A2(new_n1190), .ZN(G378));
  INV_X1    g0991(.A(KEYINPUT123), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT122), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n848), .B1(new_n915), .B2(new_n916), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n951), .B2(new_n955), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT40), .B1(new_n1195), .B2(new_n908), .ZN(new_n1196));
  OAI21_X1  g0996(.A(G330), .B1(new_n944), .B2(new_n946), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n902), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n922), .B1(new_n1199), .B2(new_n924), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n839), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n945), .A3(KEYINPUT122), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n701), .A2(new_n361), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n375), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n375), .A2(new_n1203), .ZN(new_n1206));
  OAI21_X1  g1006(.A(KEYINPUT120), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1208));
  OR2_X1    g1008(.A1(new_n375), .A2(new_n1203), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT120), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1204), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1207), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1208), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1198), .A2(new_n1202), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n1193), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1215), .A2(new_n920), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n920), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1192), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n920), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1215), .A2(new_n920), .A3(new_n1217), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(KEYINPUT123), .A3(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1184), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1188), .B1(new_n1154), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1220), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n1189), .B2(new_n1188), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n725), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1220), .A2(new_n1225), .A3(new_n770), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n771), .B1(G50), .B2(new_n853), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n778), .C2(G124), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n779), .B2(new_n783), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n803), .A2(new_n1164), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n798), .A2(new_n863), .B1(new_n855), .B2(new_n800), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(G125), .C2(new_n1046), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n807), .A2(G128), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n793), .C2(new_n856), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1238), .B1(new_n1243), .B2(KEYINPUT59), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(KEYINPUT59), .B2(new_n1243), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n783), .A2(new_n266), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1087), .B1(new_n798), .B2(new_n244), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(G116), .C2(new_n1046), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n302), .B(new_n263), .C1(new_n777), .C2(new_n811), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1249), .B(new_n1051), .C1(new_n807), .C2(G107), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(new_n440), .C2(new_n793), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT58), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n263), .A2(new_n302), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G50), .B1(new_n256), .B2(new_n302), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1251), .A2(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1245), .B(new_n1255), .C1(new_n1252), .C2(new_n1251), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1236), .B1(new_n1256), .B2(new_n773), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1216), .B2(new_n825), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT121), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1235), .A2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1234), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(G375));
  NAND2_X1  g1062(.A1(new_n917), .A2(new_n824), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n771), .B1(G68), .B2(new_n853), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n870), .A2(G116), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n803), .A2(new_n244), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1266), .B(new_n1089), .C1(G294), .C2(new_n1046), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n807), .A2(G283), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n259), .B(new_n1041), .C1(G303), .C2(new_n778), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n793), .A2(new_n242), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n870), .A2(new_n1165), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n202), .A2(new_n800), .B1(new_n802), .B2(new_n863), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G159), .B2(new_n1086), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n807), .A2(G137), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n263), .B(new_n1246), .C1(G128), .C2(new_n778), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n793), .A2(new_n855), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1270), .A2(new_n1271), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1264), .B1(new_n1279), .B2(new_n773), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1184), .A2(new_n770), .B1(new_n1263), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1185), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(new_n998), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1184), .B1(new_n887), .B2(new_n1178), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1281), .B1(new_n1283), .B2(new_n1284), .ZN(G381));
  OR2_X1    g1085(.A1(G390), .A2(G384), .ZN(new_n1286));
  OR2_X1    g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1286), .A2(G378), .A3(new_n1287), .A4(G381), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1288), .A2(new_n1059), .A3(new_n1028), .A4(new_n1261), .ZN(G407));
  INV_X1    g1089(.A(G378), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n698), .A2(G343), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1261), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1234), .A2(G378), .A3(new_n1260), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1232), .A2(new_n770), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1259), .B(new_n1297), .C1(new_n1228), .C2(new_n998), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1290), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1291), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n887), .A2(new_n1178), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(KEYINPUT60), .A3(new_n1226), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n724), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1284), .B1(KEYINPUT60), .B2(new_n1185), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G384), .B(new_n1281), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1185), .A2(KEYINPUT60), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1301), .A2(new_n1226), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n724), .A3(new_n1302), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G384), .B1(new_n1310), .B2(new_n1281), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G2897), .B(new_n1291), .C1(new_n1306), .C2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1281), .ZN(new_n1313));
  INV_X1    g1113(.A(G384), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1291), .A2(G2897), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(new_n1305), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1312), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1295), .B1(new_n1300), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(KEYINPUT126), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1321), .B(new_n1295), .C1(new_n1300), .C2(new_n1318), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1300), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT62), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1320), .A2(new_n1322), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT124), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1300), .A2(KEYINPUT124), .A3(new_n1323), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT62), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1294), .B1(new_n1326), .B2(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(G387), .B(G390), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1028), .A2(G390), .A3(new_n1059), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(KEYINPUT125), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(G393), .B(G396), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1332), .B(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT62), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1329), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT124), .B1(new_n1300), .B2(new_n1323), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1338), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  AOI22_X1  g1141(.A1(new_n1319), .A2(KEYINPUT126), .B1(new_n1324), .B2(KEYINPUT62), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(KEYINPUT127), .A4(new_n1322), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1331), .A2(new_n1337), .A3(new_n1343), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1323), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1337), .A2(new_n1345), .A3(new_n1319), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1346), .B1(KEYINPUT63), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1344), .A2(new_n1348), .ZN(G405));
  NOR2_X1   g1149(.A1(new_n1261), .A2(G378), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1296), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  XOR2_X1   g1152(.A(new_n1352), .B(new_n1323), .Z(new_n1353));
  XNOR2_X1  g1153(.A(new_n1353), .B(new_n1337), .ZN(G402));
endmodule


