//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  OR3_X1    g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n207));
  OAI21_X1  g0007(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G250), .B1(G257), .B2(G264), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n203), .A2(G50), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n212), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n220), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n201), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  OR2_X1    g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G223), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G222), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n249), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n253), .B1(new_n254), .B2(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n213), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n261), .A2(new_n265), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G169), .ZN(new_n271));
  INV_X1    g0071(.A(G179), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(new_n270), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n214), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n214), .A2(new_n277), .A3(KEYINPUT69), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G20), .B2(G33), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n274), .B1(new_n275), .B2(new_n276), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n284), .A2(new_n285), .A3(new_n213), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n284), .B2(new_n213), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n283), .A2(new_n289), .B1(new_n241), .B2(new_n291), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n286), .A2(new_n287), .A3(new_n291), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n264), .A2(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G50), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n273), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n284), .A2(new_n213), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n281), .A2(new_n275), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT15), .B(G87), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n300), .A2(new_n276), .B1(new_n214), .B2(new_n254), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT70), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n290), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n264), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n298), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G77), .A3(new_n294), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n254), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n252), .A2(G238), .ZN(new_n311));
  INV_X1    g0111(.A(G107), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n312), .B2(new_n255), .C1(new_n233), .C2(new_n257), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n262), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n267), .B1(new_n268), .B2(G244), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n319), .A3(new_n315), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n310), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n316), .A2(new_n272), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n314), .B2(new_n315), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n310), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n270), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G190), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n270), .A2(G200), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n292), .A2(KEYINPUT9), .A3(new_n295), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT9), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n296), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n336));
  AOI211_X1 g0136(.A(new_n297), .B(new_n327), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n275), .B1(new_n264), .B2(G20), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n293), .A2(new_n338), .B1(new_n291), .B2(new_n275), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT73), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n255), .B2(G20), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n202), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(G58), .B(G68), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G20), .ZN(new_n351));
  INV_X1    g0151(.A(G159), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n281), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n341), .B(new_n342), .C1(new_n349), .C2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n354), .A2(new_n298), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n342), .B1(new_n349), .B2(new_n353), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n349), .A2(new_n353), .A3(new_n342), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(KEYINPUT73), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n340), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n261), .A2(G232), .A3(new_n265), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n266), .B2(new_n265), .ZN(new_n361));
  OAI211_X1 g0161(.A(G226), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT74), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT74), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n255), .A2(new_n364), .A3(G226), .A4(G1698), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G87), .ZN(new_n366));
  OAI211_X1 g0166(.A(G223), .B(new_n249), .C1(new_n345), .C2(new_n346), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n363), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n361), .B1(new_n368), .B2(new_n262), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n272), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G169), .B2(new_n369), .ZN(new_n371));
  OR3_X1    g0171(.A1(new_n359), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n347), .B2(new_n214), .ZN(new_n373));
  NOR4_X1   g0173(.A1(new_n345), .A2(new_n346), .A3(new_n343), .A4(G20), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n278), .A2(new_n280), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(G159), .B1(new_n350), .B2(G20), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT16), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(KEYINPUT16), .A3(new_n377), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n341), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n354), .A2(new_n298), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n339), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n371), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT18), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n372), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n366), .B(new_n367), .C1(new_n362), .C2(KEYINPUT74), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n364), .B1(new_n252), .B2(G226), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n262), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n361), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n319), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(G200), .B2(new_n369), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(new_n339), .C1(new_n380), .C2(new_n381), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT76), .B1(new_n393), .B2(KEYINPUT17), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n359), .A2(new_n395), .A3(new_n396), .A4(new_n392), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT75), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT75), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n393), .A2(new_n401), .A3(KEYINPUT17), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n386), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n252), .A2(KEYINPUT71), .A3(G232), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  INV_X1    g0206(.A(G226), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n257), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT71), .B1(new_n252), .B2(G232), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n262), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n267), .B1(new_n268), .B2(G238), .ZN(new_n411));
  XOR2_X1   g0211(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n412), .B1(new_n410), .B2(new_n411), .ZN(new_n415));
  OAI21_X1  g0215(.A(G200), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n276), .A2(new_n254), .B1(new_n214), .B2(G68), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(G50), .B2(new_n376), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n288), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n419), .A2(KEYINPUT11), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT12), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n308), .B2(new_n202), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n290), .A2(KEYINPUT12), .A3(G68), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n306), .A2(G68), .A3(new_n294), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(KEYINPUT11), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n420), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n410), .A2(new_n411), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  OAI211_X1 g0230(.A(G190), .B(new_n413), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n416), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(G169), .B1(new_n414), .B2(new_n415), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(G169), .C1(new_n414), .C2(new_n415), .ZN(new_n436));
  OAI211_X1 g0236(.A(G179), .B(new_n413), .C1(new_n429), .C2(new_n430), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n432), .B1(new_n438), .B2(new_n427), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n337), .A2(new_n404), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G13), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G1), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(G20), .A3(new_n312), .ZN(new_n443));
  XOR2_X1   g0243(.A(new_n443), .B(KEYINPUT25), .Z(new_n444));
  NAND2_X1  g0244(.A1(new_n298), .A2(KEYINPUT68), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n277), .B2(G1), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n264), .A2(KEYINPUT77), .A3(G33), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n284), .A2(new_n285), .A3(new_n213), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n445), .A2(new_n449), .A3(new_n290), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n444), .B1(new_n312), .B2(new_n451), .ZN(new_n452));
  OR3_X1    g0252(.A1(new_n214), .A2(KEYINPUT23), .A3(G107), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT23), .B1(new_n214), .B2(G107), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n453), .B(new_n454), .C1(G20), .C2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n214), .B(G87), .C1(new_n345), .C2(new_n346), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT86), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n255), .A2(new_n214), .A3(G87), .A4(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n458), .A2(KEYINPUT86), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n456), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT87), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT87), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n464), .B1(new_n461), .B2(new_n462), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(KEYINPUT24), .C1(new_n470), .C2(new_n456), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n452), .B1(new_n473), .B2(new_n298), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n255), .A2(G257), .A3(G1698), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G294), .ZN(new_n476));
  OAI21_X1  g0276(.A(G250), .B1(new_n345), .B2(new_n346), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n475), .B(new_n476), .C1(G1698), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G41), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(KEYINPUT79), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n264), .B(G45), .C1(new_n479), .C2(KEYINPUT5), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n262), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n478), .A2(new_n262), .B1(new_n487), .B2(G264), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(G41), .ZN(new_n491));
  OAI211_X1 g0291(.A(KEYINPUT80), .B(new_n479), .C1(new_n481), .C2(new_n483), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n485), .A2(new_n266), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n317), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G190), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n474), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n495), .A2(new_n272), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n324), .B1(new_n488), .B2(new_n494), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT88), .B1(new_n474), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT88), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n495), .A2(G169), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n272), .B2(new_n495), .ZN(new_n505));
  INV_X1    g0305(.A(new_n298), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n470), .A2(KEYINPUT24), .A3(new_n456), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT24), .B1(new_n470), .B2(new_n456), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(KEYINPUT87), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(new_n471), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n503), .B(new_n505), .C1(new_n510), .C2(new_n452), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G1698), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(G244), .C1(new_n346), .C2(new_n345), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  INV_X1    g0316(.A(G244), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n250), .B2(new_n251), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n515), .B(new_n516), .C1(new_n518), .C2(KEYINPUT4), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n249), .B1(new_n477), .B2(KEYINPUT4), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n262), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n482), .A2(KEYINPUT79), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n523));
  AOI21_X1  g0323(.A(G41), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n261), .B(G257), .C1(new_n524), .C2(new_n485), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n521), .A2(G190), .A3(new_n494), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n494), .A2(new_n525), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(KEYINPUT81), .A3(new_n521), .A4(G190), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  AND2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n312), .A2(KEYINPUT6), .A3(G97), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n537), .A2(new_n214), .B1(new_n254), .B2(new_n281), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n312), .B1(new_n344), .B2(new_n348), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n298), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G97), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n451), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n290), .A2(G97), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n540), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(G107), .B1(new_n373), .B2(new_n374), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n535), .A2(new_n536), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G20), .B1(G77), .B2(new_n376), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n544), .B1(new_n552), .B2(new_n298), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(KEYINPUT78), .A3(new_n543), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n529), .A2(new_n521), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n531), .A2(new_n548), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n529), .A2(new_n272), .A3(new_n521), .ZN(new_n558));
  AOI21_X1  g0358(.A(G169), .B1(new_n529), .B2(new_n521), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT82), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n494), .A2(new_n525), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n477), .A2(KEYINPUT4), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n513), .B1(new_n347), .B2(new_n517), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n564), .A2(new_n515), .A3(new_n565), .A4(new_n516), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n262), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT82), .A3(new_n272), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n561), .A2(new_n568), .A3(new_n546), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n557), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n214), .B1(new_n406), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G87), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n541), .A3(new_n312), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n214), .B(G68), .C1(new_n345), .C2(new_n346), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n571), .B1(new_n406), .B2(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n298), .B1(new_n308), .B2(new_n300), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT84), .ZN(new_n580));
  INV_X1    g0380(.A(new_n300), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n293), .A2(new_n580), .A3(new_n581), .A4(new_n449), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT84), .B1(new_n451), .B2(new_n300), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G238), .B(new_n249), .C1(new_n345), .C2(new_n346), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n455), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n262), .ZN(new_n588));
  INV_X1    g0388(.A(G45), .ZN(new_n589));
  OAI21_X1  g0389(.A(G250), .B1(new_n589), .B2(G1), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n264), .A2(G45), .A3(G274), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n259), .B2(new_n260), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n324), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n584), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n592), .B1(new_n587), .B2(new_n262), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n272), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(KEYINPUT83), .A3(new_n272), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n293), .A2(G87), .A3(new_n449), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n579), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n597), .A2(new_n317), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n319), .B(new_n592), .C1(new_n587), .C2(new_n262), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n596), .A2(new_n602), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n261), .B(G270), .C1(new_n524), .C2(new_n485), .ZN(new_n609));
  OAI211_X1 g0409(.A(G264), .B(G1698), .C1(new_n345), .C2(new_n346), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n250), .A2(G303), .A3(new_n251), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n249), .C1(new_n345), .C2(new_n346), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n255), .A2(KEYINPUT85), .A3(G257), .A4(new_n249), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n494), .B(new_n609), .C1(new_n617), .C2(new_n261), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n277), .A2(G97), .ZN(new_n619));
  AOI21_X1  g0419(.A(G20), .B1(new_n619), .B2(new_n516), .ZN(new_n620));
  INV_X1    g0420(.A(G116), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n214), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n298), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(KEYINPUT20), .B(new_n298), .C1(new_n620), .C2(new_n622), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n621), .B1(new_n447), .B2(new_n448), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n621), .A2(new_n308), .B1(new_n306), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n618), .A2(new_n630), .A3(G169), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n616), .ZN(new_n634));
  INV_X1    g0434(.A(new_n612), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n261), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n494), .A2(new_n609), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n636), .A2(new_n637), .A3(new_n272), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n631), .A2(new_n632), .B1(new_n630), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n262), .ZN(new_n641));
  INV_X1    g0441(.A(new_n637), .ZN(new_n642));
  AOI21_X1  g0442(.A(G200), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n636), .A2(new_n637), .A3(G190), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n627), .B(new_n629), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n608), .A2(new_n633), .A3(new_n639), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n570), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n440), .A2(new_n498), .A3(new_n512), .A4(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n438), .A2(new_n427), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n432), .B2(new_n326), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n393), .A2(new_n401), .A3(KEYINPUT17), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n401), .B1(new_n393), .B2(KEYINPUT17), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n394), .B(new_n397), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n372), .A2(new_n385), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n335), .A2(new_n336), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n297), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n596), .A2(new_n598), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n607), .A2(new_n604), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT78), .B1(new_n553), .B2(new_n543), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n506), .B1(new_n549), .B2(new_n551), .ZN(new_n663));
  NOR4_X1   g0463(.A1(new_n663), .A2(new_n547), .A3(new_n542), .A4(new_n544), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n561), .A2(new_n568), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT89), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n558), .A2(new_n560), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT82), .B1(new_n567), .B2(G169), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n558), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n548), .A2(new_n554), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AOI211_X1 g0473(.A(KEYINPUT26), .B(new_n661), .C1(new_n667), .C2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n659), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n670), .A2(new_n546), .A3(new_n608), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(new_n661), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n474), .A2(new_n501), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n633), .A2(new_n639), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n498), .A2(new_n569), .A3(new_n557), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n440), .B1(new_n674), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n658), .A2(new_n684), .ZN(G369));
  INV_X1    g0485(.A(new_n680), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n645), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n442), .A2(new_n214), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(G213), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n630), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n680), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G330), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n693), .B1(new_n510), .B2(new_n452), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n502), .A2(new_n511), .A3(new_n498), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n679), .A2(new_n693), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n693), .B(KEYINPUT90), .Z(new_n705));
  NAND2_X1  g0505(.A1(new_n679), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n693), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n680), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(G399));
  NOR4_X1   g0510(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G1), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n210), .A2(G41), .ZN(new_n713));
  MUX2_X1   g0513(.A(new_n712), .B(new_n217), .S(new_n713), .Z(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT91), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND4_X1  g0516(.A1(new_n512), .A2(new_n647), .A3(new_n498), .A4(new_n705), .ZN(new_n717));
  AND4_X1   g0517(.A1(new_n488), .A2(new_n521), .A3(new_n529), .A4(new_n597), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n638), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n597), .A2(G179), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n495), .A2(new_n555), .A3(new_n618), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT30), .B1(new_n718), .B2(new_n638), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n693), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n705), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n717), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(new_n682), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n686), .A2(new_n502), .A3(new_n511), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n732), .A2(new_n733), .A3(new_n660), .ZN(new_n734));
  INV_X1    g0534(.A(new_n608), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n569), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT26), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n675), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n661), .B1(new_n667), .B2(new_n673), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n707), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n705), .B1(new_n683), .B2(new_n674), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n742), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n731), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n716), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n699), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n697), .A2(new_n698), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n441), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n264), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OR3_X1    g0552(.A1(new_n713), .A2(KEYINPUT92), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT92), .B1(new_n713), .B2(new_n752), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n748), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n756), .B(KEYINPUT93), .Z(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n697), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n213), .B1(G20), .B2(new_n324), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n243), .A2(G45), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n217), .A2(new_n589), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n210), .B(new_n255), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n209), .A2(G355), .A3(new_n255), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G116), .B2(new_n209), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n765), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n319), .A2(KEYINPUT96), .A3(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(KEYINPUT96), .B1(new_n319), .B2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n774), .A2(G179), .A3(new_n317), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n312), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n214), .A2(new_n319), .A3(new_n317), .A4(G179), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n347), .B(new_n777), .C1(G87), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(G20), .A2(G179), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT95), .Z(new_n781));
  NOR2_X1   g0581(.A1(new_n319), .A2(new_n317), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n319), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G50), .A2(new_n784), .B1(new_n787), .B2(G58), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n774), .A2(G179), .A3(G200), .ZN(new_n789));
  AOI21_X1  g0589(.A(KEYINPUT32), .B1(new_n789), .B2(G159), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n789), .A2(KEYINPUT32), .A3(G159), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n779), .B(new_n788), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G179), .A2(G200), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n214), .B1(new_n793), .B2(G190), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT97), .Z(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G97), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n781), .A2(new_n319), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(new_n317), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n796), .B1(new_n799), .B2(new_n254), .C1(new_n202), .C2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G322), .A2(new_n787), .B1(new_n784), .B2(G326), .ZN(new_n803));
  INV_X1    g0603(.A(G329), .ZN(new_n804));
  INV_X1    g0604(.A(new_n789), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  INV_X1    g0607(.A(new_n778), .ZN(new_n808));
  INV_X1    g0608(.A(G303), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n347), .B1(new_n794), .B2(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G283), .B2(new_n775), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT33), .B(G317), .Z(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n812), .B2(new_n799), .C1(new_n801), .C2(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n792), .A2(new_n802), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n755), .B1(new_n815), .B2(new_n764), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n763), .A2(new_n771), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n757), .A2(new_n817), .ZN(G396));
  INV_X1    g0618(.A(new_n755), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n326), .A2(new_n693), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n310), .A2(new_n693), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n326), .B1(new_n321), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n744), .B(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n819), .B1(new_n825), .B2(new_n731), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n731), .B2(new_n825), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n764), .A2(new_n758), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n755), .B1(new_n254), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n801), .A2(new_n830), .B1(new_n783), .B2(new_n809), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G116), .B2(new_n798), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT98), .Z(new_n833));
  NOR2_X1   g0633(.A1(new_n776), .A2(new_n573), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n255), .B1(new_n778), .B2(G107), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n787), .A2(G294), .B1(new_n789), .B2(G311), .ZN(new_n837));
  AND4_X1   g0637(.A1(new_n796), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G137), .A2(new_n784), .B1(new_n787), .B2(G143), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n839), .B1(new_n799), .B2(new_n352), .C1(new_n282), .C2(new_n801), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT34), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n255), .B1(new_n794), .B2(new_n201), .C1(new_n808), .C2(new_n241), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n776), .A2(new_n202), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n842), .B(new_n843), .C1(G132), .C2(new_n789), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n833), .A2(new_n838), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n764), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n829), .B1(new_n824), .B2(new_n759), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n827), .A2(new_n847), .ZN(G384));
  OR2_X1    g0648(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(G116), .A3(new_n215), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(KEYINPUT35), .B2(new_n550), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT99), .B(KEYINPUT36), .Z(new_n853));
  OAI21_X1  g0653(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n217), .A2(new_n854), .B1(G50), .B2(new_n202), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n264), .A2(G13), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n852), .A2(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  INV_X1    g0658(.A(new_n691), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n382), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n653), .B2(new_n655), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT100), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n384), .A2(new_n860), .A3(new_n393), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n860), .B2(new_n862), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n868), .A2(new_n393), .A3(new_n384), .A4(new_n860), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n858), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n867), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n356), .A2(new_n379), .A3(new_n289), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n339), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n383), .B2(new_n859), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .A3(new_n393), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(new_n859), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT38), .B(new_n877), .C1(new_n404), .C2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n427), .A2(new_n693), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n439), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n427), .B(new_n693), .C1(new_n438), .C2(new_n432), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n823), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n717), .A2(new_n727), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT101), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT40), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n878), .B1(new_n653), .B2(new_n655), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n872), .A2(new_n876), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n858), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT40), .B1(new_n891), .B2(new_n879), .ZN(new_n892));
  AND2_X1   g0692(.A1(KEYINPUT101), .A2(KEYINPUT40), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n886), .B(new_n884), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n440), .A2(new_n886), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n895), .B(new_n896), .Z(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n698), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n882), .A2(new_n883), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n705), .B(new_n824), .C1(new_n683), .C2(new_n674), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(new_n820), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n891), .A2(new_n879), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n386), .B2(new_n691), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n649), .A2(new_n693), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n871), .A2(new_n879), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n891), .B2(new_n879), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n745), .B(new_n440), .C1(new_n741), .C2(new_n742), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n658), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n909), .B(new_n911), .Z(new_n912));
  NOR2_X1   g0712(.A1(new_n898), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT102), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n898), .A2(new_n912), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n914), .B(new_n915), .C1(new_n264), .C2(new_n750), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n913), .A2(KEYINPUT102), .ZN(new_n917));
  OAI221_X1 g0717(.A(new_n857), .B1(new_n852), .B2(new_n853), .C1(new_n916), .C2(new_n917), .ZN(G367));
  INV_X1    g0718(.A(new_n704), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n557), .B(new_n569), .C1(new_n665), .C2(new_n705), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n670), .A2(new_n672), .A3(new_n728), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n604), .A2(new_n707), .ZN(new_n924));
  MUX2_X1   g0724(.A(new_n661), .B(new_n659), .S(new_n924), .Z(new_n925));
  INV_X1    g0725(.A(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n923), .B(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n703), .A2(new_n680), .A3(new_n707), .A4(new_n922), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n931));
  INV_X1    g0731(.A(new_n922), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n569), .B1(new_n932), .B2(new_n512), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n705), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n930), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n926), .B2(new_n925), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n928), .B(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n713), .B(KEYINPUT41), .Z(new_n938));
  OAI21_X1  g0738(.A(new_n706), .B1(new_n701), .B2(new_n708), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n932), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT44), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n709), .A2(new_n706), .A3(new_n922), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT45), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n945), .A3(new_n704), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n943), .B(KEYINPUT45), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n919), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n701), .A2(new_n702), .A3(new_n708), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n709), .B1(KEYINPUT103), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(KEYINPUT103), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n950), .A2(new_n951), .A3(new_n699), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n699), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n946), .A2(new_n948), .A3(new_n746), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n938), .B1(new_n955), .B2(new_n746), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n751), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n956), .A2(KEYINPUT104), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n937), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n776), .A2(new_n541), .ZN(new_n961));
  INV_X1    g0761(.A(G317), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n805), .A2(new_n962), .B1(new_n809), .B2(new_n786), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n961), .B(new_n963), .C1(G311), .C2(new_n784), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n778), .A2(G116), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT46), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n255), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n966), .B2(new_n965), .C1(new_n312), .C2(new_n794), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G294), .B2(new_n800), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n964), .B(new_n969), .C1(new_n830), .C2(new_n799), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n786), .A2(new_n282), .B1(new_n808), .B2(new_n201), .ZN(new_n971));
  INV_X1    g0771(.A(G137), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n805), .A2(new_n972), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(G143), .C2(new_n784), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n347), .B1(new_n775), .B2(G77), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT106), .Z(new_n976));
  INV_X1    g0776(.A(new_n795), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n976), .C1(new_n202), .C2(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G50), .A2(new_n798), .B1(new_n800), .B2(G159), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT105), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n970), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT47), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n764), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n925), .A2(new_n762), .ZN(new_n986));
  INV_X1    g0786(.A(new_n765), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n210), .B2(new_n581), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n210), .A2(new_n255), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n237), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n755), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n985), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n960), .A2(new_n993), .ZN(G387));
  NAND2_X1  g0794(.A1(new_n954), .A2(new_n752), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n746), .A2(new_n954), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n713), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n746), .A2(new_n954), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n234), .A2(G45), .A3(new_n347), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n275), .A2(G50), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1001));
  OAI221_X1 g0801(.A(new_n589), .B1(new_n202), .B2(new_n254), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n347), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n711), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n210), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n987), .B1(G107), .B2(new_n210), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n755), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n789), .A2(G326), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1011), .B(new_n347), .C1(new_n776), .C2(new_n621), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT111), .Z(new_n1013));
  AOI22_X1  g0813(.A1(G317), .A2(new_n787), .B1(new_n784), .B2(G322), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n809), .B2(new_n799), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G311), .B2(new_n800), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT48), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(KEYINPUT48), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n808), .A2(new_n807), .B1(new_n794), .B2(new_n830), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1020), .A2(KEYINPUT49), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(KEYINPUT49), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1013), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n977), .A2(new_n300), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G50), .B2(new_n787), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT109), .Z(new_n1026));
  AOI211_X1 g0826(.A(new_n347), .B(new_n961), .C1(new_n784), .C2(G159), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n202), .B2(new_n799), .C1(new_n275), .C2(new_n801), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n778), .A2(G77), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n805), .B2(new_n282), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT108), .Z(new_n1031));
  NOR3_X1   g0831(.A1(new_n1026), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT110), .Z(new_n1033));
  NAND2_X1  g0833(.A1(new_n1023), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1010), .B1(new_n1034), .B2(new_n764), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT112), .Z(new_n1036));
  NOR2_X1   g0836(.A1(new_n703), .A2(new_n761), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n995), .B1(new_n997), .B2(new_n998), .C1(new_n1036), .C2(new_n1037), .ZN(G393));
  NAND2_X1  g0838(.A1(new_n955), .A2(new_n713), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n946), .A2(new_n948), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n996), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n765), .B1(new_n541), .B2(new_n209), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n247), .B2(new_n989), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n347), .B1(new_n794), .B2(new_n621), .C1(new_n808), .C2(new_n830), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1044), .B(new_n777), .C1(G322), .C2(new_n789), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n812), .A2(new_n786), .B1(new_n783), .B2(new_n962), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G294), .A2(new_n798), .B1(new_n800), .B2(G303), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n255), .B1(new_n808), .B2(new_n202), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1050), .B(new_n834), .C1(G143), .C2(new_n789), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n282), .A2(new_n783), .B1(new_n786), .B2(new_n352), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n795), .A2(G77), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n275), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G50), .A2(new_n800), .B1(new_n798), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT113), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1049), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n755), .B(new_n1043), .C1(new_n1059), .C2(new_n764), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n922), .B2(new_n761), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1040), .B2(new_n751), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1041), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(G390));
  NAND2_X1  g0864(.A1(new_n882), .A2(new_n883), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n823), .A2(new_n698), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n886), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n900), .A2(new_n820), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n904), .B1(new_n1069), .B2(new_n1065), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1070), .A2(new_n906), .A3(new_n907), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n707), .B(new_n822), .C1(new_n734), .C2(new_n740), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n899), .B1(new_n1072), .B2(new_n820), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1073), .A2(new_n880), .A3(new_n904), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1068), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n440), .A2(G330), .A3(new_n886), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n910), .A2(new_n658), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n730), .A2(G330), .A3(new_n824), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n899), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n1067), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1069), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n731), .A2(new_n884), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n886), .A2(new_n1066), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n899), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1082), .A2(new_n820), .A3(new_n1072), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1077), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1072), .A2(new_n820), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n1065), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n904), .B1(new_n871), .B2(new_n879), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n907), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n871), .A2(new_n879), .A3(new_n905), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1090), .B(new_n1082), .C1(new_n1093), .C2(new_n1070), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1075), .A2(new_n1086), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT114), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1075), .A2(new_n1086), .A3(new_n1094), .A4(KEYINPUT114), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n713), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1075), .A2(new_n1094), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1077), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1100), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1099), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT115), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1101), .B2(new_n751), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1075), .A2(new_n1094), .A3(KEYINPUT115), .A4(new_n752), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1091), .A2(new_n758), .A3(new_n1092), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n828), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n819), .B1(new_n1056), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n255), .B(new_n843), .C1(G87), .C2(new_n778), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n805), .A2(new_n807), .B1(new_n621), .B2(new_n786), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G283), .B2(new_n784), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G97), .A2(new_n798), .B1(new_n800), .B2(G107), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1054), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  AOI22_X1  g0918(.A1(new_n798), .A2(new_n1118), .B1(new_n795), .B2(G159), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n972), .B2(new_n801), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n255), .B1(new_n776), .B2(new_n241), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT116), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT53), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n808), .B2(new_n282), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n778), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G132), .A2(new_n787), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n784), .A2(G128), .B1(new_n789), .B2(G125), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1123), .A2(new_n1124), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1117), .B1(new_n1120), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1112), .B1(new_n1131), .B2(new_n764), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT117), .Z(new_n1133));
  AOI22_X1  g0933(.A1(new_n1108), .A2(new_n1109), .B1(new_n1110), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1106), .A2(new_n1134), .ZN(G378));
  OAI21_X1  g0935(.A(new_n819), .B1(G50), .B2(new_n1111), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n787), .A2(G128), .B1(new_n778), .B2(new_n1118), .ZN(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n783), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n799), .A2(new_n972), .B1(new_n977), .B2(new_n282), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(G132), .C2(new_n800), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n277), .B(new_n479), .C1(new_n776), .C2(new_n352), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G124), .B2(new_n789), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n775), .A2(G58), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n312), .B2(new_n786), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n255), .A2(G41), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1029), .B(new_n1150), .C1(new_n783), .C2(new_n621), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G68), .B2(new_n795), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n541), .B2(new_n801), .C1(new_n300), .C2(new_n799), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1149), .B(new_n1153), .C1(G283), .C2(new_n789), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT118), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1147), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n241), .B1(G33), .B2(G41), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1157), .B1(new_n1156), .B2(new_n1155), .C1(new_n1150), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1136), .B1(new_n1159), .B2(new_n764), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n297), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n296), .A2(new_n859), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n657), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n657), .B2(new_n1161), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  OR3_X1    g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n758), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1160), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n698), .B1(new_n888), .B2(new_n894), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1169), .B1(new_n903), .B2(new_n908), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n903), .A2(new_n908), .A3(new_n1169), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1176), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1178), .A2(new_n1174), .A3(new_n1172), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1171), .B1(new_n1180), .B2(new_n751), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1077), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT57), .B1(new_n1186), .B2(new_n1180), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1181), .B1(new_n1188), .B2(new_n713), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G375));
  INV_X1    g0990(.A(new_n938), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1081), .A2(new_n1085), .A3(new_n1077), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1104), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n899), .A2(new_n758), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n789), .A2(G128), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1148), .B(new_n255), .C1(new_n352), .C2(new_n808), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(G137), .C2(new_n787), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n799), .A2(new_n282), .B1(new_n977), .B2(new_n241), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n800), .B2(new_n1118), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n784), .A2(G132), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT120), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1197), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n255), .B1(new_n775), .B2(G77), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT119), .Z(new_n1204));
  OAI22_X1  g1004(.A1(new_n805), .A2(new_n809), .B1(new_n807), .B2(new_n783), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n786), .A2(new_n830), .B1(new_n808), .B2(new_n541), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1024), .B1(new_n798), .B2(G107), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n800), .A2(G116), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1204), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n846), .B1(new_n1202), .B2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n755), .B(new_n1211), .C1(new_n202), .C2(new_n828), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1102), .A2(new_n752), .B1(new_n1194), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1193), .A2(new_n1213), .ZN(G381));
  NAND3_X1  g1014(.A1(new_n960), .A2(new_n993), .A3(new_n1063), .ZN(new_n1215));
  OR2_X1    g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1215), .A2(G384), .A3(new_n1216), .A4(G381), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT121), .Z(new_n1218));
  INV_X1    g1018(.A(KEYINPUT122), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G378), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1106), .A2(new_n1134), .A3(KEYINPUT122), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G375), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1218), .A2(new_n1223), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n692), .A2(G213), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(G407), .A2(G213), .A3(new_n1227), .ZN(G409));
  AOI21_X1  g1028(.A(new_n1183), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1186), .A2(new_n1180), .A3(KEYINPUT57), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n713), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1181), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(G378), .A3(new_n1232), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1106), .A2(new_n1134), .A3(KEYINPUT122), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT122), .B1(new_n1106), .B2(new_n1134), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1186), .A2(new_n1180), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1191), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1232), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1226), .B1(new_n1233), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G384), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1104), .A2(new_n713), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1192), .A2(KEYINPUT60), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1192), .A2(KEYINPUT60), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1213), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1242), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1244), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1192), .A2(KEYINPUT60), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n713), .B(new_n1104), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(G384), .A3(new_n1213), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1248), .A2(new_n1252), .A3(KEYINPUT124), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1255), .A2(G2897), .A3(new_n1226), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1226), .A2(G2897), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1248), .A2(new_n1252), .A3(KEYINPUT124), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT124), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT125), .B1(new_n1241), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1257), .A2(new_n1261), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1189), .A2(G378), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1264), .B(new_n1265), .C1(new_n1266), .C2(new_n1226), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n937), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n959), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n752), .B1(new_n956), .B2(KEYINPUT104), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(G390), .B1(new_n1272), .B2(new_n992), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(G393), .B(G396), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1273), .A2(new_n1215), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1273), .B2(new_n1215), .ZN(new_n1276));
  OR3_X1    g1076(.A1(new_n1275), .A2(new_n1276), .A3(KEYINPUT61), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1226), .B(new_n1253), .C1(new_n1233), .C2(new_n1240), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(KEYINPUT63), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1253), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1100), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1281));
  INV_X1    g1081(.A(G378), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1181), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1181), .B1(new_n1237), .B2(new_n1191), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1222), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1225), .B(new_n1280), .C1(new_n1283), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT123), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1287), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1268), .B(new_n1279), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1265), .B1(new_n1266), .B2(new_n1226), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1233), .A2(new_n1240), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1225), .A4(new_n1280), .ZN(new_n1297));
  XOR2_X1   g1097(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1298));
  NAND3_X1  g1098(.A1(new_n1294), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1278), .A2(new_n1296), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1291), .A2(new_n1301), .ZN(G405));
  OAI21_X1  g1102(.A(new_n1233), .B1(new_n1189), .B2(new_n1222), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1292), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1293), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1280), .A2(KEYINPUT127), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1308), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(G402));
endmodule


