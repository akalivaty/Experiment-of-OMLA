

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U549 ( .A1(G299), .A2(n646), .ZN(n612) );
  NAND2_X1 U550 ( .A1(n702), .A2(n594), .ZN(n657) );
  NOR2_X2 U551 ( .A1(n535), .A2(n534), .ZN(G160) );
  AND2_X1 U552 ( .A1(n637), .A2(G2072), .ZN(n608) );
  INV_X1 U553 ( .A(KEYINPUT97), .ZN(n596) );
  NAND2_X1 U554 ( .A1(n673), .A2(n672), .ZN(n721) );
  NOR2_X2 U555 ( .A1(G2105), .A2(n525), .ZN(n869) );
  NOR2_X1 U556 ( .A1(n542), .A2(G651), .ZN(n782) );
  AND2_X1 U557 ( .A1(G2105), .A2(n525), .ZN(n874) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n746) );
  NOR2_X1 U559 ( .A1(n745), .A2(n744), .ZN(n747) );
  NOR2_X1 U560 ( .A1(G543), .A2(G651), .ZN(n778) );
  NAND2_X1 U561 ( .A1(G91), .A2(n778), .ZN(n514) );
  XNOR2_X1 U562 ( .A(n514), .B(KEYINPUT72), .ZN(n523) );
  XOR2_X1 U563 ( .A(KEYINPUT0), .B(G543), .Z(n542) );
  NAND2_X1 U564 ( .A1(n782), .A2(G53), .ZN(n517) );
  XNOR2_X1 U565 ( .A(KEYINPUT67), .B(G651), .ZN(n518) );
  NOR2_X1 U566 ( .A1(G543), .A2(n518), .ZN(n515) );
  XOR2_X1 U567 ( .A(KEYINPUT1), .B(n515), .Z(n783) );
  NAND2_X1 U568 ( .A1(G65), .A2(n783), .ZN(n516) );
  NAND2_X1 U569 ( .A1(n517), .A2(n516), .ZN(n521) );
  NOR2_X1 U570 ( .A1(n542), .A2(n518), .ZN(n779) );
  NAND2_X1 U571 ( .A1(G78), .A2(n779), .ZN(n519) );
  XNOR2_X1 U572 ( .A(KEYINPUT73), .B(n519), .ZN(n520) );
  NOR2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n523), .A2(n522), .ZN(G299) );
  XOR2_X1 U575 ( .A(KEYINPUT64), .B(G2104), .Z(n525) );
  NAND2_X1 U576 ( .A1(G125), .A2(n874), .ZN(n524) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n524), .Z(n529) );
  NAND2_X1 U578 ( .A1(G101), .A2(n869), .ZN(n527) );
  INV_X1 U579 ( .A(KEYINPUT23), .ZN(n526) );
  XNOR2_X1 U580 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XOR2_X1 U583 ( .A(n530), .B(KEYINPUT66), .Z(n531) );
  XNOR2_X1 U584 ( .A(KEYINPUT17), .B(n531), .ZN(n867) );
  NAND2_X1 U585 ( .A1(G137), .A2(n867), .ZN(n533) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n873) );
  NAND2_X1 U587 ( .A1(n873), .A2(G113), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  AND2_X1 U589 ( .A1(n874), .A2(G126), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G138), .A2(n867), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G114), .A2(n873), .ZN(n537) );
  NAND2_X1 U592 ( .A1(G102), .A2(n869), .ZN(n536) );
  AND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U596 ( .A1(G74), .A2(G651), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G87), .A2(n542), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U599 ( .A1(n783), .A2(n545), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n782), .A2(G49), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(G288) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(KEYINPUT80), .ZN(n560) );
  NAND2_X1 U603 ( .A1(n778), .A2(G89), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G76), .A2(n779), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n551), .B(KEYINPUT5), .ZN(n558) );
  XNOR2_X1 U608 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G63), .A2(n783), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT78), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G51), .A2(n782), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n560), .B(n559), .ZN(G168) );
  NAND2_X1 U616 ( .A1(G64), .A2(n783), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n561), .B(KEYINPUT70), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G52), .A2(n782), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G90), .A2(n778), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G77), .A2(n779), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U623 ( .A(KEYINPUT71), .B(n566), .ZN(n567) );
  XNOR2_X1 U624 ( .A(n567), .B(KEYINPUT9), .ZN(n568) );
  NOR2_X1 U625 ( .A1(n569), .A2(n568), .ZN(G171) );
  XOR2_X1 U626 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U627 ( .A1(G88), .A2(n778), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G75), .A2(n779), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U630 ( .A1(n782), .A2(G50), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G62), .A2(n783), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U633 ( .A1(n575), .A2(n574), .ZN(G166) );
  INV_X1 U634 ( .A(G166), .ZN(G303) );
  NAND2_X1 U635 ( .A1(n778), .A2(G86), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G61), .A2(n783), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U638 ( .A(n578), .B(KEYINPUT89), .ZN(n580) );
  NAND2_X1 U639 ( .A1(G48), .A2(n782), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n779), .A2(G73), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT2), .B(n581), .Z(n582) );
  NOR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U644 ( .A(KEYINPUT90), .B(n584), .Z(G305) );
  NAND2_X1 U645 ( .A1(n779), .A2(G72), .ZN(n585) );
  XNOR2_X1 U646 ( .A(n585), .B(KEYINPUT68), .ZN(n592) );
  NAND2_X1 U647 ( .A1(n778), .A2(G85), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G60), .A2(n783), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G47), .A2(n782), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT69), .B(n588), .ZN(n589) );
  NOR2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U653 ( .A1(n592), .A2(n591), .ZN(G290) );
  NOR2_X1 U654 ( .A1(G164), .A2(G1384), .ZN(n702) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n701) );
  INV_X1 U656 ( .A(n701), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G8), .A2(n657), .ZN(n725) );
  NOR2_X1 U658 ( .A1(G1976), .A2(G288), .ZN(n675) );
  NAND2_X1 U659 ( .A1(n675), .A2(KEYINPUT33), .ZN(n595) );
  NOR2_X1 U660 ( .A1(n725), .A2(n595), .ZN(n683) );
  NOR2_X1 U661 ( .A1(G1966), .A2(n725), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n597), .B(n596), .ZN(n669) );
  NOR2_X1 U663 ( .A1(G2084), .A2(n657), .ZN(n666) );
  NOR2_X1 U664 ( .A1(n669), .A2(n666), .ZN(n598) );
  XOR2_X1 U665 ( .A(n598), .B(KEYINPUT103), .Z(n599) );
  NAND2_X1 U666 ( .A1(G8), .A2(n599), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT30), .ZN(n601) );
  NOR2_X1 U668 ( .A1(n601), .A2(G168), .ZN(n605) );
  XNOR2_X1 U669 ( .A(G2078), .B(KEYINPUT25), .ZN(n933) );
  XNOR2_X1 U670 ( .A(n657), .B(KEYINPUT98), .ZN(n609) );
  INV_X1 U671 ( .A(n609), .ZN(n637) );
  NAND2_X1 U672 ( .A1(n933), .A2(n637), .ZN(n603) );
  INV_X1 U673 ( .A(G1961), .ZN(n984) );
  NAND2_X1 U674 ( .A1(n657), .A2(n984), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n652) );
  NOR2_X1 U676 ( .A1(G171), .A2(n652), .ZN(n604) );
  NOR2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT31), .B(n606), .Z(n656) );
  XOR2_X1 U679 ( .A(KEYINPUT27), .B(KEYINPUT99), .Z(n607) );
  XNOR2_X1 U680 ( .A(n608), .B(n607), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n609), .A2(G1956), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n646) );
  XOR2_X1 U683 ( .A(KEYINPUT102), .B(n612), .Z(n645) );
  NAND2_X1 U684 ( .A1(G92), .A2(n778), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G79), .A2(n779), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n782), .A2(G54), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G66), .A2(n783), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U691 ( .A(KEYINPUT15), .B(n619), .Z(n985) );
  NAND2_X1 U692 ( .A1(n778), .A2(G81), .ZN(n620) );
  XNOR2_X1 U693 ( .A(n620), .B(KEYINPUT12), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G68), .A2(n779), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U696 ( .A(KEYINPUT13), .B(n623), .Z(n627) );
  NAND2_X1 U697 ( .A1(n783), .A2(G56), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(KEYINPUT75), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT14), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n782), .A2(G43), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n992) );
  INV_X1 U703 ( .A(G1996), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n657), .A2(n630), .ZN(n632) );
  XNOR2_X1 U705 ( .A(KEYINPUT26), .B(KEYINPUT101), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n632), .B(n631), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n657), .A2(G1341), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U709 ( .A1(n992), .A2(n635), .ZN(n636) );
  OR2_X1 U710 ( .A1(n985), .A2(n636), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n985), .A2(n636), .ZN(n641) );
  NAND2_X1 U712 ( .A1(G2067), .A2(n637), .ZN(n639) );
  NAND2_X1 U713 ( .A1(G1348), .A2(n657), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n650) );
  NAND2_X1 U718 ( .A1(n646), .A2(G299), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT28), .ZN(n648) );
  XNOR2_X1 U720 ( .A(KEYINPUT100), .B(n648), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT29), .B(n651), .Z(n654) );
  NAND2_X1 U723 ( .A1(G171), .A2(n652), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n667) );
  NAND2_X1 U726 ( .A1(n667), .A2(G286), .ZN(n662) );
  NOR2_X1 U727 ( .A1(G1971), .A2(n725), .ZN(n659) );
  NOR2_X1 U728 ( .A1(G2090), .A2(n657), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U730 ( .A1(n660), .A2(G303), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n663), .B(KEYINPUT104), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n664), .A2(G8), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n665), .B(KEYINPUT32), .ZN(n673) );
  NAND2_X1 U735 ( .A1(G8), .A2(n666), .ZN(n671) );
  INV_X1 U736 ( .A(n667), .ZN(n668) );
  NOR2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U739 ( .A1(G1971), .A2(G303), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n1000) );
  INV_X1 U741 ( .A(KEYINPUT33), .ZN(n676) );
  AND2_X1 U742 ( .A1(n1000), .A2(n676), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n721), .A2(n677), .ZN(n681) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n995) );
  INV_X1 U745 ( .A(n995), .ZN(n678) );
  NOR2_X1 U746 ( .A1(n678), .A2(n725), .ZN(n679) );
  OR2_X1 U747 ( .A1(KEYINPUT33), .A2(n679), .ZN(n680) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n717) );
  XOR2_X1 U750 ( .A(G1981), .B(G305), .Z(n981) );
  XNOR2_X1 U751 ( .A(KEYINPUT93), .B(G1986), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n684), .B(G290), .ZN(n997) );
  NAND2_X1 U753 ( .A1(n873), .A2(G117), .ZN(n686) );
  NAND2_X1 U754 ( .A1(G141), .A2(n867), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n869), .A2(G105), .ZN(n687) );
  XOR2_X1 U757 ( .A(KEYINPUT38), .B(n687), .Z(n688) );
  NOR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n874), .A2(G129), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n863) );
  NAND2_X1 U761 ( .A1(G1996), .A2(n863), .ZN(n692) );
  XOR2_X1 U762 ( .A(KEYINPUT96), .B(n692), .Z(n700) );
  NAND2_X1 U763 ( .A1(n869), .A2(G95), .ZN(n694) );
  NAND2_X1 U764 ( .A1(G131), .A2(n867), .ZN(n693) );
  NAND2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n698) );
  NAND2_X1 U766 ( .A1(G107), .A2(n873), .ZN(n696) );
  NAND2_X1 U767 ( .A1(G119), .A2(n874), .ZN(n695) );
  NAND2_X1 U768 ( .A1(n696), .A2(n695), .ZN(n697) );
  OR2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n860) );
  AND2_X1 U770 ( .A1(n860), .A2(G1991), .ZN(n699) );
  NOR2_X1 U771 ( .A1(n700), .A2(n699), .ZN(n730) );
  NAND2_X1 U772 ( .A1(n997), .A2(n730), .ZN(n703) );
  NOR2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n740) );
  NAND2_X1 U774 ( .A1(n703), .A2(n740), .ZN(n715) );
  XNOR2_X1 U775 ( .A(G2067), .B(KEYINPUT37), .ZN(n737) );
  NAND2_X1 U776 ( .A1(n869), .A2(G104), .ZN(n705) );
  NAND2_X1 U777 ( .A1(G140), .A2(n867), .ZN(n704) );
  NAND2_X1 U778 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U779 ( .A(KEYINPUT34), .B(n706), .ZN(n713) );
  NAND2_X1 U780 ( .A1(n873), .A2(G116), .ZN(n707) );
  XNOR2_X1 U781 ( .A(n707), .B(KEYINPUT94), .ZN(n709) );
  NAND2_X1 U782 ( .A1(G128), .A2(n874), .ZN(n708) );
  NAND2_X1 U783 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U784 ( .A(KEYINPUT35), .B(n710), .ZN(n711) );
  XNOR2_X1 U785 ( .A(KEYINPUT95), .B(n711), .ZN(n712) );
  NOR2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U787 ( .A(KEYINPUT36), .B(n714), .ZN(n880) );
  NOR2_X1 U788 ( .A1(n737), .A2(n880), .ZN(n959) );
  NAND2_X1 U789 ( .A1(n959), .A2(n740), .ZN(n735) );
  AND2_X1 U790 ( .A1(n715), .A2(n735), .ZN(n728) );
  AND2_X1 U791 ( .A1(n981), .A2(n728), .ZN(n716) );
  AND2_X1 U792 ( .A1(n717), .A2(n716), .ZN(n745) );
  NAND2_X1 U793 ( .A1(G8), .A2(G166), .ZN(n718) );
  NOR2_X1 U794 ( .A1(G2090), .A2(n718), .ZN(n719) );
  XNOR2_X1 U795 ( .A(n719), .B(KEYINPUT105), .ZN(n720) );
  NAND2_X1 U796 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U797 ( .A1(n722), .A2(n725), .ZN(n727) );
  NOR2_X1 U798 ( .A1(G1981), .A2(G305), .ZN(n723) );
  XOR2_X1 U799 ( .A(n723), .B(KEYINPUT24), .Z(n724) );
  OR2_X1 U800 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n743) );
  NOR2_X1 U803 ( .A1(G1996), .A2(n863), .ZN(n954) );
  INV_X1 U804 ( .A(n730), .ZN(n958) );
  NOR2_X1 U805 ( .A1(G1986), .A2(G290), .ZN(n731) );
  NOR2_X1 U806 ( .A1(G1991), .A2(n860), .ZN(n961) );
  NOR2_X1 U807 ( .A1(n731), .A2(n961), .ZN(n732) );
  NOR2_X1 U808 ( .A1(n958), .A2(n732), .ZN(n733) );
  NOR2_X1 U809 ( .A1(n954), .A2(n733), .ZN(n734) );
  XNOR2_X1 U810 ( .A(KEYINPUT39), .B(n734), .ZN(n736) );
  NAND2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n737), .A2(n880), .ZN(n956) );
  NAND2_X1 U813 ( .A1(n738), .A2(n956), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U815 ( .A(KEYINPUT106), .B(n741), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U817 ( .A(n747), .B(n746), .ZN(G329) );
  AND2_X1 U818 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U819 ( .A1(G123), .A2(n874), .ZN(n748) );
  XOR2_X1 U820 ( .A(KEYINPUT18), .B(n748), .Z(n749) );
  XNOR2_X1 U821 ( .A(n749), .B(KEYINPUT85), .ZN(n751) );
  NAND2_X1 U822 ( .A1(G135), .A2(n867), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U824 ( .A(KEYINPUT86), .B(n752), .ZN(n755) );
  NAND2_X1 U825 ( .A1(G111), .A2(n873), .ZN(n753) );
  XNOR2_X1 U826 ( .A(KEYINPUT87), .B(n753), .ZN(n754) );
  NOR2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n869), .A2(G99), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n757), .A2(n756), .ZN(n962) );
  XNOR2_X1 U830 ( .A(G2096), .B(n962), .ZN(n758) );
  OR2_X1 U831 ( .A1(G2100), .A2(n758), .ZN(G156) );
  INV_X1 U832 ( .A(G57), .ZN(G237) );
  INV_X1 U833 ( .A(G82), .ZN(G220) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U835 ( .A(n759), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n816) );
  NAND2_X1 U837 ( .A1(n816), .A2(G567), .ZN(n760) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n760), .Z(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n768) );
  OR2_X1 U840 ( .A1(n992), .A2(n768), .ZN(n761) );
  XNOR2_X1 U841 ( .A(KEYINPUT76), .B(n761), .ZN(G153) );
  INV_X1 U842 ( .A(G171), .ZN(G301) );
  NOR2_X1 U843 ( .A1(n985), .A2(G868), .ZN(n762) );
  XNOR2_X1 U844 ( .A(n762), .B(KEYINPUT77), .ZN(n764) );
  NAND2_X1 U845 ( .A1(G868), .A2(G301), .ZN(n763) );
  NAND2_X1 U846 ( .A1(n764), .A2(n763), .ZN(G284) );
  INV_X1 U847 ( .A(G868), .ZN(n799) );
  NAND2_X1 U848 ( .A1(G299), .A2(n799), .ZN(n766) );
  NAND2_X1 U849 ( .A1(G868), .A2(G286), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U851 ( .A(KEYINPUT81), .B(n767), .Z(G297) );
  NAND2_X1 U852 ( .A1(n768), .A2(G559), .ZN(n769) );
  NAND2_X1 U853 ( .A1(n769), .A2(n985), .ZN(n770) );
  XNOR2_X1 U854 ( .A(n770), .B(KEYINPUT16), .ZN(n771) );
  XNOR2_X1 U855 ( .A(KEYINPUT82), .B(n771), .ZN(G148) );
  NOR2_X1 U856 ( .A1(G868), .A2(n992), .ZN(n772) );
  XOR2_X1 U857 ( .A(KEYINPUT83), .B(n772), .Z(n775) );
  NAND2_X1 U858 ( .A1(G868), .A2(n985), .ZN(n773) );
  NOR2_X1 U859 ( .A1(G559), .A2(n773), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U861 ( .A(KEYINPUT84), .B(n776), .ZN(G282) );
  NAND2_X1 U862 ( .A1(n985), .A2(G559), .ZN(n797) );
  XNOR2_X1 U863 ( .A(n992), .B(n797), .ZN(n777) );
  NOR2_X1 U864 ( .A1(G860), .A2(n777), .ZN(n789) );
  NAND2_X1 U865 ( .A1(G93), .A2(n778), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G80), .A2(n779), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n787) );
  NAND2_X1 U868 ( .A1(n782), .A2(G55), .ZN(n785) );
  NAND2_X1 U869 ( .A1(G67), .A2(n783), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n800) );
  XOR2_X1 U872 ( .A(n800), .B(KEYINPUT88), .Z(n788) );
  XNOR2_X1 U873 ( .A(n789), .B(n788), .ZN(G145) );
  XNOR2_X1 U874 ( .A(KEYINPUT91), .B(KEYINPUT19), .ZN(n791) );
  XNOR2_X1 U875 ( .A(G299), .B(G166), .ZN(n790) );
  XNOR2_X1 U876 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U877 ( .A(n792), .B(G288), .ZN(n794) );
  XNOR2_X1 U878 ( .A(n800), .B(G290), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n794), .B(n793), .ZN(n795) );
  XNOR2_X1 U880 ( .A(G305), .B(n795), .ZN(n796) );
  XNOR2_X1 U881 ( .A(n796), .B(n992), .ZN(n887) );
  XOR2_X1 U882 ( .A(n887), .B(n797), .Z(n798) );
  NOR2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n802) );
  NOR2_X1 U884 ( .A1(G868), .A2(n800), .ZN(n801) );
  NOR2_X1 U885 ( .A1(n802), .A2(n801), .ZN(G295) );
  NAND2_X1 U886 ( .A1(G2078), .A2(G2084), .ZN(n803) );
  XOR2_X1 U887 ( .A(KEYINPUT20), .B(n803), .Z(n804) );
  NAND2_X1 U888 ( .A1(G2090), .A2(n804), .ZN(n805) );
  XNOR2_X1 U889 ( .A(KEYINPUT21), .B(n805), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n806), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U891 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U892 ( .A(KEYINPUT74), .B(G132), .Z(G219) );
  NOR2_X1 U893 ( .A1(G219), .A2(G220), .ZN(n807) );
  XOR2_X1 U894 ( .A(KEYINPUT22), .B(n807), .Z(n808) );
  XNOR2_X1 U895 ( .A(n808), .B(KEYINPUT92), .ZN(n809) );
  NOR2_X1 U896 ( .A1(G218), .A2(n809), .ZN(n810) );
  NAND2_X1 U897 ( .A1(G96), .A2(n810), .ZN(n820) );
  NAND2_X1 U898 ( .A1(n820), .A2(G2106), .ZN(n814) );
  NAND2_X1 U899 ( .A1(G69), .A2(G120), .ZN(n811) );
  NOR2_X1 U900 ( .A1(G237), .A2(n811), .ZN(n812) );
  NAND2_X1 U901 ( .A1(G108), .A2(n812), .ZN(n821) );
  NAND2_X1 U902 ( .A1(n821), .A2(G567), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n814), .A2(n813), .ZN(n822) );
  NAND2_X1 U904 ( .A1(G483), .A2(G661), .ZN(n815) );
  NOR2_X1 U905 ( .A1(n822), .A2(n815), .ZN(n819) );
  NAND2_X1 U906 ( .A1(n819), .A2(G36), .ZN(G176) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U909 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(G188) );
  XNOR2_X1 U912 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G69), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  INV_X1 U918 ( .A(n822), .ZN(G319) );
  XOR2_X1 U919 ( .A(KEYINPUT41), .B(G1991), .Z(n824) );
  XNOR2_X1 U920 ( .A(G1966), .B(G1996), .ZN(n823) );
  XNOR2_X1 U921 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U922 ( .A(n825), .B(KEYINPUT111), .Z(n827) );
  XNOR2_X1 U923 ( .A(G1971), .B(G1986), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U925 ( .A(G1976), .B(G1981), .Z(n829) );
  XNOR2_X1 U926 ( .A(G1961), .B(G1956), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U929 ( .A(KEYINPUT112), .B(G2474), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(G229) );
  XOR2_X1 U931 ( .A(G2096), .B(KEYINPUT43), .Z(n835) );
  XNOR2_X1 U932 ( .A(G2090), .B(KEYINPUT110), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n836), .B(G2678), .Z(n838) );
  XNOR2_X1 U935 ( .A(G2072), .B(G2067), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U937 ( .A(KEYINPUT42), .B(G2100), .Z(n840) );
  XNOR2_X1 U938 ( .A(G2078), .B(G2084), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(G227) );
  NAND2_X1 U941 ( .A1(n873), .A2(G112), .ZN(n844) );
  NAND2_X1 U942 ( .A1(G136), .A2(n867), .ZN(n843) );
  NAND2_X1 U943 ( .A1(n844), .A2(n843), .ZN(n850) );
  NAND2_X1 U944 ( .A1(G124), .A2(n874), .ZN(n845) );
  XOR2_X1 U945 ( .A(KEYINPUT44), .B(n845), .Z(n846) );
  XNOR2_X1 U946 ( .A(n846), .B(KEYINPUT113), .ZN(n848) );
  NAND2_X1 U947 ( .A1(G100), .A2(n869), .ZN(n847) );
  NAND2_X1 U948 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U949 ( .A1(n850), .A2(n849), .ZN(G162) );
  NAND2_X1 U950 ( .A1(n869), .A2(G106), .ZN(n851) );
  XOR2_X1 U951 ( .A(KEYINPUT115), .B(n851), .Z(n853) );
  NAND2_X1 U952 ( .A1(G142), .A2(n867), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n854), .B(KEYINPUT45), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G118), .A2(n873), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n874), .A2(G130), .ZN(n857) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(n857), .Z(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n866) );
  XOR2_X1 U960 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n862) );
  XOR2_X1 U961 ( .A(G164), .B(n860), .Z(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n882) );
  NAND2_X1 U965 ( .A1(G139), .A2(n867), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n868), .B(KEYINPUT116), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G103), .A2(n869), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U969 ( .A(KEYINPUT117), .B(n872), .Z(n879) );
  NAND2_X1 U970 ( .A1(G115), .A2(n873), .ZN(n876) );
  NAND2_X1 U971 ( .A1(G127), .A2(n874), .ZN(n875) );
  NAND2_X1 U972 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n964) );
  XNOR2_X1 U975 ( .A(n880), .B(n964), .ZN(n881) );
  XNOR2_X1 U976 ( .A(n882), .B(n881), .ZN(n885) );
  XNOR2_X1 U977 ( .A(G160), .B(G162), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n883), .B(n962), .ZN(n884) );
  XOR2_X1 U979 ( .A(n885), .B(n884), .Z(n886) );
  NOR2_X1 U980 ( .A1(G37), .A2(n886), .ZN(G395) );
  XNOR2_X1 U981 ( .A(n985), .B(G286), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U983 ( .A(n889), .B(G171), .ZN(n890) );
  NOR2_X1 U984 ( .A1(G37), .A2(n890), .ZN(G397) );
  XOR2_X1 U985 ( .A(G2451), .B(G2443), .Z(n892) );
  XNOR2_X1 U986 ( .A(G2427), .B(G2454), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U988 ( .A(n893), .B(G2446), .Z(n895) );
  XNOR2_X1 U989 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U991 ( .A(G2435), .B(KEYINPUT108), .Z(n897) );
  XNOR2_X1 U992 ( .A(G2430), .B(G2438), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(n899), .B(n898), .Z(n900) );
  NAND2_X1 U995 ( .A1(G14), .A2(n900), .ZN(n906) );
  NAND2_X1 U996 ( .A1(G319), .A2(n906), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n901) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  INV_X1 U1004 ( .A(n906), .ZN(G401) );
  XNOR2_X1 U1005 ( .A(G1986), .B(G24), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(G1971), .B(G22), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(G1976), .B(G23), .ZN(n907) );
  NOR2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(KEYINPUT127), .B(n909), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT58), .B(n912), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(G1966), .B(G21), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(G1961), .B(G5), .ZN(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n926) );
  XOR2_X1 U1016 ( .A(G1348), .B(KEYINPUT59), .Z(n917) );
  XNOR2_X1 U1017 ( .A(G4), .B(n917), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(G20), .B(G1956), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(G1341), .B(G19), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(G1981), .B(G6), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT60), .B(n924), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1026 ( .A(KEYINPUT61), .B(n927), .Z(n928) );
  NOR2_X1 U1027 ( .A1(G16), .A2(n928), .ZN(n951) );
  XOR2_X1 U1028 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n976) );
  XOR2_X1 U1029 ( .A(G2084), .B(G34), .Z(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT54), .B(n929), .ZN(n944) );
  XNOR2_X1 U1031 ( .A(G2090), .B(G35), .ZN(n942) );
  XOR2_X1 U1032 ( .A(G25), .B(G1991), .Z(n930) );
  NAND2_X1 U1033 ( .A1(n930), .A2(G28), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(G2072), .B(G33), .ZN(n932) );
  XNOR2_X1 U1035 ( .A(G1996), .B(G32), .ZN(n931) );
  NOR2_X1 U1036 ( .A1(n932), .A2(n931), .ZN(n937) );
  XOR2_X1 U1037 ( .A(n933), .B(G27), .Z(n935) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n934) );
  NOR2_X1 U1039 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1040 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1041 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(KEYINPUT53), .B(n940), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(n945), .B(KEYINPUT121), .ZN(n946) );
  XOR2_X1 U1046 ( .A(n976), .B(n946), .Z(n948) );
  INV_X1 U1047 ( .A(G29), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n949), .A2(G11), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n980) );
  XOR2_X1 U1051 ( .A(G2090), .B(G162), .Z(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT118), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1054 ( .A(KEYINPUT51), .B(n955), .Z(n957) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n974) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n972) );
  XOR2_X1 U1057 ( .A(G2084), .B(G160), .Z(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G2072), .B(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G164), .B(G2078), .ZN(n965) );
  NAND2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1063 ( .A(KEYINPUT119), .B(n967), .Z(n968) );
  XNOR2_X1 U1064 ( .A(KEYINPUT50), .B(n968), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(KEYINPUT52), .B(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n978), .A2(G29), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n1011) );
  XOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .Z(n1009) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(KEYINPUT57), .B(n983), .ZN(n991) );
  XNOR2_X1 U1076 ( .A(G301), .B(n984), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n985), .B(G1348), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n986), .B(KEYINPUT122), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT123), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n1006) );
  XNOR2_X1 U1082 ( .A(n992), .B(G1341), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT125), .ZN(n1004) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n999) );
  XOR2_X1 U1086 ( .A(G1956), .B(G299), .Z(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(KEYINPUT124), .B(n1002), .Z(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(KEYINPUT126), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1095 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1012), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1097 ( .A(G311), .ZN(G150) );
endmodule

