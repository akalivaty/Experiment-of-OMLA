

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X2 U559 ( .A1(n750), .A2(n720), .ZN(n722) );
  XNOR2_X1 U560 ( .A(n595), .B(n594), .ZN(n894) );
  NOR2_X2 U561 ( .A1(n694), .A2(n797), .ZN(n729) );
  XOR2_X1 U562 ( .A(KEYINPUT0), .B(G543), .Z(n653) );
  XNOR2_X1 U563 ( .A(KEYINPUT64), .B(n530), .ZN(n658) );
  OR2_X1 U564 ( .A1(n894), .A2(n716), .ZN(n936) );
  INV_X1 U565 ( .A(KEYINPUT70), .ZN(n594) );
  INV_X1 U566 ( .A(G651), .ZN(n532) );
  AND2_X2 U567 ( .A1(n546), .A2(G2104), .ZN(n866) );
  NOR2_X1 U568 ( .A1(n551), .A2(n550), .ZN(G160) );
  NOR2_X1 U569 ( .A1(G543), .A2(G651), .ZN(n641) );
  NAND2_X1 U570 ( .A1(G89), .A2(n641), .ZN(n525) );
  XOR2_X1 U571 ( .A(KEYINPUT4), .B(n525), .Z(n526) );
  XNOR2_X1 U572 ( .A(n526), .B(KEYINPUT73), .ZN(n528) );
  NOR2_X1 U573 ( .A1(n653), .A2(n532), .ZN(n645) );
  NAND2_X1 U574 ( .A1(G76), .A2(n645), .ZN(n527) );
  NAND2_X1 U575 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n529), .B(KEYINPUT5), .ZN(n540) );
  XNOR2_X1 U577 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n538) );
  NOR2_X1 U578 ( .A1(n653), .A2(G651), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G51), .A2(n658), .ZN(n531) );
  XNOR2_X1 U580 ( .A(n531), .B(KEYINPUT74), .ZN(n536) );
  NOR2_X1 U581 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n533), .Z(n534) );
  XNOR2_X2 U583 ( .A(KEYINPUT66), .B(n534), .ZN(n657) );
  NAND2_X1 U584 ( .A1(G63), .A2(n657), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U586 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U587 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U588 ( .A(KEYINPUT7), .B(n541), .Z(n948) );
  XNOR2_X1 U589 ( .A(n948), .B(KEYINPUT8), .ZN(G286) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n870) );
  NAND2_X1 U591 ( .A1(G113), .A2(n870), .ZN(n544) );
  NOR2_X1 U592 ( .A1(G2105), .A2(G2104), .ZN(n542) );
  XOR2_X1 U593 ( .A(KEYINPUT17), .B(n542), .Z(n867) );
  NAND2_X1 U594 ( .A1(G137), .A2(n867), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n544), .A2(n543), .ZN(n551) );
  INV_X1 U596 ( .A(G2105), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n866), .A2(G101), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(n545), .Z(n548) );
  NOR2_X1 U599 ( .A1(G2104), .A2(n546), .ZN(n871) );
  NAND2_X1 U600 ( .A1(n871), .A2(G125), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U602 ( .A(KEYINPUT65), .B(n549), .Z(n550) );
  NAND2_X1 U603 ( .A1(G85), .A2(n641), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G72), .A2(n645), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U606 ( .A1(G60), .A2(n657), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G47), .A2(n658), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n556) );
  OR2_X1 U609 ( .A1(n557), .A2(n556), .ZN(G290) );
  XNOR2_X1 U610 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U611 ( .A(G2435), .B(G2427), .Z(n559) );
  XNOR2_X1 U612 ( .A(G2446), .B(G2454), .ZN(n558) );
  XNOR2_X1 U613 ( .A(n559), .B(n558), .ZN(n565) );
  XOR2_X1 U614 ( .A(G2451), .B(G2430), .Z(n561) );
  XNOR2_X1 U615 ( .A(G1348), .B(G1341), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U617 ( .A(G2438), .B(G2443), .Z(n562) );
  XNOR2_X1 U618 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U619 ( .A(n565), .B(n564), .Z(n566) );
  AND2_X1 U620 ( .A1(G14), .A2(n566), .ZN(G401) );
  AND2_X1 U621 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  NAND2_X1 U625 ( .A1(G90), .A2(n641), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G77), .A2(n645), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U628 ( .A(KEYINPUT9), .B(n569), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n657), .A2(G64), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n658), .A2(G52), .ZN(n570) );
  AND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n574) );
  XOR2_X1 U634 ( .A(n574), .B(KEYINPUT10), .Z(n928) );
  NAND2_X1 U635 ( .A1(n928), .A2(G567), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U637 ( .A1(n657), .A2(G56), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n576), .Z(n583) );
  NAND2_X1 U639 ( .A1(G81), .A2(n641), .ZN(n577) );
  XNOR2_X1 U640 ( .A(n577), .B(KEYINPUT12), .ZN(n578) );
  XNOR2_X1 U641 ( .A(n578), .B(KEYINPUT68), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G68), .A2(n645), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G43), .A2(n658), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(n932) );
  INV_X1 U648 ( .A(G860), .ZN(n609) );
  OR2_X1 U649 ( .A1(n932), .A2(n609), .ZN(G153) );
  NAND2_X1 U650 ( .A1(G54), .A2(n658), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n645), .A2(G79), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G66), .A2(n657), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U654 ( .A1(G92), .A2(n641), .ZN(n588) );
  XNOR2_X1 U655 ( .A(KEYINPUT69), .B(n588), .ZN(n589) );
  NOR2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n593), .Z(n595) );
  NOR2_X1 U659 ( .A1(G868), .A2(n894), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(KEYINPUT71), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(n599), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n641), .ZN(n601) );
  NAND2_X1 U665 ( .A1(G78), .A2(n645), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U667 ( .A1(G65), .A2(n657), .ZN(n602) );
  XNOR2_X1 U668 ( .A(KEYINPUT67), .B(n602), .ZN(n603) );
  NOR2_X1 U669 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U670 ( .A1(G53), .A2(n658), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n606), .A2(n605), .ZN(G299) );
  INV_X1 U672 ( .A(G868), .ZN(n668) );
  NOR2_X1 U673 ( .A1(G286), .A2(n668), .ZN(n608) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U675 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n610), .A2(n894), .ZN(n611) );
  XNOR2_X1 U678 ( .A(n611), .B(KEYINPUT76), .ZN(n612) );
  XNOR2_X1 U679 ( .A(KEYINPUT16), .B(n612), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n932), .ZN(n615) );
  NAND2_X1 U681 ( .A1(n894), .A2(G868), .ZN(n613) );
  NOR2_X1 U682 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U683 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G99), .A2(n866), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G111), .A2(n870), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n623) );
  NAND2_X1 U687 ( .A1(n871), .A2(G123), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n618), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U689 ( .A1(G135), .A2(n867), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U691 ( .A(KEYINPUT77), .B(n621), .Z(n622) );
  NOR2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n1010) );
  XOR2_X1 U693 ( .A(G2096), .B(n1010), .Z(n624) );
  NOR2_X1 U694 ( .A1(G2100), .A2(n624), .ZN(n625) );
  XOR2_X1 U695 ( .A(KEYINPUT78), .B(n625), .Z(G156) );
  NAND2_X1 U696 ( .A1(n641), .A2(G93), .ZN(n627) );
  NAND2_X1 U697 ( .A1(G67), .A2(n657), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U699 ( .A1(G80), .A2(n645), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G55), .A2(n658), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n669) );
  NAND2_X1 U703 ( .A1(n894), .A2(G559), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n632), .B(n932), .ZN(n666) );
  XOR2_X1 U705 ( .A(KEYINPUT79), .B(n666), .Z(n633) );
  NOR2_X1 U706 ( .A1(G860), .A2(n633), .ZN(n634) );
  XOR2_X1 U707 ( .A(n669), .B(n634), .Z(G145) );
  NAND2_X1 U708 ( .A1(G88), .A2(n641), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G75), .A2(n645), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U711 ( .A1(G62), .A2(n657), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G50), .A2(n658), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(G166) );
  NAND2_X1 U715 ( .A1(n641), .A2(G86), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n642), .B(KEYINPUT80), .ZN(n644) );
  NAND2_X1 U717 ( .A1(G61), .A2(n657), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n649) );
  NAND2_X1 U719 ( .A1(G73), .A2(n645), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT81), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(KEYINPUT2), .ZN(n648) );
  NOR2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(KEYINPUT82), .ZN(n652) );
  NAND2_X1 U724 ( .A1(G48), .A2(n658), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G87), .A2(n653), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U730 ( .A1(G49), .A2(n658), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(G288) );
  XNOR2_X1 U732 ( .A(G166), .B(G290), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n669), .B(G299), .ZN(n661) );
  XNOR2_X1 U734 ( .A(G305), .B(n661), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(n664), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(G288), .ZN(n895) );
  XNOR2_X1 U738 ( .A(n666), .B(n895), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U746 ( .A1(n675), .A2(G2072), .ZN(G158) );
  NAND2_X1 U747 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U748 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U749 ( .A1(G108), .A2(n677), .ZN(n849) );
  NAND2_X1 U750 ( .A1(G567), .A2(n849), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n678), .B(KEYINPUT83), .ZN(n683) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n679) );
  XNOR2_X1 U753 ( .A(KEYINPUT22), .B(n679), .ZN(n680) );
  NAND2_X1 U754 ( .A1(n680), .A2(G96), .ZN(n681) );
  OR2_X1 U755 ( .A1(G218), .A2(n681), .ZN(n850) );
  AND2_X1 U756 ( .A1(G2106), .A2(n850), .ZN(n682) );
  NOR2_X1 U757 ( .A1(n683), .A2(n682), .ZN(G319) );
  INV_X1 U758 ( .A(G319), .ZN(n686) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n684) );
  XNOR2_X1 U760 ( .A(KEYINPUT84), .B(n684), .ZN(n685) );
  NOR2_X1 U761 ( .A1(n686), .A2(n685), .ZN(n848) );
  NAND2_X1 U762 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U763 ( .A1(n870), .A2(G114), .ZN(n689) );
  NAND2_X1 U764 ( .A1(G102), .A2(n866), .ZN(n687) );
  XOR2_X1 U765 ( .A(KEYINPUT85), .B(n687), .Z(n688) );
  NAND2_X1 U766 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U767 ( .A1(G138), .A2(n867), .ZN(n691) );
  NAND2_X1 U768 ( .A1(G126), .A2(n871), .ZN(n690) );
  NAND2_X1 U769 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U770 ( .A1(n693), .A2(n692), .ZN(G164) );
  XOR2_X1 U771 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n798) );
  INV_X1 U773 ( .A(n798), .ZN(n694) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n797) );
  INV_X1 U775 ( .A(n729), .ZN(n750) );
  NAND2_X1 U776 ( .A1(G8), .A2(n750), .ZN(n787) );
  NOR2_X1 U777 ( .A1(G1966), .A2(n787), .ZN(n759) );
  NOR2_X1 U778 ( .A1(G2084), .A2(n750), .ZN(n760) );
  NOR2_X1 U779 ( .A1(n759), .A2(n760), .ZN(n695) );
  NAND2_X1 U780 ( .A1(G8), .A2(n695), .ZN(n696) );
  XNOR2_X1 U781 ( .A(KEYINPUT99), .B(n696), .ZN(n697) );
  XNOR2_X1 U782 ( .A(n697), .B(KEYINPUT30), .ZN(n698) );
  NAND2_X1 U783 ( .A1(n698), .A2(n948), .ZN(n708) );
  XOR2_X1 U784 ( .A(G2078), .B(KEYINPUT25), .Z(n983) );
  NOR2_X1 U785 ( .A1(n750), .A2(n983), .ZN(n699) );
  XNOR2_X1 U786 ( .A(n699), .B(KEYINPUT93), .ZN(n703) );
  INV_X1 U787 ( .A(KEYINPUT92), .ZN(n700) );
  NOR2_X1 U788 ( .A1(G1961), .A2(n700), .ZN(n701) );
  NAND2_X1 U789 ( .A1(n750), .A2(n701), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U791 ( .A1(G1961), .A2(n729), .ZN(n704) );
  NOR2_X1 U792 ( .A1(KEYINPUT92), .A2(n704), .ZN(n705) );
  NOR2_X1 U793 ( .A1(n706), .A2(n705), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(G301), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n710) );
  XOR2_X1 U796 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n709) );
  XNOR2_X1 U797 ( .A(n710), .B(n709), .ZN(n748) );
  NAND2_X1 U798 ( .A1(G1956), .A2(n750), .ZN(n711) );
  XNOR2_X1 U799 ( .A(KEYINPUT94), .B(n711), .ZN(n714) );
  NAND2_X1 U800 ( .A1(n729), .A2(G2072), .ZN(n712) );
  XOR2_X1 U801 ( .A(KEYINPUT27), .B(n712), .Z(n713) );
  NAND2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n736) );
  NAND2_X1 U803 ( .A1(G299), .A2(n736), .ZN(n715) );
  XNOR2_X1 U804 ( .A(KEYINPUT28), .B(n715), .ZN(n742) );
  INV_X1 U805 ( .A(G1348), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n936), .A2(KEYINPUT26), .ZN(n717) );
  NOR2_X1 U807 ( .A1(G1341), .A2(n717), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n729), .A2(n718), .ZN(n728) );
  INV_X1 U809 ( .A(n894), .ZN(n929) );
  AND2_X1 U810 ( .A1(G2067), .A2(n729), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n929), .A2(n719), .ZN(n724) );
  XOR2_X1 U812 ( .A(G1996), .B(KEYINPUT95), .Z(n993) );
  NAND2_X1 U813 ( .A1(KEYINPUT26), .A2(n993), .ZN(n720) );
  OR2_X1 U814 ( .A1(KEYINPUT26), .A2(n993), .ZN(n721) );
  AND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n723) );
  AND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n726) );
  INV_X1 U817 ( .A(n932), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n734) );
  NAND2_X1 U820 ( .A1(G1348), .A2(n750), .ZN(n731) );
  NAND2_X1 U821 ( .A1(G2067), .A2(n729), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U823 ( .A1(n732), .A2(n929), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U825 ( .A(KEYINPUT96), .B(n735), .ZN(n739) );
  NOR2_X1 U826 ( .A1(G299), .A2(n736), .ZN(n737) );
  XNOR2_X1 U827 ( .A(KEYINPUT97), .B(n737), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U829 ( .A(KEYINPUT98), .B(n740), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U831 ( .A(n743), .B(KEYINPUT29), .ZN(n746) );
  NOR2_X1 U832 ( .A1(G301), .A2(n744), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n758) );
  INV_X1 U835 ( .A(n758), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n749), .A2(G286), .ZN(n755) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n787), .ZN(n752) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n750), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n753), .A2(G303), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n756), .A2(G8), .ZN(n757) );
  XNOR2_X1 U843 ( .A(KEYINPUT32), .B(n757), .ZN(n765) );
  NOR2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U845 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U847 ( .A(KEYINPUT101), .B(n763), .Z(n764) );
  NAND2_X1 U848 ( .A1(n765), .A2(n764), .ZN(n772) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n766) );
  NAND2_X1 U850 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U851 ( .A1(n772), .A2(n767), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n768), .A2(n787), .ZN(n783) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n775) );
  NOR2_X1 U854 ( .A1(G303), .A2(G1971), .ZN(n769) );
  NOR2_X1 U855 ( .A1(n775), .A2(n769), .ZN(n938) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n770) );
  AND2_X1 U857 ( .A1(n938), .A2(n770), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n781) );
  INV_X1 U859 ( .A(n787), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n942) );
  AND2_X1 U861 ( .A1(n773), .A2(n942), .ZN(n774) );
  NOR2_X1 U862 ( .A1(KEYINPUT33), .A2(n774), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n775), .A2(KEYINPUT33), .ZN(n776) );
  NOR2_X1 U864 ( .A1(n776), .A2(n787), .ZN(n777) );
  NOR2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U866 ( .A(G1981), .B(G305), .Z(n949) );
  AND2_X1 U867 ( .A1(n779), .A2(n949), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n832) );
  NOR2_X1 U870 ( .A1(G1981), .A2(G305), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(KEYINPUT91), .ZN(n785) );
  XNOR2_X1 U872 ( .A(KEYINPUT24), .B(n785), .ZN(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n830) );
  NAND2_X1 U874 ( .A1(G104), .A2(n866), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G140), .A2(n867), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n790), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G116), .A2(n870), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G128), .A2(n871), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U883 ( .A(KEYINPUT36), .B(n796), .Z(n890) );
  XOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .Z(n799) );
  OR2_X1 U885 ( .A1(n890), .A2(n799), .ZN(n1030) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n833) );
  NAND2_X1 U887 ( .A1(n799), .A2(n890), .ZN(n800) );
  XNOR2_X1 U888 ( .A(n800), .B(KEYINPUT87), .ZN(n1014) );
  NAND2_X1 U889 ( .A1(n833), .A2(n1014), .ZN(n835) );
  XOR2_X1 U890 ( .A(KEYINPUT39), .B(KEYINPUT102), .Z(n825) );
  NAND2_X1 U891 ( .A1(G105), .A2(n866), .ZN(n801) );
  XNOR2_X1 U892 ( .A(n801), .B(KEYINPUT38), .ZN(n808) );
  NAND2_X1 U893 ( .A1(G117), .A2(n870), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G141), .A2(n867), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U896 ( .A1(G129), .A2(n871), .ZN(n804) );
  XNOR2_X1 U897 ( .A(KEYINPUT89), .B(n804), .ZN(n805) );
  NOR2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n881) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n881), .ZN(n1028) );
  NAND2_X1 U901 ( .A1(G1996), .A2(n881), .ZN(n809) );
  XOR2_X1 U902 ( .A(KEYINPUT90), .B(n809), .Z(n818) );
  NAND2_X1 U903 ( .A1(G107), .A2(n870), .ZN(n811) );
  NAND2_X1 U904 ( .A1(G119), .A2(n871), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U906 ( .A(KEYINPUT88), .B(n812), .ZN(n816) );
  NAND2_X1 U907 ( .A1(G95), .A2(n866), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G131), .A2(n867), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  OR2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n886) );
  AND2_X1 U911 ( .A1(n886), .A2(G1991), .ZN(n817) );
  NOR2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n1016) );
  INV_X1 U913 ( .A(n1016), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n833), .ZN(n834) );
  INV_X1 U915 ( .A(n834), .ZN(n822) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n886), .ZN(n1011) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n1011), .A2(n820), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n1028), .A2(n823), .ZN(n824) );
  XOR2_X1 U921 ( .A(n825), .B(n824), .Z(n826) );
  NAND2_X1 U922 ( .A1(n835), .A2(n826), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n1030), .A2(n827), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n828), .A2(n833), .ZN(n839) );
  INV_X1 U925 ( .A(n839), .ZN(n829) );
  OR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n841) );
  XNOR2_X1 U928 ( .A(G1986), .B(G290), .ZN(n934) );
  AND2_X1 U929 ( .A1(n934), .A2(n833), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n836) );
  OR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(n838) );
  AND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(n840) );
  NOR2_X1 U933 ( .A1(n841), .A2(n840), .ZN(n843) );
  XOR2_X1 U934 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n842) );
  XNOR2_X1 U935 ( .A(n843), .B(n842), .ZN(G329) );
  INV_X1 U936 ( .A(n948), .ZN(G168) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n928), .ZN(G217) );
  INV_X1 U938 ( .A(G661), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G2), .A2(G15), .ZN(n844) );
  NOR2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U941 ( .A(KEYINPUT104), .B(n846), .Z(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U943 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  INV_X1 U947 ( .A(G69), .ZN(G235) );
  NOR2_X1 U948 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  NAND2_X1 U950 ( .A1(G124), .A2(n871), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n866), .A2(G100), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U954 ( .A1(G112), .A2(n870), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G136), .A2(n867), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U957 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U958 ( .A1(G106), .A2(n866), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G142), .A2(n867), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(KEYINPUT45), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G118), .A2(n870), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n871), .A2(G130), .ZN(n863) );
  XOR2_X1 U965 ( .A(KEYINPUT108), .B(n863), .Z(n864) );
  NOR2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n885) );
  NAND2_X1 U967 ( .A1(G103), .A2(n866), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G139), .A2(n867), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G115), .A2(n870), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G127), .A2(n871), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(n874), .ZN(n875) );
  XNOR2_X1 U974 ( .A(KEYINPUT47), .B(n875), .ZN(n876) );
  NOR2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n1020) );
  XOR2_X1 U976 ( .A(KEYINPUT110), .B(KEYINPUT48), .Z(n879) );
  XNOR2_X1 U977 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n1020), .B(n880), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n881), .B(G162), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U982 ( .A(n885), .B(n884), .Z(n888) );
  XOR2_X1 U983 ( .A(G164), .B(n886), .Z(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(n1010), .Z(n892) );
  XNOR2_X1 U986 ( .A(G160), .B(n890), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U988 ( .A1(G37), .A2(n893), .ZN(G395) );
  XOR2_X1 U989 ( .A(n894), .B(n932), .Z(n896) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U991 ( .A(n897), .B(KEYINPUT113), .Z(n899) );
  XOR2_X1 U992 ( .A(G301), .B(KEYINPUT112), .Z(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(G286), .ZN(n901) );
  NOR2_X1 U995 ( .A1(G37), .A2(n901), .ZN(G397) );
  XOR2_X1 U996 ( .A(G1976), .B(G1981), .Z(n903) );
  XNOR2_X1 U997 ( .A(G1956), .B(G1971), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U999 ( .A(G1961), .B(G1966), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G1996), .B(G1991), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1002 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1003 ( .A(KEYINPUT107), .B(G2474), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1005 ( .A(G1986), .B(KEYINPUT41), .Z(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(G229) );
  XOR2_X1 U1007 ( .A(KEYINPUT43), .B(G2678), .Z(n913) );
  XNOR2_X1 U1008 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n917) );
  XOR2_X1 U1010 ( .A(KEYINPUT42), .B(G2090), .Z(n915) );
  XNOR2_X1 U1011 ( .A(G2067), .B(G2072), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(n917), .B(n916), .Z(n919) );
  XNOR2_X1 U1014 ( .A(G2096), .B(G2100), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n921) );
  XOR2_X1 U1016 ( .A(G2084), .B(G2078), .Z(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(G227) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n922) );
  XNOR2_X1 U1019 ( .A(n922), .B(KEYINPUT114), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n923), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G401), .A2(n924), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(G229), .A2(G227), .ZN(n925) );
  XOR2_X1 U1023 ( .A(KEYINPUT49), .B(n925), .Z(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  INV_X1 U1027 ( .A(n928), .ZN(G223) );
  INV_X1 U1028 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1029 ( .A(G171), .B(G1961), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n929), .A2(G1348), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n947) );
  XNOR2_X1 U1032 ( .A(G1341), .B(n932), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(G303), .A2(G1971), .ZN(n937) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(G1956), .B(G299), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1040 ( .A(KEYINPUT123), .B(n943), .Z(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n955) );
  XOR2_X1 U1043 ( .A(G1966), .B(n948), .Z(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(n951), .B(KEYINPUT122), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n953), .B(n952), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G16), .B(KEYINPUT56), .Z(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n1008) );
  XOR2_X1 U1051 ( .A(G1966), .B(G21), .Z(n968) );
  XOR2_X1 U1052 ( .A(G1348), .B(G4), .Z(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT59), .B(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G19), .B(G1341), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G1956), .B(G20), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G1981), .B(G6), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1060 ( .A(KEYINPUT124), .B(n965), .Z(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT60), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G5), .B(G1961), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT125), .B(n971), .ZN(n979) );
  XOR2_X1 U1066 ( .A(G1986), .B(G24), .Z(n975) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(G23), .B(G1976), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(KEYINPUT126), .B(n976), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(KEYINPUT58), .B(n977), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1074 ( .A(KEYINPUT61), .B(n980), .Z(n981) );
  NOR2_X1 U1075 ( .A1(G16), .A2(n981), .ZN(n1005) );
  XOR2_X1 U1076 ( .A(G2084), .B(G34), .Z(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT54), .B(n982), .ZN(n1000) );
  XNOR2_X1 U1078 ( .A(G2090), .B(G35), .ZN(n998) );
  XNOR2_X1 U1079 ( .A(G27), .B(n983), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(KEYINPUT119), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G2067), .B(G26), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(G2072), .B(G33), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(G28), .A2(n987), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(G25), .B(G1991), .ZN(n988) );
  XNOR2_X1 U1086 ( .A(KEYINPUT118), .B(n988), .ZN(n989) );
  NOR2_X1 U1087 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(G32), .B(n993), .ZN(n994) );
  NOR2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(KEYINPUT53), .B(n996), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(n1001), .B(KEYINPUT120), .ZN(n1002) );
  XNOR2_X1 U1095 ( .A(n1002), .B(KEYINPUT55), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(G29), .A2(n1003), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(G11), .A2(n1006), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(n1009), .B(KEYINPUT127), .ZN(n1039) );
  INV_X1 U1101 ( .A(G29), .ZN(n1037) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT115), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1106 ( .A(G160), .B(G2084), .Z(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT116), .B(n1019), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(n1020), .B(KEYINPUT117), .Z(n1021) );
  XOR2_X1 U1110 ( .A(G2072), .B(n1021), .Z(n1023) );
  XOR2_X1 U1111 ( .A(G164), .B(G2078), .Z(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(KEYINPUT50), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(G2090), .B(G162), .Z(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(KEYINPUT51), .B(n1029), .Z(n1031) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1120 ( .A(KEYINPUT52), .B(n1034), .Z(n1035) );
  NOR2_X1 U1121 ( .A1(KEYINPUT55), .A2(n1035), .ZN(n1036) );
  NOR2_X1 U1122 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1123 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1040), .Z(G150) );
  INV_X1 U1125 ( .A(G150), .ZN(G311) );
endmodule

