

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579;

  XOR2_X1 U324 ( .A(G64GAT), .B(G92GAT), .Z(n292) );
  INV_X1 U325 ( .A(KEYINPUT46), .ZN(n377) );
  INV_X1 U326 ( .A(KEYINPUT31), .ZN(n371) );
  XNOR2_X1 U327 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U328 ( .A(n374), .B(n373), .ZN(n375) );
  NOR2_X1 U329 ( .A1(n525), .A2(n444), .ZN(n557) );
  XNOR2_X1 U330 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n445) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(G1348GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT68), .B(G1GAT), .Z(n294) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(G197GAT), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n307) );
  XNOR2_X1 U335 ( .A(G50GAT), .B(G22GAT), .ZN(n295) );
  XNOR2_X1 U336 ( .A(n295), .B(G141GAT), .ZN(n326) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G8GAT), .Z(n413) );
  XOR2_X1 U338 ( .A(n326), .B(n413), .Z(n297) );
  NAND2_X1 U339 ( .A1(G229GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U341 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n299) );
  XNOR2_X1 U342 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U344 ( .A(n301), .B(n300), .Z(n305) );
  XNOR2_X1 U345 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n302), .B(KEYINPUT7), .ZN(n382) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G15GAT), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n303), .B(G113GAT), .ZN(n316) );
  XNOR2_X1 U349 ( .A(n382), .B(n316), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n565) );
  XNOR2_X1 U352 ( .A(KEYINPUT69), .B(n565), .ZN(n526) );
  XOR2_X1 U353 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n309) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U356 ( .A(n310), .B(G176GAT), .Z(n314) );
  XNOR2_X1 U357 ( .A(G134GAT), .B(G127GAT), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n311), .B(KEYINPUT0), .ZN(n433) );
  XNOR2_X1 U359 ( .A(G99GAT), .B(G71GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n312), .B(G120GAT), .ZN(n362) );
  XNOR2_X1 U361 ( .A(n433), .B(n362), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n321) );
  XOR2_X1 U364 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n318) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G183GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n320) );
  XOR2_X1 U367 ( .A(G190GAT), .B(KEYINPUT17), .Z(n319) );
  XOR2_X1 U368 ( .A(n320), .B(n319), .Z(n419) );
  XOR2_X2 U369 ( .A(n321), .B(n419), .Z(n525) );
  XOR2_X1 U370 ( .A(G211GAT), .B(KEYINPUT21), .Z(n323) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G218GAT), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n418) );
  XOR2_X1 U373 ( .A(n418), .B(KEYINPUT24), .Z(n325) );
  NAND2_X1 U374 ( .A1(G228GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n339) );
  XOR2_X1 U376 ( .A(KEYINPUT23), .B(G106GAT), .Z(n328) );
  XOR2_X1 U377 ( .A(KEYINPUT74), .B(G162GAT), .Z(n394) );
  XNOR2_X1 U378 ( .A(n326), .B(n394), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U380 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n330) );
  XNOR2_X1 U381 ( .A(G204GAT), .B(KEYINPUT86), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U383 ( .A(n332), .B(n331), .Z(n337) );
  XNOR2_X1 U384 ( .A(G78GAT), .B(KEYINPUT71), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n333), .B(G148GAT), .ZN(n367) );
  XOR2_X1 U386 ( .A(G155GAT), .B(KEYINPUT3), .Z(n335) );
  XNOR2_X1 U387 ( .A(KEYINPUT87), .B(KEYINPUT2), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n432) );
  XNOR2_X1 U389 ( .A(n367), .B(n432), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n456) );
  XOR2_X1 U392 ( .A(KEYINPUT12), .B(KEYINPUT82), .Z(n341) );
  XNOR2_X1 U393 ( .A(KEYINPUT79), .B(KEYINPUT14), .ZN(n340) );
  XNOR2_X1 U394 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U395 ( .A(G57GAT), .B(KEYINPUT13), .Z(n370) );
  XOR2_X1 U396 ( .A(n370), .B(G64GAT), .Z(n343) );
  XNOR2_X1 U397 ( .A(G183GAT), .B(G127GAT), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U399 ( .A(n345), .B(n344), .Z(n347) );
  NAND2_X1 U400 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U402 ( .A(G211GAT), .B(G78GAT), .Z(n349) );
  XNOR2_X1 U403 ( .A(G15GAT), .B(G71GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U405 ( .A(n351), .B(n350), .Z(n359) );
  XOR2_X1 U406 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n353) );
  XNOR2_X1 U407 ( .A(KEYINPUT15), .B(KEYINPUT80), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U409 ( .A(G155GAT), .B(G8GAT), .Z(n355) );
  XNOR2_X1 U410 ( .A(G1GAT), .B(G22GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n359), .B(n358), .Z(n572) );
  INV_X1 U414 ( .A(n572), .ZN(n553) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(G85GAT), .ZN(n360) );
  XOR2_X1 U416 ( .A(n360), .B(KEYINPUT72), .Z(n381) );
  INV_X1 U417 ( .A(n381), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n376) );
  XOR2_X1 U419 ( .A(KEYINPUT70), .B(KEYINPUT73), .Z(n364) );
  NAND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U422 ( .A(n365), .B(KEYINPUT33), .Z(n369) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(G204GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n292), .B(n366), .ZN(n416) );
  XNOR2_X1 U425 ( .A(n367), .B(n416), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n370), .B(KEYINPUT32), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n568) );
  XOR2_X1 U429 ( .A(KEYINPUT41), .B(n568), .Z(n540) );
  OR2_X1 U430 ( .A1(n540), .A2(n565), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U432 ( .A1(n553), .A2(n379), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n380), .B(KEYINPUT114), .ZN(n403) );
  XOR2_X1 U434 ( .A(n382), .B(n381), .Z(n402) );
  XOR2_X1 U435 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n384) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(KEYINPUT9), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U438 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n386) );
  XNOR2_X1 U439 ( .A(KEYINPUT10), .B(KEYINPUT76), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U441 ( .A(n388), .B(n387), .Z(n400) );
  XOR2_X1 U442 ( .A(KEYINPUT64), .B(G92GAT), .Z(n390) );
  XNOR2_X1 U443 ( .A(G190GAT), .B(G134GAT), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n398) );
  XOR2_X1 U445 ( .A(G218GAT), .B(G99GAT), .Z(n392) );
  XNOR2_X1 U446 ( .A(G43GAT), .B(G50GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U448 ( .A(n394), .B(n393), .Z(n396) );
  NAND2_X1 U449 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U453 ( .A(n402), .B(n401), .Z(n558) );
  INV_X1 U454 ( .A(n558), .ZN(n546) );
  NAND2_X1 U455 ( .A1(n403), .A2(n546), .ZN(n404) );
  XNOR2_X1 U456 ( .A(n404), .B(KEYINPUT47), .ZN(n411) );
  XOR2_X1 U457 ( .A(KEYINPUT45), .B(KEYINPUT65), .Z(n406) );
  XOR2_X1 U458 ( .A(KEYINPUT36), .B(n546), .Z(n575) );
  NAND2_X1 U459 ( .A1(n553), .A2(n575), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U461 ( .A(KEYINPUT115), .B(n407), .ZN(n408) );
  NAND2_X1 U462 ( .A1(n408), .A2(n568), .ZN(n409) );
  NOR2_X1 U463 ( .A1(n409), .A2(n526), .ZN(n410) );
  NOR2_X1 U464 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U465 ( .A(KEYINPUT48), .B(n412), .ZN(n521) );
  XOR2_X1 U466 ( .A(KEYINPUT90), .B(n413), .Z(n415) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U469 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U470 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U471 ( .A(n421), .B(n420), .Z(n510) );
  XOR2_X1 U472 ( .A(n510), .B(KEYINPUT119), .Z(n422) );
  NOR2_X1 U473 ( .A1(n521), .A2(n422), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n423), .B(KEYINPUT54), .ZN(n442) );
  XOR2_X1 U475 ( .A(KEYINPUT1), .B(G57GAT), .Z(n425) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(G141GAT), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n441) );
  XOR2_X1 U478 ( .A(G85GAT), .B(G148GAT), .Z(n427) );
  XNOR2_X1 U479 ( .A(G113GAT), .B(G120GAT), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U481 ( .A(G29GAT), .B(G162GAT), .Z(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n437) );
  XNOR2_X1 U483 ( .A(KEYINPUT89), .B(KEYINPUT5), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n430), .B(KEYINPUT4), .ZN(n431) );
  XOR2_X1 U485 ( .A(n431), .B(KEYINPUT6), .Z(n435) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n437), .B(n436), .ZN(n439) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n507) );
  NAND2_X1 U492 ( .A1(n442), .A2(n507), .ZN(n563) );
  NOR2_X1 U493 ( .A1(n456), .A2(n563), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n443), .B(KEYINPUT55), .ZN(n444) );
  NAND2_X1 U495 ( .A1(n526), .A2(n557), .ZN(n446) );
  NOR2_X1 U496 ( .A1(n558), .A2(n572), .ZN(n447) );
  XNOR2_X1 U497 ( .A(KEYINPUT16), .B(n447), .ZN(n465) );
  XOR2_X1 U498 ( .A(n510), .B(KEYINPUT91), .Z(n448) );
  XNOR2_X1 U499 ( .A(n448), .B(KEYINPUT27), .ZN(n458) );
  NOR2_X1 U500 ( .A1(n458), .A2(n507), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT92), .B(n449), .Z(n520) );
  XNOR2_X1 U502 ( .A(KEYINPUT85), .B(n525), .ZN(n450) );
  NOR2_X1 U503 ( .A1(n520), .A2(n450), .ZN(n451) );
  XOR2_X1 U504 ( .A(n456), .B(KEYINPUT28), .Z(n523) );
  NAND2_X1 U505 ( .A1(n451), .A2(n523), .ZN(n464) );
  OR2_X1 U506 ( .A1(n525), .A2(n510), .ZN(n452) );
  XNOR2_X1 U507 ( .A(KEYINPUT93), .B(n452), .ZN(n453) );
  NOR2_X1 U508 ( .A1(n456), .A2(n453), .ZN(n454) );
  XOR2_X1 U509 ( .A(KEYINPUT94), .B(n454), .Z(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(n455), .ZN(n460) );
  NAND2_X1 U511 ( .A1(n525), .A2(n456), .ZN(n457) );
  XOR2_X1 U512 ( .A(n457), .B(KEYINPUT26), .Z(n538) );
  INV_X1 U513 ( .A(n538), .ZN(n564) );
  NOR2_X1 U514 ( .A1(n564), .A2(n458), .ZN(n459) );
  NOR2_X1 U515 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT95), .B(n461), .ZN(n462) );
  NAND2_X1 U517 ( .A1(n462), .A2(n507), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n464), .A2(n463), .ZN(n475) );
  NAND2_X1 U519 ( .A1(n465), .A2(n475), .ZN(n466) );
  XOR2_X1 U520 ( .A(n466), .B(KEYINPUT96), .Z(n494) );
  AND2_X1 U521 ( .A1(n526), .A2(n568), .ZN(n479) );
  NAND2_X1 U522 ( .A1(n494), .A2(n479), .ZN(n473) );
  NOR2_X1 U523 ( .A1(n507), .A2(n473), .ZN(n467) );
  XOR2_X1 U524 ( .A(n467), .B(KEYINPUT34), .Z(n468) );
  XNOR2_X1 U525 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NOR2_X1 U526 ( .A1(n510), .A2(n473), .ZN(n470) );
  XNOR2_X1 U527 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(G1325GAT) );
  NOR2_X1 U529 ( .A1(n525), .A2(n473), .ZN(n472) );
  XNOR2_X1 U530 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n472), .B(n471), .ZN(G1326GAT) );
  NOR2_X1 U532 ( .A1(n523), .A2(n473), .ZN(n474) );
  XOR2_X1 U533 ( .A(G22GAT), .B(n474), .Z(G1327GAT) );
  NAND2_X1 U534 ( .A1(n575), .A2(n475), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n553), .A2(n476), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT37), .B(KEYINPUT98), .ZN(n477) );
  XOR2_X1 U537 ( .A(n478), .B(n477), .Z(n505) );
  NAND2_X1 U538 ( .A1(n505), .A2(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(KEYINPUT38), .B(n480), .ZN(n489) );
  NOR2_X1 U540 ( .A1(n489), .A2(n507), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT39), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G29GAT), .B(n482), .ZN(G1328GAT) );
  NOR2_X1 U543 ( .A1(n489), .A2(n510), .ZN(n484) );
  XNOR2_X1 U544 ( .A(G36GAT), .B(KEYINPUT99), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(G1329GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n486) );
  XNOR2_X1 U547 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n488) );
  NOR2_X1 U549 ( .A1(n489), .A2(n525), .ZN(n487) );
  XOR2_X1 U550 ( .A(n488), .B(n487), .Z(G1330GAT) );
  XNOR2_X1 U551 ( .A(KEYINPUT103), .B(KEYINPUT102), .ZN(n491) );
  NOR2_X1 U552 ( .A1(n523), .A2(n489), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G50GAT), .B(n492), .ZN(G1331GAT) );
  XOR2_X1 U555 ( .A(n540), .B(KEYINPUT104), .Z(n548) );
  NAND2_X1 U556 ( .A1(n565), .A2(n548), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(KEYINPUT105), .ZN(n506) );
  NAND2_X1 U558 ( .A1(n506), .A2(n494), .ZN(n501) );
  NOR2_X1 U559 ( .A1(n507), .A2(n501), .ZN(n496) );
  XNOR2_X1 U560 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n495) );
  XNOR2_X1 U561 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n497), .Z(G1332GAT) );
  NOR2_X1 U563 ( .A1(n510), .A2(n501), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(G1333GAT) );
  NOR2_X1 U566 ( .A1(n525), .A2(n501), .ZN(n500) );
  XOR2_X1 U567 ( .A(G71GAT), .B(n500), .Z(G1334GAT) );
  NOR2_X1 U568 ( .A1(n523), .A2(n501), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(n504), .ZN(G1335GAT) );
  NAND2_X1 U572 ( .A1(n506), .A2(n505), .ZN(n516) );
  NOR2_X1 U573 ( .A1(n507), .A2(n516), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n516), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n516), .ZN(n514) );
  XOR2_X1 U581 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n515), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n523), .A2(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT116), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n523), .A2(n537), .ZN(n524) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n534), .A2(n526), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT117), .B(n527), .Z(n528) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U595 ( .A1(n534), .A2(n548), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n532) );
  NAND2_X1 U598 ( .A1(n534), .A2(n553), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n533), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U602 ( .A1(n534), .A2(n558), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n565), .A2(n545), .ZN(n539) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n539), .Z(G1344GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n545), .ZN(n542) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n572), .A2(n545), .ZN(n544) );
  XOR2_X1 U612 ( .A(G155GAT), .B(n544), .Z(G1346GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(G162GAT), .B(n547), .Z(G1347GAT) );
  XOR2_X1 U615 ( .A(G176GAT), .B(KEYINPUT57), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n557), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1349GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n555) );
  NAND2_X1 U621 ( .A1(n557), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G183GAT), .B(n556), .ZN(G1350GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n560), .ZN(G1351GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n562) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n567) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n576) );
  INV_X1 U631 ( .A(n576), .ZN(n571) );
  NOR2_X1 U632 ( .A1(n565), .A2(n571), .ZN(n566) );
  XOR2_X1 U633 ( .A(n567), .B(n566), .Z(G1352GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n571), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n578) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(G218GAT), .B(n579), .Z(G1355GAT) );
endmodule

