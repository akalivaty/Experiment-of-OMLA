//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(KEYINPUT67), .A3(new_n196), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT0), .A4(G128), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT0), .B(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n200), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n203), .A2(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n201), .A2(G143), .ZN(new_n215));
  OAI211_X1 g029(.A(G128), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n202), .B(new_n204), .C1(KEYINPUT1), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n188), .A2(G137), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n190), .A2(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n196), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n223), .A3(KEYINPUT69), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n218), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n196), .A2(new_n222), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n224), .A2(KEYINPUT30), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n199), .A2(KEYINPUT68), .A3(new_n200), .A4(new_n209), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n212), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT2), .A2(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT2), .A3(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G119), .ZN(new_n243));
  INV_X1    g057(.A(G119), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT66), .A3(G116), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(G119), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n245), .A2(new_n246), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(new_n239), .A3(new_n236), .A4(new_n243), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n209), .A2(new_n197), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n219), .B1(new_n223), .B2(KEYINPUT64), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n196), .A2(new_n222), .A3(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n231), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n224), .A2(new_n251), .A3(new_n228), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n212), .A2(new_n259), .A3(new_n230), .ZN(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT31), .B1(new_n258), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n266), .B(KEYINPUT71), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n248), .A2(new_n250), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n255), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n260), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n219), .B2(new_n223), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT28), .B1(new_n276), .B2(new_n210), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n271), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n260), .A2(new_n266), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT31), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n231), .A2(new_n257), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n260), .A3(new_n266), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n270), .A2(new_n278), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n278), .A2(new_n282), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n269), .B(new_n280), .C1(new_n279), .C2(new_n281), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT70), .B1(new_n283), .B2(KEYINPUT31), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n286), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n288), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n290), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n281), .A2(new_n260), .ZN(new_n299));
  INV_X1    g113(.A(new_n266), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n271), .A2(new_n277), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n304), .B2(new_n275), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n260), .A2(new_n274), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT72), .B(new_n303), .C1(new_n306), .C2(new_n272), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n301), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n277), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n212), .A2(new_n230), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n224), .A2(new_n228), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n212), .A2(new_n230), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n311), .A2(new_n259), .B1(new_n313), .B2(new_n273), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n310), .B1(new_n314), .B2(new_n272), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G472), .B1(new_n308), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n296), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n289), .A2(new_n298), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT9), .B(G234), .ZN(new_n321));
  OAI21_X1  g135(.A(G221), .B1(new_n321), .B2(G902), .ZN(new_n322));
  OAI21_X1  g136(.A(G214), .B1(G237), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G210), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G122), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT8), .ZN(new_n328));
  INV_X1    g142(.A(G104), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT3), .B1(new_n329), .B2(G107), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n331));
  INV_X1    g145(.A(G107), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G104), .ZN(new_n333));
  INV_X1    g147(.A(G101), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(G107), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n329), .A2(G107), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n332), .A2(G104), .ZN(new_n338));
  OAI21_X1  g152(.A(G101), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT5), .A4(new_n246), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n242), .A2(G119), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT5), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n238), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AND4_X1   g158(.A1(new_n250), .A2(new_n336), .A3(new_n339), .A4(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n250), .A2(new_n344), .B1(new_n336), .B2(new_n339), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n328), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n348));
  INV_X1    g162(.A(G125), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n213), .A2(G128), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(new_n206), .ZN(new_n351));
  INV_X1    g165(.A(new_n218), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n348), .B(new_n349), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n208), .A2(G125), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G125), .B1(new_n216), .B2(new_n218), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n348), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n262), .A2(G224), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT85), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT7), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n355), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n356), .A2(new_n348), .B1(G125), .B2(new_n208), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n226), .A2(new_n349), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT83), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n347), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n327), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n330), .A2(new_n333), .A3(new_n335), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT77), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n330), .A2(new_n333), .A3(new_n371), .A4(new_n335), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n334), .A2(KEYINPUT4), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n370), .A2(KEYINPUT78), .A3(new_n372), .A4(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n370), .A2(G101), .A3(new_n372), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n336), .A2(KEYINPUT4), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n379), .A2(new_n380), .B1(new_n250), .B2(new_n248), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n345), .B(new_n368), .C1(new_n378), .C2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n309), .B1(new_n367), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT86), .B(new_n309), .C1(new_n367), .C2(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n363), .A2(new_n365), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n359), .B(KEYINPUT84), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n345), .B1(new_n378), .B2(new_n381), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n327), .A2(KEYINPUT82), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n382), .A2(new_n391), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n392), .A2(new_n391), .A3(new_n394), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n326), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n390), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n392), .A2(new_n327), .ZN(new_n401));
  INV_X1    g215(.A(new_n392), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n401), .A2(KEYINPUT6), .B1(new_n402), .B2(new_n393), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n400), .B1(new_n403), .B2(new_n396), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(new_n325), .A3(new_n386), .A4(new_n385), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n324), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G469), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n194), .A2(KEYINPUT67), .A3(new_n196), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT67), .B1(new_n194), .B2(new_n196), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n336), .A2(new_n339), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n226), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n216), .A2(new_n336), .A3(new_n339), .A4(new_n218), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI211_X1 g228(.A(KEYINPUT79), .B(KEYINPUT12), .C1(new_n410), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n200), .A3(new_n199), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT12), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n414), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n197), .A2(KEYINPUT12), .ZN(new_n421));
  OAI22_X1  g235(.A1(new_n415), .A2(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G140), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n262), .A2(G227), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n208), .B1(new_n379), .B2(new_n380), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n378), .A2(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n410), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n378), .A2(new_n426), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n428), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n433), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g250(.A(KEYINPUT81), .B(new_n425), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n434), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n410), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n429), .A2(new_n430), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT81), .B1(new_n442), .B2(new_n425), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n407), .B(new_n309), .C1(new_n438), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(G469), .A2(G902), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n436), .B1(new_n431), .B2(KEYINPUT80), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n435), .B2(new_n425), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n425), .B(KEYINPUT76), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n420), .A2(new_n421), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n417), .A2(new_n418), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT79), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n417), .A2(new_n416), .A3(new_n418), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n455), .B2(new_n435), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n456), .A3(G469), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n444), .A2(new_n445), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G217), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n321), .A2(new_n459), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G128), .B(G143), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT95), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n188), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(KEYINPUT13), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n203), .A2(G128), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(G134), .C1(KEYINPUT13), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G122), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G116), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n242), .A2(G122), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(G107), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n464), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n332), .B1(new_n469), .B2(KEYINPUT14), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n471), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT95), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n462), .B(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G134), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n464), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n461), .B1(new_n473), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n475), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n477), .A2(G134), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n463), .A2(new_n188), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n464), .A2(new_n467), .A3(new_n472), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n460), .ZN(new_n486));
  AOI21_X1  g300(.A(G902), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n487), .B(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(G237), .A2(G953), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n203), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(G143), .A3(G214), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(KEYINPUT88), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT18), .A3(G131), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT18), .A2(G131), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n493), .A2(KEYINPUT88), .A3(new_n497), .A4(new_n494), .ZN(new_n498));
  INV_X1    g312(.A(G140), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G125), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n349), .A2(G140), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G146), .ZN(new_n503));
  XNOR2_X1  g317(.A(G125), .B(G140), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n201), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n503), .B2(new_n505), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n496), .B(new_n498), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(G113), .B(G122), .Z(new_n510));
  XOR2_X1   g324(.A(KEYINPUT90), .B(G104), .Z(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT16), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n349), .A2(KEYINPUT16), .A3(G140), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(G146), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G146), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  OAI21_X1  g331(.A(KEYINPUT92), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n515), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n491), .A2(G143), .A3(G214), .ZN(new_n523));
  AOI21_X1  g337(.A(G143), .B1(new_n491), .B2(G214), .ZN(new_n524));
  OAI21_X1  g338(.A(G131), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n518), .B(new_n521), .C1(new_n522), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n493), .A2(new_n195), .A3(new_n494), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n529), .B2(KEYINPUT17), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT93), .A4(new_n522), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n509), .B(new_n512), .C1(new_n526), .C2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n525), .A2(new_n522), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n516), .A2(new_n517), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n520), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n537), .A2(new_n518), .A3(new_n530), .A4(new_n531), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n512), .B1(new_n538), .B2(new_n509), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n309), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT94), .B(G475), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT19), .B1(new_n504), .B2(KEYINPUT89), .ZN(new_n543));
  AND4_X1   g357(.A1(KEYINPUT89), .A2(new_n500), .A3(new_n501), .A4(KEYINPUT19), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n529), .B(new_n515), .C1(new_n545), .C2(G146), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n509), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n512), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT91), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n550), .B(new_n512), .C1(new_n509), .C2(new_n546), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n533), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n490), .B(new_n542), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n262), .A2(G952), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(G234), .B2(G237), .ZN(new_n559));
  NAND2_X1  g373(.A1(G234), .A2(G237), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(G902), .A3(G953), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n561), .B(KEYINPUT96), .Z(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT21), .B(G898), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n559), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  AND4_X1   g380(.A1(new_n322), .A2(new_n406), .A3(new_n458), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n459), .B1(G234), .B2(new_n309), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n217), .A2(G119), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n244), .A2(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT74), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT74), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT24), .B(G110), .Z(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT75), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n572), .A2(new_n578), .A3(new_n574), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n581));
  INV_X1    g395(.A(new_n569), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n570), .B(new_n581), .C1(new_n582), .C2(KEYINPUT23), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n519), .A2(new_n515), .B1(G110), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n583), .A2(G110), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n575), .B1(new_n572), .B2(new_n574), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n515), .B(new_n505), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT22), .B(G137), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n585), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n585), .B2(new_n588), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT25), .B1(new_n595), .B2(new_n309), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n588), .ZN(new_n597));
  INV_X1    g411(.A(new_n591), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n309), .A3(new_n592), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT25), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n568), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n568), .A2(G902), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n320), .A2(new_n567), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  INV_X1    g423(.A(new_n565), .ZN(new_n610));
  INV_X1    g424(.A(new_n541), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n509), .B1(new_n526), .B2(new_n532), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n548), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n533), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(new_n309), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n552), .A2(new_n554), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT20), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n480), .A2(new_n486), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n480), .A2(new_n486), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(G478), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n488), .A2(new_n309), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n487), .B2(new_n488), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n406), .A2(new_n610), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n285), .A2(new_n309), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n292), .A2(new_n293), .ZN(new_n634));
  INV_X1    g448(.A(new_n291), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n295), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n285), .B2(new_n309), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n638), .B2(KEYINPUT97), .ZN(new_n639));
  INV_X1    g453(.A(new_n322), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n422), .A2(new_n441), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n641), .A2(new_n450), .B1(new_n446), .B2(new_n448), .ZN(new_n642));
  OAI21_X1  g456(.A(G469), .B1(new_n642), .B2(G902), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n640), .B(new_n606), .C1(new_n643), .C2(new_n444), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n629), .A2(new_n633), .A3(new_n639), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  NAND2_X1  g461(.A1(new_n399), .A2(new_n405), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n323), .ZN(new_n649));
  INV_X1    g463(.A(new_n489), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n487), .B(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(new_n542), .C1(new_n555), .C2(new_n556), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n649), .A2(new_n565), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n653), .A2(new_n633), .A3(new_n639), .A4(new_n644), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT98), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  NAND2_X1  g471(.A1(new_n458), .A2(new_n322), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n649), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n598), .A2(KEYINPUT36), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n597), .B(new_n661), .Z(new_n662));
  INV_X1    g476(.A(new_n604), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n603), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n568), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n595), .A2(KEYINPUT25), .A3(new_n309), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n600), .A2(new_n601), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n662), .A2(new_n663), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT99), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n672), .A2(new_n565), .A3(new_n557), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n659), .A2(new_n633), .A3(new_n639), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  AND2_X1   g490(.A1(new_n320), .A2(new_n659), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n665), .A2(new_n671), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n559), .B(KEYINPUT100), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(G900), .B2(new_n562), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n679), .B1(new_n652), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n619), .A2(KEYINPUT101), .A3(new_n651), .A4(new_n681), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n678), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  XOR2_X1   g501(.A(new_n648), .B(KEYINPUT38), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n617), .A2(new_n618), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n490), .B1(new_n689), .B2(new_n542), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  OR3_X1    g505(.A1(new_n688), .A2(new_n324), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n640), .B1(new_n643), .B2(new_n444), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n681), .B(KEYINPUT39), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n603), .A2(new_n664), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n313), .A2(new_n273), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n260), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n699), .A2(new_n271), .B1(new_n279), .B2(new_n281), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n289), .A2(new_n298), .A3(new_n319), .A4(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n692), .A2(new_n696), .A3(new_n697), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n203), .ZN(G45));
  OR2_X1    g519(.A1(new_n619), .A2(new_n627), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n706), .A2(new_n672), .A3(new_n682), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n677), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  AND3_X1   g523(.A1(new_n285), .A2(KEYINPUT73), .A3(new_n296), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT73), .B1(new_n285), .B2(new_n296), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n277), .B1(new_n699), .B2(KEYINPUT28), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n301), .A2(new_n305), .A3(new_n307), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n637), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n287), .B2(new_n288), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n606), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n309), .B1(new_n438), .B2(new_n443), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n322), .A3(new_n444), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n724), .A3(new_n322), .A4(new_n444), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n719), .A2(new_n629), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND3_X1  g543(.A1(new_n719), .A2(new_n653), .A3(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NAND4_X1  g545(.A1(new_n678), .A2(new_n610), .A3(new_n490), .A4(new_n619), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n718), .B2(new_n712), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n723), .A2(new_n406), .A3(new_n725), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  XNOR2_X1  g550(.A(KEYINPUT104), .B(G472), .ZN(new_n737));
  INV_X1    g551(.A(new_n271), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n268), .B1(new_n713), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n315), .A2(new_n271), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n268), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n743), .A3(new_n282), .ZN(new_n744));
  AOI221_X4 g558(.A(new_n606), .B1(new_n630), .B2(new_n737), .C1(new_n744), .C2(new_n286), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n649), .A2(new_n691), .A3(new_n565), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n726), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR2_X1   g562(.A1(new_n706), .A2(new_n682), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n723), .A2(new_n749), .A3(new_n406), .A4(new_n725), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n744), .A2(new_n286), .B1(new_n630), .B2(new_n737), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n697), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n349), .ZN(G27));
  NAND3_X1  g568(.A1(new_n399), .A2(new_n323), .A3(new_n405), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AND4_X1   g570(.A1(KEYINPUT42), .A2(new_n749), .A3(new_n693), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n285), .A2(new_n296), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n318), .B(new_n758), .C1(new_n636), .C2(KEYINPUT32), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n759), .A2(KEYINPUT105), .A3(new_n607), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT105), .B1(new_n759), .B2(new_n607), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n658), .A2(new_n755), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n320), .A2(new_n607), .A3(new_n763), .A4(new_n749), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  AND2_X1   g582(.A1(new_n683), .A2(new_n684), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n320), .A2(new_n607), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NAND2_X1  g585(.A1(new_n449), .A2(new_n456), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n407), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n642), .A2(KEYINPUT45), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n445), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n445), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n444), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n322), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n689), .A2(new_n542), .A3(new_n624), .A4(new_n626), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(new_n697), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n633), .A2(new_n639), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(KEYINPUT44), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT44), .B1(new_n790), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n755), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n786), .A2(new_n694), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n785), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n322), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n749), .A2(new_n606), .A3(new_n756), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n800), .A2(new_n320), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  NAND2_X1  g617(.A1(new_n721), .A2(new_n444), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT107), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT49), .Z(new_n806));
  NOR3_X1   g620(.A1(new_n787), .A2(new_n640), .A3(new_n324), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n688), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n607), .A3(new_n703), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n558), .B(KEYINPUT116), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n788), .A2(new_n680), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n745), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n813), .B2(new_n734), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n726), .A2(new_n756), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n760), .A2(new_n761), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n811), .ZN(new_n818));
  NAND2_X1  g632(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n703), .A2(new_n607), .A3(new_n559), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(KEYINPUT115), .A3(new_n821), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n824), .A2(new_n628), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n827));
  AOI211_X1 g641(.A(new_n820), .B(new_n826), .C1(new_n818), .C2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n798), .B(new_n799), .C1(new_n322), .C2(new_n805), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n756), .A3(new_n813), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n697), .A2(new_n816), .A3(new_n751), .A4(new_n811), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n726), .A2(new_n324), .A3(new_n688), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(new_n812), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT50), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n824), .A2(new_n619), .A3(new_n627), .A4(new_n825), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n830), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT51), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT51), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n828), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n746), .A2(new_n725), .A3(new_n723), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n842), .A2(new_n745), .B1(new_n733), .B2(new_n734), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n751), .A2(new_n763), .A3(new_n697), .A4(new_n749), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n672), .A2(new_n557), .A3(new_n682), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n320), .A2(new_n763), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n770), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n719), .B(new_n726), .C1(new_n629), .C2(new_n653), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n767), .A2(new_n843), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n608), .A2(new_n645), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT108), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n654), .A2(new_n674), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT108), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n608), .A2(new_n645), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT109), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n608), .A2(new_n854), .A3(new_n645), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n854), .B1(new_n608), .B2(new_n645), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n858), .A2(new_n859), .A3(new_n852), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT109), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n848), .A2(new_n735), .A3(new_n747), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n770), .A2(new_n844), .A3(new_n846), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n762), .B2(new_n766), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n320), .B(new_n659), .C1(new_n685), .C2(new_n707), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n406), .A2(new_n690), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n658), .A2(new_n682), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n702), .A2(new_n789), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n867), .B1(new_n873), .B2(new_n753), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n734), .A2(new_n697), .A3(new_n749), .A4(new_n751), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n868), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n866), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(KEYINPUT110), .A3(new_n876), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT110), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n883), .B(new_n867), .C1(new_n873), .C2(new_n753), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n849), .A2(new_n879), .A3(new_n856), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT112), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n882), .A2(new_n884), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n862), .A4(new_n864), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT112), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n880), .A2(new_n881), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n866), .A2(new_n879), .A3(new_n885), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n857), .A2(new_n865), .B1(new_n874), .B2(new_n876), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n894), .B(KEYINPUT54), .C1(new_n879), .C2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(KEYINPUT111), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n878), .A2(KEYINPUT53), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT111), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT54), .A4(new_n894), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n841), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n809), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n262), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n309), .B1(new_n880), .B2(new_n892), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT56), .B1(new_n906), .B2(G210), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n403), .A2(new_n396), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n390), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n404), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n905), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n907), .B2(new_n913), .ZN(G51));
  OR2_X1    g729(.A1(new_n438), .A2(new_n443), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT112), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n917), .A2(new_n918), .B1(new_n895), .B2(KEYINPUT53), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT54), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n920), .A2(new_n893), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n445), .B(KEYINPUT57), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  INV_X1    g738(.A(new_n779), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n906), .B2(new_n925), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n878), .A2(new_n879), .B1(new_n888), .B2(new_n891), .ZN(new_n927));
  NOR4_X1   g741(.A1(new_n927), .A2(KEYINPUT119), .A3(new_n309), .A4(new_n779), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n904), .B1(new_n923), .B2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  INV_X1    g745(.A(new_n552), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n904), .ZN(G60));
  AND2_X1   g749(.A1(new_n621), .A2(new_n623), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n625), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n920), .B2(new_n893), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n897), .A2(new_n900), .A3(new_n939), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n904), .B(new_n941), .C1(new_n942), .C2(new_n936), .ZN(G63));
  INV_X1    g757(.A(new_n595), .ZN(new_n944));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n927), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n946), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n662), .B(KEYINPUT121), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n919), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n905), .A3(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(KEYINPUT122), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n919), .A2(new_n948), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n904), .B1(new_n956), .B2(new_n944), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(KEYINPUT122), .A3(new_n952), .A4(new_n950), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n955), .A2(new_n958), .ZN(G66));
  INV_X1    g773(.A(G224), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n564), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n860), .A2(new_n862), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n963), .B2(G953), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n908), .B1(G898), .B2(new_n262), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT123), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G69));
  AOI21_X1  g781(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AOI22_X1  g783(.A1(new_n311), .A2(new_n229), .B1(new_n256), .B2(new_n255), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(new_n545), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n875), .A2(new_n868), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n704), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT62), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n976));
  AOI211_X1 g790(.A(new_n755), .B(new_n695), .C1(new_n706), .C2(new_n652), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n719), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT125), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n795), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n976), .B1(new_n795), .B2(new_n979), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n802), .B(new_n975), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n972), .B1(new_n982), .B2(new_n262), .ZN(new_n983));
  INV_X1    g797(.A(new_n973), .ZN(new_n984));
  AND4_X1   g798(.A1(new_n767), .A2(new_n795), .A3(new_n770), .A4(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n786), .A2(new_n694), .A3(new_n817), .A4(new_n870), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n802), .A2(new_n262), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(G900), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n972), .B1(new_n988), .B2(new_n262), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(KEYINPUT127), .B(new_n969), .C1(new_n983), .C2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n969), .A2(KEYINPUT127), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n987), .B2(new_n990), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n982), .A2(new_n262), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n993), .B(new_n995), .C1(new_n996), .C2(new_n972), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n992), .A2(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n982), .B2(new_n962), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n300), .B1(new_n281), .B2(new_n260), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n802), .A2(new_n986), .A3(new_n985), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1000), .B1(new_n1004), .B2(new_n962), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n299), .A2(new_n266), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n898), .A2(new_n894), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1000), .ZN(new_n1009));
  NOR4_X1   g823(.A1(new_n1008), .A2(new_n1006), .A3(new_n1009), .A4(new_n1002), .ZN(new_n1010));
  NOR4_X1   g824(.A1(new_n1003), .A2(new_n1007), .A3(new_n1010), .A4(new_n904), .ZN(G57));
endmodule


