//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  OR3_X1    g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT92), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT92), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n210), .B(new_n211), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT91), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT15), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n216), .A2(new_n217), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(G43gat), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT93), .B(G43gat), .Z(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G50gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n221), .B1(new_n228), .B2(new_n215), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  AOI21_X1  g031(.A(G1gat), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(KEYINPUT94), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n233), .B(new_n234), .Z(new_n235));
  XOR2_X1   g034(.A(KEYINPUT95), .B(G8gat), .Z(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT95), .A2(G8gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n229), .A2(KEYINPUT17), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n230), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n239), .A2(new_n229), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n207), .B1(new_n246), .B2(KEYINPUT96), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT18), .A4(new_n243), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n239), .B(new_n229), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n243), .B(KEYINPUT13), .Z(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n247), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(G176gat), .B(G204gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT98), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT7), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(G85gat), .A3(G92gat), .A4(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G85gat), .ZN(new_n264));
  INV_X1    g063(.A(G92gat), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n259), .B(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267));
  AOI22_X1  g066(.A1(KEYINPUT8), .A2(new_n267), .B1(new_n264), .B2(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G99gat), .B(G106gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT99), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n273), .A2(KEYINPUT99), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G71gat), .B(G78gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT97), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G57gat), .B(G64gat), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n277), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(KEYINPUT10), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n271), .ZN(new_n287));
  INV_X1    g086(.A(new_n285), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n275), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(new_n289), .B2(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n291), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n258), .B1(new_n296), .B2(KEYINPUT102), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT102), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n298), .A3(new_n257), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n254), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G134gat), .B(G162gat), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT101), .Z(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n275), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(new_n229), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT100), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n230), .A2(new_n240), .A3(new_n307), .ZN(new_n311));
  XNOR2_X1  g110(.A(G190gat), .B(G218gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(new_n310), .B2(new_n311), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n305), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(new_n311), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n312), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT101), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(new_n320), .A3(new_n314), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n285), .A2(KEYINPUT21), .ZN(new_n324));
  XNOR2_X1  g123(.A(G127gat), .B(G155gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(G211gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n326), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT21), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n239), .B1(new_n332), .B2(new_n288), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n331), .B(new_n335), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n323), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  AND2_X1   g141(.A1(G211gat), .A2(G218gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(KEYINPUT22), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n348), .B(KEYINPUT71), .Z(new_n349));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  INV_X1    g152(.A(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT65), .ZN(new_n357));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n357), .A2(new_n363), .A3(KEYINPUT25), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n356), .A2(KEYINPUT65), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n353), .A2(KEYINPUT64), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n367), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n366), .A2(new_n368), .A3(new_n352), .A4(new_n355), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n364), .A2(new_n365), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT27), .B(G183gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n354), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT28), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n376), .A3(new_n354), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT66), .B(KEYINPUT26), .ZN(new_n380));
  INV_X1    g179(.A(new_n358), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT66), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(KEYINPUT26), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT26), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT66), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT67), .B(new_n358), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n362), .B1(new_n358), .B2(new_n385), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n382), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n350), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n378), .B1(new_n391), .B2(KEYINPUT68), .ZN(new_n392));
  INV_X1    g191(.A(new_n350), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n358), .B1(new_n384), .B2(new_n386), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n388), .B1(new_n394), .B2(new_n379), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n395), .B2(new_n387), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT68), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n372), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n347), .B(new_n349), .C1(new_n399), .C2(KEYINPUT29), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n364), .A2(new_n365), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n370), .A2(new_n371), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n378), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n396), .B2(new_n397), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n390), .A2(new_n397), .A3(new_n350), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(G226gat), .A3(G233gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n397), .B1(new_n390), .B2(new_n350), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n406), .A2(new_n411), .A3(new_n378), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n412), .B2(new_n372), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n347), .B1(new_n413), .B2(new_n349), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n346), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n416));
  INV_X1    g215(.A(new_n349), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n413), .A2(new_n348), .B1(new_n407), .B2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n344), .B(new_n345), .Z(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n416), .B1(new_n415), .B2(new_n420), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n341), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n341), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n415), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT30), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n415), .A2(new_n427), .A3(new_n420), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(new_n264), .ZN(new_n431));
  XNOR2_X1  g230(.A(KEYINPUT0), .B(G57gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G120gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G113gat), .ZN(new_n436));
  INV_X1    g235(.A(G113gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G120gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n440));
  INV_X1    g239(.A(G134gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G127gat), .ZN(new_n442));
  INV_X1    g241(.A(G127gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(G134gat), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n439), .A2(new_n440), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n444), .ZN(new_n446));
  XNOR2_X1  g245(.A(G113gat), .B(G120gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G141gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(G148gat), .ZN(new_n452));
  INV_X1    g251(.A(G148gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G141gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(G155gat), .A2(G162gat), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n452), .A2(new_n454), .B1(KEYINPUT2), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT74), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n459));
  INV_X1    g258(.A(G155gat), .ZN(new_n460));
  INV_X1    g259(.A(G162gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT75), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT75), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n458), .A2(new_n462), .A3(new_n465), .A4(new_n459), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n456), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n455), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n462), .A2(KEYINPUT76), .A3(new_n455), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n470), .A2(new_n456), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n450), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT3), .B1(new_n467), .B2(new_n472), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT77), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n467), .C2(new_n472), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT4), .B1(new_n473), .B2(new_n450), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT4), .ZN(new_n483));
  NOR4_X1   g282(.A1(new_n467), .A2(new_n472), .A3(new_n449), .A4(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G225gat), .A2(G233gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n481), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n488));
  INV_X1    g287(.A(new_n486), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n450), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n467), .A2(new_n472), .A3(new_n449), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT5), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n493), .B1(new_n487), .B2(new_n488), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n434), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n487), .A2(new_n488), .ZN(new_n498));
  INV_X1    g297(.A(new_n493), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n494), .A3(new_n433), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n500), .A2(KEYINPUT6), .A3(new_n494), .A4(new_n433), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n423), .A2(new_n429), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G78gat), .B(G106gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G50gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n467), .A2(new_n472), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n410), .A3(new_n419), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n515), .A2(G228gat), .A3(G233gat), .A4(new_n477), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n410), .B1(new_n514), .B2(new_n474), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n419), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT29), .B1(new_n473), .B2(new_n475), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT84), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G228gat), .A2(G233gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT83), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n517), .A2(new_n346), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n473), .A2(new_n346), .A3(KEYINPUT29), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n473), .A2(new_n475), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(G22gat), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n477), .A2(G228gat), .A3(G233gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n521), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n346), .B1(new_n520), .B2(KEYINPUT84), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n515), .B1(new_n473), .B2(new_n475), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n419), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n524), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G22gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n531), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n513), .B1(new_n542), .B2(KEYINPUT82), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT82), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n544), .B(new_n512), .C1(new_n531), .C2(new_n541), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n510), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n522), .A2(new_n530), .A3(G22gat), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n540), .B1(new_n536), .B2(new_n539), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT82), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n512), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n542), .A2(KEYINPUT82), .A3(new_n513), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n509), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n407), .A2(new_n449), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n399), .A2(new_n450), .ZN(new_n554));
  AND2_X1   g353(.A1(G227gat), .A2(G233gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT34), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(KEYINPUT34), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G43gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G99gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  AOI21_X1  g363(.A(new_n556), .B1(new_n553), .B2(new_n554), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(KEYINPUT33), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n566), .A2(new_n568), .ZN(new_n571));
  OAI211_X1 g370(.A(KEYINPUT69), .B(new_n561), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n566), .A2(new_n568), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n559), .B2(new_n560), .ZN(new_n575));
  INV_X1    g374(.A(new_n560), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(KEYINPUT69), .A3(new_n558), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n573), .A2(new_n575), .A3(new_n577), .A4(new_n569), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n546), .A2(new_n552), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n423), .A2(new_n429), .A3(new_n505), .A4(KEYINPUT80), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n508), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n581), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT90), .B1(new_n581), .B2(KEYINPUT35), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT85), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n423), .B2(new_n429), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n399), .A2(new_n348), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n417), .B1(new_n407), .B2(new_n410), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n347), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n399), .A2(KEYINPUT29), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT72), .B1(new_n590), .B2(new_n417), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n419), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n418), .A2(new_n419), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT73), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n415), .A2(new_n416), .A3(new_n420), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n596), .A2(new_n341), .B1(new_n426), .B2(new_n428), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n584), .ZN(new_n598));
  INV_X1    g397(.A(new_n504), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n503), .B2(KEYINPUT88), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT88), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n497), .A2(new_n501), .A3(new_n601), .A4(new_n502), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT35), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AND4_X1   g402(.A1(new_n586), .A2(new_n579), .A3(new_n598), .A4(new_n603), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n582), .A2(new_n583), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n546), .A2(new_n552), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT80), .B1(new_n597), .B2(new_n505), .ZN(new_n608));
  AND4_X1   g407(.A1(KEYINPUT80), .A2(new_n423), .A3(new_n429), .A4(new_n505), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n572), .A2(new_n578), .ZN(new_n611));
  NAND2_X1  g410(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n612));
  OR2_X1    g411(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n572), .A2(new_n578), .A3(KEYINPUT70), .A4(KEYINPUT36), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618));
  INV_X1    g417(.A(new_n481), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n482), .A2(new_n484), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n618), .B(new_n489), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n621), .A2(KEYINPUT86), .A3(new_n434), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT86), .B1(new_n621), .B2(new_n434), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n489), .B1(new_n619), .B2(new_n620), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n490), .A2(new_n491), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n625), .B(KEYINPUT39), .C1(new_n489), .C2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(KEYINPUT40), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n628), .A2(new_n501), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n627), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT87), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n423), .A2(new_n429), .A3(new_n584), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n633), .B(new_n634), .C1(new_n585), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT89), .B(KEYINPUT38), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n341), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n419), .B1(new_n409), .B2(new_n414), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n418), .B2(new_n346), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n415), .A2(new_n641), .A3(new_n420), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n600), .A2(new_n425), .A3(new_n602), .A4(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT37), .B1(new_n421), .B2(new_n422), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n644), .A2(new_n341), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n638), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n606), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n632), .B(new_n629), .C1(new_n635), .C2(new_n585), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(KEYINPUT87), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n617), .B1(new_n636), .B2(new_n652), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n301), .B(new_n338), .C1(new_n605), .C2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT90), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n604), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n581), .A2(KEYINPUT90), .A3(KEYINPUT35), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n636), .ZN(new_n662));
  INV_X1    g461(.A(new_n617), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n301), .A4(new_n338), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n656), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n505), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT104), .B(G1gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1324gat));
  NOR2_X1   g470(.A1(new_n635), .A2(new_n585), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(G8gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n656), .B2(new_n666), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT105), .B(KEYINPUT16), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G8gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(KEYINPUT42), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT42), .B1(new_n676), .B2(new_n678), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n675), .B(new_n679), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n673), .A3(new_n678), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(KEYINPUT106), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n675), .A2(new_n679), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(KEYINPUT106), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n680), .A2(new_n681), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n692), .ZN(G1325gat));
  AOI21_X1  g492(.A(G15gat), .B1(new_n667), .B2(new_n611), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n614), .A2(new_n615), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n667), .B2(new_n696), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n667), .A2(new_n607), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n700), .B2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1327gat));
  AOI21_X1  g505(.A(new_n322), .B1(new_n661), .B2(new_n664), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n254), .A2(new_n300), .A3(new_n336), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n505), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n708), .B(KEYINPUT111), .Z(new_n713));
  NAND2_X1  g512(.A1(new_n665), .A2(new_n323), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(KEYINPUT44), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n505), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n712), .A2(new_n720), .ZN(G1328gat));
  NOR3_X1   g520(.A1(new_n709), .A2(G36gat), .A3(new_n672), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n719), .B2(new_n672), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  AOI21_X1  g524(.A(new_n226), .B1(new_n718), .B2(new_n695), .ZN(new_n726));
  INV_X1    g525(.A(new_n709), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n727), .A2(new_n226), .A3(new_n611), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n606), .B1(new_n709), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n731), .B2(new_n709), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n224), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n718), .A2(G50gat), .A3(new_n607), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n734), .A2(KEYINPUT48), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT48), .B1(new_n734), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  INV_X1    g537(.A(new_n300), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n253), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n665), .A2(new_n338), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n668), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n741), .B(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(new_n673), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  INV_X1    g551(.A(new_n611), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n741), .A2(KEYINPUT114), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT114), .B1(new_n741), .B2(new_n753), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(G71gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n746), .A2(new_n695), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n752), .B(new_n758), .C1(new_n759), .C2(new_n757), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n746), .B2(new_n695), .ZN(new_n761));
  AOI21_X1  g560(.A(G71gat), .B1(new_n754), .B2(new_n755), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT50), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n760), .A2(new_n763), .ZN(G1334gat));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n607), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g565(.A1(new_n715), .A2(new_n717), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n254), .A2(new_n337), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT115), .Z(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n739), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n505), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n714), .B2(new_n769), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n769), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n707), .A2(KEYINPUT51), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n300), .A2(new_n264), .A3(new_n668), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n771), .B2(new_n672), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n672), .A2(G92gat), .A3(new_n739), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n782), .B(new_n783), .C1(new_n779), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n775), .A2(KEYINPUT116), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n774), .A2(new_n788), .A3(new_n777), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n789), .A3(new_n784), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n782), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n791), .B2(new_n783), .ZN(G1337gat));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n300), .A2(new_n793), .A3(new_n611), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT117), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n775), .B2(new_n778), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n771), .A2(new_n616), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n793), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT118), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n800), .B(new_n796), .C1(new_n797), .C2(new_n793), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1338gat));
  OAI21_X1  g601(.A(G106gat), .B1(new_n771), .B2(new_n606), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n739), .A2(new_n606), .A3(G106gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n803), .B(new_n804), .C1(new_n779), .C2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n789), .A3(new_n805), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n803), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(new_n804), .ZN(G1339gat));
  NAND4_X1  g609(.A1(new_n246), .A2(new_n207), .A3(new_n248), .A4(new_n251), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n249), .A2(new_n250), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n243), .B1(new_n241), .B2(new_n242), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n206), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n300), .A2(new_n816), .B1(new_n317), .B2(new_n321), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n293), .B(new_n286), .C1(new_n289), .C2(KEYINPUT10), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n292), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n257), .B1(new_n292), .B2(KEYINPUT54), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR3_X1    g621(.A1(new_n820), .A2(new_n821), .A3(new_n818), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n296), .A2(new_n258), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n253), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n336), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n822), .A3(new_n824), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n323), .B1(new_n827), .B2(new_n815), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n253), .A2(new_n300), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n826), .A2(new_n828), .B1(new_n338), .B2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n607), .A3(new_n753), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(new_n668), .A3(new_n672), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n253), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n300), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g635(.A1(new_n832), .A2(new_n336), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT119), .B(G127gat), .Z(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(G1342gat));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n832), .B(new_n323), .C1(new_n840), .C2(new_n441), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n441), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(G1343gat));
  NOR3_X1   g642(.A1(new_n673), .A2(new_n505), .A3(new_n695), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n828), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n338), .A2(new_n829), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n847), .B2(new_n607), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n830), .A2(new_n849), .A3(new_n606), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n844), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n254), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n830), .A2(new_n606), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n844), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n451), .A3(new_n253), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n847), .A2(KEYINPUT57), .A3(new_n607), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n849), .B1(new_n830), .B2(new_n606), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n844), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n254), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n858), .B1(new_n865), .B2(new_n451), .ZN(new_n866));
  INV_X1    g665(.A(new_n864), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT120), .B1(new_n863), .B2(new_n844), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n253), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT121), .A3(G141gat), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n866), .A2(new_n870), .A3(new_n856), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n857), .B1(new_n871), .B2(new_n853), .ZN(G1344gat));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n453), .A3(new_n300), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT122), .B1(new_n861), .B2(new_n862), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n862), .A2(KEYINPUT122), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n300), .A3(new_n844), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n874), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n860), .A2(new_n864), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT59), .B(new_n453), .C1(new_n881), .C2(new_n300), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n873), .B1(new_n880), .B2(new_n882), .ZN(G1345gat));
  AOI21_X1  g682(.A(G155gat), .B1(new_n855), .B2(new_n336), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n336), .A2(G155gat), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT123), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n881), .B2(new_n886), .ZN(G1346gat));
  NAND3_X1  g686(.A1(new_n855), .A2(new_n461), .A3(new_n323), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n322), .B1(new_n860), .B2(new_n864), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n461), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n672), .A2(new_n668), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n831), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n253), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n300), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n336), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n328), .ZN(new_n898));
  OAI221_X1 g697(.A(new_n898), .B1(KEYINPUT124), .B2(KEYINPUT60), .C1(new_n373), .C2(new_n897), .ZN(new_n899));
  NAND2_X1  g698(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n899), .B(new_n900), .ZN(G1350gat));
  NAND2_X1  g700(.A1(new_n892), .A2(new_n323), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G190gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(KEYINPUT125), .A3(KEYINPUT61), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(KEYINPUT61), .B2(new_n903), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT125), .B1(new_n903), .B2(KEYINPUT61), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n905), .A2(new_n906), .B1(G190gat), .B2(new_n902), .ZN(G1351gat));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n616), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n854), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT126), .Z(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n203), .A3(new_n253), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n877), .A2(new_n908), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n253), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n203), .ZN(G1352gat));
  NAND3_X1  g715(.A1(new_n878), .A2(new_n300), .A3(new_n909), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G204gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n910), .A2(G204gat), .A3(new_n739), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT62), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1353gat));
  INV_X1    g720(.A(G211gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n911), .A2(new_n922), .A3(new_n336), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n913), .A2(new_n336), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n924), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT63), .B1(new_n924), .B2(G211gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(G1354gat));
  AOI21_X1  g726(.A(G218gat), .B1(new_n911), .B2(new_n323), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n323), .A2(G218gat), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT127), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n913), .B2(new_n930), .ZN(G1355gat));
endmodule


