//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  NAND2_X1  g000(.A1(KEYINPUT82), .A2(G104), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT82), .A2(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT3), .A2(G107), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n188), .A2(new_n189), .A3(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT3), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n191), .B2(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT82), .A2(G104), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n195), .A3(new_n187), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(G104), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .A4(new_n192), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT4), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n205), .B(G101), .C1(new_n191), .C2(new_n197), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G119), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n211), .A3(G116), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n208), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G113), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n212), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n212), .A2(new_n219), .A3(KEYINPUT68), .A4(new_n214), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n212), .A2(new_n214), .ZN(new_n224));
  INV_X1    g038(.A(new_n219), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT84), .B1(new_n207), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n225), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT67), .B(G119), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n213), .B1(new_n229), .B2(G116), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT68), .B1(new_n230), .B2(new_n219), .ZN(new_n231));
  INV_X1    g045(.A(new_n223), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT84), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n206), .A4(new_n204), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n227), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n223), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n199), .A2(new_n194), .A3(new_n187), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n201), .B1(G104), .B2(G107), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n203), .A2(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT85), .B(KEYINPUT5), .Z(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(G116), .A3(new_n229), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G113), .C1(new_n224), .C2(new_n242), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n237), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT86), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n237), .A2(new_n241), .A3(new_n244), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n236), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G110), .B(G122), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n236), .A2(new_n249), .A3(new_n251), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(KEYINPUT6), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n259), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n262), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT64), .B1(new_n270), .B2(new_n266), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n262), .B2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n270), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n269), .A2(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n265), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  INV_X1    g091(.A(G224), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI221_X1 g094(.A(new_n265), .B1(new_n278), .B2(G953), .C1(new_n276), .C2(new_n264), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n250), .A2(new_n283), .A3(new_n252), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n255), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n279), .A2(KEYINPUT7), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n280), .B2(new_n281), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n203), .A2(new_n240), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n237), .A2(new_n244), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT5), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n243), .B(G113), .C1(new_n291), .C2(new_n224), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n237), .B2(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n251), .B(KEYINPUT8), .Z(new_n294));
  NOR3_X1   g108(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n277), .A2(new_n287), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n288), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n297), .B2(new_n254), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n285), .A2(new_n286), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT87), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n285), .A2(new_n301), .A3(new_n298), .A4(new_n286), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n285), .A2(new_n298), .ZN(new_n303));
  INV_X1    g117(.A(new_n286), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT91), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n264), .A2(G140), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT74), .ZN(new_n313));
  OR3_X1    g127(.A1(new_n264), .A2(KEYINPUT74), .A3(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  NOR2_X1   g133(.A1(G237), .A2(G953), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(G143), .A3(G214), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(G143), .B1(new_n320), .B2(G214), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n323), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n321), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT17), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n315), .A2(new_n257), .A3(new_n317), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n321), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT17), .A3(G131), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n319), .A2(new_n329), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n313), .A2(G146), .A3(new_n314), .ZN(new_n334));
  AND4_X1   g148(.A1(KEYINPUT76), .A2(new_n311), .A3(new_n312), .A4(new_n257), .ZN(new_n335));
  XNOR2_X1  g149(.A(G125), .B(G140), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT76), .B1(new_n336), .B2(new_n257), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n331), .A2(KEYINPUT18), .A3(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT18), .A2(G131), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n325), .A2(new_n321), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT89), .B(G104), .Z(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n333), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT90), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n333), .A2(new_n342), .A3(new_n349), .A4(new_n346), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n324), .A2(new_n327), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT19), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n313), .B2(new_n314), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n336), .A2(KEYINPUT19), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n257), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n319), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n342), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT88), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n360), .A3(new_n342), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n345), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n309), .B1(new_n351), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G475), .A2(G902), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n351), .A2(new_n362), .A3(new_n309), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n351), .A2(new_n362), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n365), .A2(KEYINPUT92), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n365), .A2(KEYINPUT92), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT20), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n367), .A2(KEYINPUT20), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n333), .A2(new_n342), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n351), .B1(new_n346), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G902), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n376), .A2(G475), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(G234), .A2(G237), .ZN(new_n379));
  INV_X1    g193(.A(G953), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(G952), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(G902), .A3(G953), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT21), .B(G898), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT15), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G478), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT9), .B(G234), .ZN(new_n390));
  INV_X1    g204(.A(G217), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(new_n391), .A3(G953), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G122), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT93), .B1(new_n394), .B2(G116), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n396));
  INV_X1    g210(.A(G116), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT14), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(G116), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n399), .A2(KEYINPUT14), .ZN(new_n403));
  OAI21_X1  g217(.A(G107), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n399), .A2(new_n401), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n260), .A2(G128), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n260), .A2(G128), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n407), .A2(G134), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G134), .B1(new_n407), .B2(new_n408), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n405), .A2(new_n194), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT13), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n406), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT94), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n406), .B2(new_n413), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n406), .A2(new_n415), .A3(new_n413), .ZN(new_n418));
  OAI21_X1  g232(.A(G134), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n405), .A2(new_n194), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n399), .A2(new_n194), .A3(new_n401), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n419), .B(new_n409), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT95), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n412), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n412), .B2(new_n422), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n393), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n412), .A2(new_n422), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT95), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n392), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(KEYINPUT96), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT96), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n432), .B(G902), .C1(new_n426), .C2(new_n429), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n389), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n433), .A2(new_n389), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n378), .A2(new_n387), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  INV_X1    g254(.A(G227), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n440), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n276), .A2(new_n204), .A3(new_n206), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n259), .B(new_n270), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n241), .A2(KEYINPUT10), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT10), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n263), .B2(new_n289), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT83), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT69), .ZN(new_n452));
  INV_X1    g266(.A(G134), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT11), .B1(new_n453), .B2(G137), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT11), .ZN(new_n455));
  INV_X1    g269(.A(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(G134), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT66), .B1(new_n456), .B2(G134), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT66), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n453), .A3(G137), .ZN(new_n461));
  AND4_X1   g275(.A1(new_n326), .A2(new_n458), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n459), .A2(new_n461), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n326), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n452), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G131), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n326), .A3(new_n458), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(KEYINPUT69), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n445), .A2(new_n447), .A3(new_n449), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n451), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n450), .A2(new_n470), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n444), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n241), .A2(new_n446), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n263), .A2(new_n289), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n469), .B(new_n465), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT12), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n263), .B(new_n289), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n462), .A2(new_n464), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(new_n480), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n484), .A2(new_n474), .A3(new_n443), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n439), .B(new_n375), .C1(new_n476), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n473), .A2(new_n475), .A3(new_n444), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n443), .B1(new_n484), .B2(new_n474), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(G469), .ZN(new_n489));
  NAND2_X1  g303(.A1(G469), .A2(G902), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G221), .B1(new_n390), .B2(G902), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n308), .A2(new_n438), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(G472), .A2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT32), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n465), .A2(new_n276), .A3(new_n469), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n453), .A2(G137), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n456), .A2(G134), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n446), .A2(new_n468), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n501), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n505), .ZN(new_n509));
  INV_X1    g323(.A(new_n276), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n510), .B2(new_n482), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n508), .A2(new_n233), .A3(new_n509), .A4(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n501), .A2(new_n226), .A3(new_n505), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n320), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n514), .A2(new_n515), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n515), .B1(new_n514), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n501), .A2(new_n505), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT28), .A3(new_n226), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n511), .A2(new_n233), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT28), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n520), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT71), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n514), .A2(new_n521), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT31), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n514), .A2(new_n515), .A3(new_n521), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n535), .A2(KEYINPUT71), .A3(new_n532), .A4(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n500), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n497), .B1(new_n533), .B2(new_n538), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n499), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n535), .A2(new_n532), .A3(new_n536), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n537), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n516), .B2(new_n528), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n525), .A2(new_n226), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n529), .A3(new_n526), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT29), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n531), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n530), .A2(new_n520), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n514), .A2(new_n531), .A3(new_n516), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n556), .B1(KEYINPUT29), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G472), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n541), .A2(new_n543), .A3(new_n548), .A4(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n337), .A2(new_n335), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n319), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n208), .A2(new_n256), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n229), .B2(new_n256), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT24), .B(G110), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G110), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n229), .B2(G128), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n570), .B(new_n572), .C1(new_n566), .C2(new_n571), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n573), .A3(KEYINPUT75), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n564), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n572), .B1(new_n566), .B2(new_n571), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G110), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n568), .B2(new_n567), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n319), .A2(new_n330), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT22), .B(G137), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n380), .A2(G221), .A3(G234), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(KEYINPUT77), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n578), .B2(new_n584), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n596), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n589), .A2(new_n591), .A3(new_n598), .A4(new_n594), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n391), .B1(G234), .B2(new_n375), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT79), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT79), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n597), .A2(new_n603), .A3(new_n599), .A4(new_n600), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n589), .A2(new_n591), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n600), .A2(G902), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT80), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n602), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n562), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT81), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT73), .B1(new_n547), .B2(new_n500), .ZN(new_n613));
  INV_X1    g427(.A(new_n500), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n540), .B(new_n614), .C1(new_n546), .C2(new_n537), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n542), .A2(new_n499), .B1(G472), .B2(new_n560), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n609), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT81), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n496), .B1(new_n612), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n201), .ZN(G3));
  AOI21_X1  g436(.A(new_n498), .B1(new_n546), .B2(new_n537), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n547), .A2(new_n375), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(G472), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n494), .A2(new_n609), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(KEYINPUT97), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n546), .B2(new_n537), .ZN(new_n629));
  INV_X1    g443(.A(G472), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n542), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n493), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n305), .A2(new_n299), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n307), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT33), .B1(new_n426), .B2(new_n429), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n427), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n393), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n427), .A2(new_n640), .A3(new_n392), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(G478), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(G902), .ZN(new_n647));
  INV_X1    g461(.A(new_n430), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n645), .A2(new_n647), .B1(new_n648), .B2(new_n646), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n387), .C1(new_n372), .C2(new_n377), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n637), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n635), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT99), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  INV_X1    g470(.A(new_n366), .ZN(new_n657));
  INV_X1    g471(.A(new_n365), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n657), .A2(new_n363), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT20), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n367), .A2(KEYINPUT20), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n377), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n436), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n664), .A2(new_n637), .A3(new_n386), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n635), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NOR2_X1   g482(.A1(new_n308), .A2(new_n494), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n579), .A2(new_n585), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n607), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n602), .A2(new_n604), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n438), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n669), .A2(new_n676), .A3(new_n625), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  NOR2_X1   g493(.A1(new_n637), .A2(new_n494), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n384), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT100), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(KEYINPUT100), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n381), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n664), .A2(new_n675), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n562), .A2(new_n680), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  OAI21_X1  g503(.A(new_n436), .B1(new_n372), .B2(new_n377), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n685), .B(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n493), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n691), .B(new_n307), .C1(new_n695), .C2(KEYINPUT40), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(KEYINPUT40), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n541), .A2(new_n548), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n551), .A2(new_n531), .A3(new_n516), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n375), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n531), .B1(new_n514), .B2(new_n516), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n702), .B1(new_n623), .B2(KEYINPUT32), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n306), .B(KEYINPUT38), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n697), .A2(new_n705), .A3(new_n675), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  NAND2_X1  g522(.A1(new_n368), .A2(new_n371), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n659), .B2(new_n660), .ZN(new_n710));
  INV_X1    g524(.A(new_n377), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n649), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n685), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n675), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n561), .B1(new_n623), .B2(KEYINPUT32), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n714), .B(new_n680), .C1(new_n698), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  OR2_X1    g531(.A1(new_n476), .A2(new_n485), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n375), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n492), .A3(new_n486), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n562), .A2(new_n610), .A3(new_n652), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT102), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n723), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n562), .A2(new_n610), .A3(new_n665), .A4(new_n722), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR2_X1   g542(.A1(new_n637), .A2(new_n721), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n562), .A2(new_n676), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NOR2_X1   g545(.A1(new_n553), .A2(new_n520), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n535), .A2(new_n536), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n497), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n624), .B2(G472), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n637), .A2(new_n690), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n721), .A2(new_n386), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n610), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  OAI211_X1 g554(.A(new_n674), .B(new_n734), .C1(new_n629), .C2(new_n630), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n713), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n729), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  AND3_X1   g558(.A1(new_n300), .A2(new_n302), .A3(new_n305), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n489), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT103), .A4(G469), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n486), .A3(new_n490), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n492), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n745), .A2(KEYINPUT104), .A3(new_n307), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n300), .A2(new_n305), .A3(new_n307), .A4(new_n302), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n753), .B1(new_n754), .B2(new_n750), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n713), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n562), .A3(new_n610), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT105), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n618), .A2(new_n761), .A3(new_n757), .A4(new_n756), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n543), .A2(new_n539), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT106), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n543), .A2(new_n766), .A3(new_n539), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n561), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n713), .A2(new_n760), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n610), .A3(new_n756), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NOR2_X1   g586(.A1(new_n664), .A2(new_n686), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n618), .A2(new_n773), .A3(new_n756), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  NAND2_X1  g589(.A1(new_n378), .A2(new_n650), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT43), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n625), .B2(new_n675), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n631), .A2(KEYINPUT108), .A3(new_n674), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n781), .A3(KEYINPUT44), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n487), .A2(new_n488), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n439), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(new_n490), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n486), .B1(new_n791), .B2(KEYINPUT46), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n492), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n693), .A3(new_n754), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n786), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  XOR2_X1   g611(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n794), .B(new_n798), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n713), .A2(new_n610), .A3(new_n754), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n799), .A2(new_n562), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n310), .ZN(G42));
  NAND2_X1  g616(.A1(new_n736), .A2(new_n610), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n777), .A2(new_n803), .A3(new_n381), .ZN(new_n804));
  INV_X1    g618(.A(new_n307), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n722), .B(new_n805), .C1(KEYINPUT114), .C2(KEYINPUT50), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n706), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n741), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n777), .A2(new_n381), .A3(new_n721), .A4(new_n754), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n720), .A2(new_n486), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n799), .B1(new_n492), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n804), .A2(new_n754), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n816), .A2(new_n817), .B1(new_n808), .B2(new_n810), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n754), .A2(new_n721), .A3(new_n609), .A4(new_n381), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n704), .A2(new_n819), .A3(new_n378), .A4(new_n649), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT115), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n814), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT51), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n768), .A2(new_n610), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n813), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT48), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n704), .A2(new_n819), .A3(new_n712), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(G952), .A3(new_n380), .ZN(new_n828));
  INV_X1    g642(.A(new_n804), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(new_n729), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT116), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT111), .B1(new_n308), .B2(new_n651), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n437), .A2(new_n372), .A3(new_n377), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n387), .A3(new_n307), .A4(new_n306), .ZN(new_n836));
  INV_X1    g650(.A(new_n651), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n307), .A4(new_n306), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n834), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n727), .B1(new_n840), .B2(new_n634), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n723), .A2(new_n730), .A3(new_n677), .A4(new_n739), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n621), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n562), .A2(new_n756), .A3(new_n610), .A4(new_n773), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n756), .A2(new_n742), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n436), .A2(new_n686), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n493), .A3(new_n663), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n675), .A3(new_n754), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n562), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n844), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n846), .A4(new_n850), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n843), .A2(new_n771), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n749), .A2(new_n492), .A3(new_n685), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n637), .A2(new_n690), .A3(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n675), .B(new_n858), .C1(new_n698), .C2(new_n703), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n688), .A2(new_n716), .A3(new_n859), .A4(new_n743), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT113), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n562), .B(new_n680), .C1(new_n687), .C2(new_n714), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(KEYINPUT52), .A3(new_n743), .A4(new_n859), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n862), .B(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n856), .A2(new_n866), .A3(KEYINPUT53), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n860), .A2(new_n861), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n864), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n843), .A2(new_n771), .A3(new_n854), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n867), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n856), .A2(new_n866), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n872), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n877), .B2(new_n868), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n833), .A2(new_n878), .B1(G952), .B2(G953), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n815), .A2(KEYINPUT49), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT110), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n492), .A2(new_n307), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n815), .B2(KEYINPUT49), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n610), .ZN(new_n884));
  OR4_X1    g698(.A1(new_n706), .A2(new_n881), .A3(new_n776), .A4(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n879), .B1(new_n705), .B2(new_n885), .ZN(G75));
  NAND2_X1  g700(.A1(new_n867), .A2(new_n873), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(G210), .A3(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n255), .A2(new_n284), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT117), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT118), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n282), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n888), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n888), .B2(new_n889), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n380), .A2(G952), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G51));
  XOR2_X1   g712(.A(new_n490), .B(KEYINPUT57), .Z(new_n899));
  INV_X1    g713(.A(new_n874), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n868), .B1(new_n867), .B2(new_n873), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n718), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n887), .A2(G902), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n904), .A2(new_n790), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n897), .B1(new_n903), .B2(new_n905), .ZN(G54));
  NOR2_X1   g720(.A1(new_n657), .A2(new_n363), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(KEYINPUT58), .A2(G475), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n897), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(G60));
  XOR2_X1   g728(.A(new_n645), .B(KEYINPUT119), .Z(new_n915));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT59), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n915), .B(new_n917), .C1(new_n900), .C2(new_n901), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n911), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n878), .B2(new_n917), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT60), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n862), .A2(new_n865), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n860), .A2(KEYINPUT113), .A3(new_n861), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n926), .A2(new_n855), .A3(new_n872), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n871), .A2(new_n872), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n605), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n897), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT121), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n887), .A2(new_n932), .A3(new_n672), .A4(new_n923), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n672), .B(new_n923), .C1(new_n927), .C2(new_n928), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n931), .A2(KEYINPUT61), .A3(new_n934), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(G66));
  NOR3_X1   g754(.A1(new_n385), .A2(new_n278), .A3(new_n380), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n843), .B2(new_n380), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n891), .B1(G898), .B2(new_n380), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT122), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(G69));
  NAND2_X1  g759(.A1(new_n612), .A2(new_n620), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n835), .A2(new_n712), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n947), .A2(new_n695), .A3(new_n754), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n801), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n863), .A2(new_n743), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n707), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n796), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n951), .A2(new_n955), .A3(new_n707), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT124), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n380), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n794), .A2(new_n693), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n824), .A2(new_n737), .A3(new_n961), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT125), .Z(new_n963));
  NOR3_X1   g777(.A1(new_n801), .A2(new_n845), .A3(new_n950), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n771), .A3(new_n796), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n380), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n508), .A2(new_n509), .A3(new_n513), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n354), .A2(new_n355), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n681), .B2(G953), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n960), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(G953), .B1(new_n441), .B2(new_n681), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n958), .A2(KEYINPUT123), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n969), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n971), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G72));
  INV_X1    g791(.A(new_n843), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n954), .A2(new_n978), .A3(new_n957), .ZN(new_n979));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n701), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n965), .A2(new_n978), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n982), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n911), .B(new_n983), .C1(new_n985), .C2(new_n558), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n558), .A2(new_n981), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n877), .A2(new_n701), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n986), .A2(new_n988), .ZN(G57));
endmodule


