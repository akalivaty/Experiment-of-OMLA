//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT88), .ZN(new_n205));
  XOR2_X1   g004(.A(G169gat), .B(G197gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT12), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n207), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT89), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT89), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n216), .A2(KEYINPUT15), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT14), .ZN(new_n222));
  NAND2_X1  g021(.A1(G29gat), .A2(G36gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT92), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G43gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT91), .B(G50gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT90), .B(G43gat), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n226), .A2(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n220), .B(new_n225), .C1(KEYINPUT15), .C2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n216), .A2(KEYINPUT15), .ZN(new_n232));
  INV_X1    g031(.A(new_n223), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n222), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(new_n219), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G15gat), .B(G22gat), .ZN(new_n237));
  INV_X1    g036(.A(G1gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT16), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n238), .B2(new_n237), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(G8gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n231), .A2(new_n235), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT17), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n231), .A2(new_n235), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n247), .B2(new_n241), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT18), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n231), .A2(new_n235), .A3(new_n245), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n245), .B1(new_n231), .B2(new_n235), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n241), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n241), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n243), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n253), .A2(KEYINPUT18), .A3(new_n249), .A4(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n249), .B(KEYINPUT13), .Z(new_n257));
  NOR2_X1   g056(.A1(new_n254), .A2(new_n243), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n242), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n214), .B1(new_n250), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT18), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(new_n255), .ZN(new_n263));
  INV_X1    g062(.A(new_n249), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n265), .A2(new_n256), .A3(new_n213), .A4(new_n259), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G211gat), .B(G218gat), .ZN(new_n270));
  INV_X1    g069(.A(G204gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G197gat), .ZN(new_n272));
  INV_X1    g071(.A(G197gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G204gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n277));
  OAI21_X1  g076(.A(G211gat), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n270), .B1(new_n280), .B2(KEYINPUT78), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT78), .ZN(new_n282));
  AOI211_X1 g081(.A(new_n282), .B(new_n275), .C1(new_n278), .C2(new_n279), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n287), .A2(new_n282), .A3(new_n270), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT79), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n282), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n280), .A2(KEYINPUT78), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n270), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n281), .A2(new_n283), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT79), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G226gat), .A2(G233gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT26), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303));
  NAND2_X1  g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n306), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G190gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT27), .B1(new_n306), .B2(KEYINPUT69), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT28), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT27), .B(G183gat), .Z(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n311), .A2(new_n312), .A3(G190gat), .ZN(new_n313));
  OAI221_X1 g112(.A(new_n299), .B1(new_n302), .B2(new_n305), .C1(new_n310), .C2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT23), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n304), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n321), .A3(new_n304), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT25), .B1(new_n300), .B2(KEYINPUT23), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT24), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT67), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT67), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT24), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n326), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n315), .B1(new_n323), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n329), .A2(KEYINPUT24), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n327), .A2(KEYINPUT67), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n299), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n333), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n324), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n318), .A2(new_n321), .A3(new_n304), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n321), .B1(new_n318), .B2(new_n304), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n343), .A3(KEYINPUT68), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT64), .B1(new_n326), .B2(KEYINPUT24), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT64), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n299), .A2(new_n348), .A3(new_n327), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n333), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n301), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n304), .A3(new_n318), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n345), .B(new_n346), .C1(new_n350), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n344), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n346), .B1(new_n350), .B2(new_n353), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n356), .A2(KEYINPUT65), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n314), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n298), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(KEYINPUT65), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n361), .A2(new_n354), .A3(new_n335), .A4(new_n344), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n297), .B1(new_n362), .B2(new_n314), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n296), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G8gat), .B(G36gat), .Z(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT80), .ZN(new_n366));
  XOR2_X1   g165(.A(G64gat), .B(G92gat), .Z(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n296), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n358), .A2(new_n298), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n362), .B2(new_n314), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n369), .B(new_n370), .C1(new_n298), .C2(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n364), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n368), .B1(new_n364), .B2(new_n372), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n375), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT87), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n372), .ZN(new_n380));
  INV_X1    g179(.A(new_n368), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n368), .A3(new_n372), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(KEYINPUT30), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT87), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n377), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G127gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G134gat), .ZN(new_n390));
  XOR2_X1   g189(.A(KEYINPUT70), .B(G134gat), .Z(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(new_n389), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n393));
  INV_X1    g192(.A(G113gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(G120gat), .ZN(new_n395));
  INV_X1    g194(.A(G120gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(G113gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT71), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n394), .B2(G120gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(KEYINPUT72), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT72), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G113gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n406), .A3(G120gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n409));
  INV_X1    g208(.A(G134gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G127gat), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n390), .B2(new_n411), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n390), .A2(new_n411), .A3(new_n409), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n408), .B(new_n393), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G148gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417));
  INV_X1    g216(.A(G141gat), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(G148gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(G148gat), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT2), .ZN(new_n422));
  INV_X1    g221(.A(G155gat), .ZN(new_n423));
  INV_X1    g222(.A(G162gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n415), .A2(G141gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(G148gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n422), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n423), .A2(new_n424), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n426), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n421), .A2(new_n427), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n399), .A2(new_n414), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n415), .A2(G141gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n428), .B1(new_n438), .B2(new_n417), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n439), .A2(new_n416), .B1(new_n426), .B2(new_n425), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n433), .B1(new_n422), .B2(new_n430), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT82), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n421), .A2(new_n427), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n431), .A2(new_n434), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(KEYINPUT3), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n437), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n414), .A2(new_n435), .A3(new_n399), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n414), .A2(new_n435), .A3(new_n399), .A4(KEYINPUT4), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n388), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n454), .A2(KEYINPUT39), .ZN(new_n455));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT0), .ZN(new_n457));
  XNOR2_X1  g256(.A(G57gat), .B(G85gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  NAND2_X1  g258(.A1(new_n414), .A2(new_n399), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n449), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n463), .A2(new_n388), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n454), .A3(KEYINPUT39), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n455), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n437), .A2(new_n447), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(new_n387), .A3(new_n451), .A4(new_n452), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n463), .A2(new_n388), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n459), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n470), .A2(new_n473), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n468), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n466), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n379), .A2(new_n386), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  XOR2_X1   g282(.A(G78gat), .B(G106gat), .Z(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT31), .B(G50gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G228gat), .A2(G233gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n435), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n359), .B1(new_n489), .B2(KEYINPUT3), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n289), .A2(new_n295), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n292), .A2(new_n293), .A3(new_n359), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n462), .B1(new_n492), .B2(new_n436), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n491), .B1(new_n493), .B2(KEYINPUT85), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n495));
  AOI211_X1 g294(.A(new_n495), .B(new_n462), .C1(new_n492), .C2(new_n436), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n488), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G22gat), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n492), .A2(new_n436), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n487), .B(new_n491), .C1(new_n499), .C2(new_n435), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n498), .B1(new_n497), .B2(new_n500), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n483), .B(new_n486), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(new_n500), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G22gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n486), .A2(new_n483), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n483), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n380), .A2(KEYINPUT37), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(new_n364), .B2(new_n372), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n368), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT38), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT38), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n516), .B(new_n368), .C1(new_n511), .C2(new_n513), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n476), .B1(new_n475), .B2(new_n477), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n478), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n475), .A2(new_n477), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n476), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n374), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n515), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n482), .A2(new_n510), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n358), .A2(new_n461), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n362), .A2(new_n460), .A3(new_n314), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G227gat), .A2(G233gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT34), .ZN(new_n532));
  INV_X1    g331(.A(G227gat), .ZN(new_n533));
  INV_X1    g332(.A(G233gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n526), .B2(new_n527), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT34), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT74), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n532), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n526), .A2(new_n535), .A3(new_n527), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT32), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G15gat), .B(G43gat), .Z(new_n545));
  XNOR2_X1  g344(.A(G71gat), .B(G99gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n547), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n541), .B(KEYINPUT32), .C1(new_n543), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n540), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n532), .A2(new_n538), .A3(new_n539), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n550), .A3(new_n548), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT36), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT75), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n540), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n560), .B2(KEYINPUT36), .ZN(new_n561));
  INV_X1    g360(.A(new_n518), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n562), .A2(KEYINPUT84), .A3(new_n521), .A4(new_n478), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT84), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n520), .B(new_n476), .C1(new_n564), .C2(KEYINPUT6), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n384), .A2(new_n377), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n503), .A2(new_n509), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n525), .A2(new_n561), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n558), .A2(new_n503), .A3(new_n509), .A4(new_n559), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT35), .B1(new_n572), .B2(new_n568), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n379), .A2(new_n386), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n552), .A2(new_n554), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n519), .A2(new_n522), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(KEYINPUT35), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n574), .A2(new_n510), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n269), .B1(new_n571), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G183gat), .B(G211gat), .Z(new_n581));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT96), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT94), .A2(G57gat), .A3(G64gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(KEYINPUT94), .A2(G57gat), .ZN(new_n592));
  INV_X1    g391(.A(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n589), .A2(G71gat), .A3(G78gat), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n591), .B(new_n594), .C1(new_n595), .C2(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  AND2_X1   g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g407(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n602), .A2(new_n603), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n607), .B1(new_n610), .B2(new_n604), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n584), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n608), .B1(new_n605), .B2(new_n606), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n604), .A3(new_n607), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n583), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n254), .B1(new_n601), .B2(KEYINPUT21), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n612), .B2(new_n615), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n581), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n612), .A2(new_n615), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n616), .ZN(new_n623));
  INV_X1    g422(.A(new_n581), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n627));
  XNOR2_X1  g426(.A(G99gat), .B(G106gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT98), .ZN(new_n629));
  NAND2_X1  g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT7), .ZN(new_n631));
  NAND2_X1  g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(G85gat), .ZN(new_n633));
  INV_X1    g432(.A(G92gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(KEYINPUT8), .A2(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n628), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n631), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n251), .B2(new_n252), .ZN(new_n644));
  XNOR2_X1  g443(.A(G190gat), .B(G218gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT99), .ZN(new_n646));
  NAND2_X1  g445(.A1(G232gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n243), .A2(new_n642), .B1(KEYINPUT41), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n644), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n646), .B1(new_n644), .B2(new_n649), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n627), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(KEYINPUT100), .A3(new_n650), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(new_n655), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n627), .B(new_n659), .C1(new_n651), .C2(new_n652), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n626), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n641), .A2(new_n637), .A3(new_n598), .A4(new_n600), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n639), .B1(new_n636), .B2(KEYINPUT101), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n629), .A2(new_n669), .A3(new_n640), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n590), .A2(new_n596), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n667), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n642), .A2(new_n601), .A3(KEYINPUT10), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n666), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n667), .A2(new_n672), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n666), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT103), .ZN(new_n680));
  XOR2_X1   g479(.A(G176gat), .B(G204gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n674), .A2(KEYINPUT102), .A3(new_n675), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n674), .B2(new_n675), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n665), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n677), .A2(new_n666), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n682), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n664), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n580), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n566), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n574), .ZN(new_n696));
  INV_X1    g495(.A(G8gat), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT42), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g499(.A(KEYINPUT42), .B(new_n698), .S(new_n700), .Z(G1325gat));
  OAI21_X1  g500(.A(G15gat), .B1(new_n695), .B2(new_n561), .ZN(new_n702));
  INV_X1    g501(.A(new_n575), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n695), .B2(new_n704), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n691), .A2(new_n569), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT104), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  AND2_X1   g508(.A1(new_n621), .A2(new_n625), .ZN(new_n710));
  INV_X1    g509(.A(new_n689), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n663), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n580), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n566), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT45), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n571), .A2(new_n579), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n571), .A2(new_n579), .A3(KEYINPUT105), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n663), .A2(KEYINPUT44), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n661), .A2(new_n662), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT44), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n267), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n566), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(KEYINPUT106), .ZN(new_n731));
  OAI21_X1  g530(.A(G29gat), .B1(new_n730), .B2(KEYINPUT106), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n716), .B1(new_n731), .B2(new_n732), .ZN(G1328gat));
  NOR3_X1   g532(.A1(new_n714), .A2(G36gat), .A3(new_n574), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n729), .A2(new_n574), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n736), .B2(KEYINPUT107), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n703), .A2(new_n228), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n580), .A2(new_n713), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n561), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n743), .A3(new_n728), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n744), .B2(new_n228), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT47), .B1(new_n741), .B2(KEYINPUT108), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT109), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n745), .B(new_n747), .ZN(G1330gat));
  NAND2_X1  g547(.A1(new_n569), .A2(new_n227), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n714), .A2(new_n510), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n729), .A2(new_n749), .B1(new_n227), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g551(.A1(new_n719), .A2(new_n720), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n664), .A2(new_n267), .A3(new_n711), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n692), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  INV_X1    g557(.A(new_n574), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n761), .B2(new_n760), .ZN(G1333gat));
  OAI21_X1  g563(.A(G71gat), .B1(new_n755), .B2(new_n561), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n703), .A2(G71gat), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n755), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g567(.A1(new_n756), .A2(new_n569), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n626), .A2(new_n267), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n689), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n722), .B2(new_n725), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774), .B2(new_n566), .ZN(new_n775));
  AND4_X1   g574(.A1(KEYINPUT51), .A2(new_n717), .A3(new_n723), .A4(new_n771), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n663), .B1(new_n571), .B2(new_n579), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n778), .B2(new_n771), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n692), .A2(new_n633), .A3(new_n689), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT110), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n775), .B1(new_n782), .B2(new_n784), .ZN(G1336gat));
  NAND3_X1  g584(.A1(new_n759), .A2(new_n634), .A3(new_n689), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n777), .B2(new_n780), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n773), .A2(new_n759), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n789), .B(new_n791), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n774), .B2(new_n561), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n703), .A2(G99gat), .A3(new_n711), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n782), .B2(new_n794), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n510), .A2(G106gat), .A3(new_n711), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n776), .B2(new_n779), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n510), .B(new_n772), .C1(new_n722), .C2(new_n725), .ZN(new_n799));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n796), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n797), .C1(new_n776), .C2(new_n779), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n802), .B(new_n804), .C1(new_n799), .C2(new_n800), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT113), .B1(new_n805), .B2(KEYINPUT53), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n801), .B1(new_n806), .B2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n682), .B1(new_n676), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n674), .A2(new_n675), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT102), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n674), .A2(KEYINPUT102), .A3(new_n675), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n666), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n674), .A2(new_n666), .A3(new_n675), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT54), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n809), .B(new_n811), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n818), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n686), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n809), .B1(new_n822), .B2(new_n811), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n267), .B(new_n688), .C1(new_n820), .C2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n248), .A2(new_n249), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n242), .A2(new_n258), .A3(new_n257), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n210), .B(new_n208), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n689), .A2(new_n266), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n723), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n688), .B1(new_n820), .B2(new_n823), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n266), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n830), .A2(new_n663), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n710), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n626), .A2(new_n727), .A3(new_n663), .A4(new_n711), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(new_n692), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n574), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n572), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(new_n404), .A3(new_n406), .A4(new_n267), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n703), .A2(new_n569), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n841), .A2(new_n845), .A3(new_n269), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(new_n394), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n842), .B2(new_n689), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n841), .A2(new_n845), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n711), .A2(new_n396), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1341gat));
  NAND3_X1  g650(.A1(new_n842), .A2(new_n389), .A3(new_n626), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n841), .A2(new_n845), .A3(new_n710), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n389), .ZN(G1342gat));
  NOR2_X1   g653(.A1(new_n759), .A2(new_n663), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n391), .A3(new_n572), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n856), .B2(new_n845), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n743), .A2(new_n510), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n839), .A3(new_n692), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT118), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(new_n839), .A3(new_n867), .A4(new_n692), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n759), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n269), .A2(G141gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n743), .A2(new_n759), .A3(new_n566), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n836), .A2(new_n569), .A3(new_n838), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n828), .B1(new_n269), .B2(new_n830), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n832), .B1(new_n877), .B2(new_n663), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n626), .ZN(new_n879));
  INV_X1    g678(.A(new_n834), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT57), .B(new_n569), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n874), .B1(new_n873), .B2(new_n875), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n872), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G141gat), .B1(new_n884), .B2(new_n269), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AND4_X1   g686(.A1(new_n574), .A2(new_n840), .A3(new_n870), .A4(new_n864), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n267), .B(new_n872), .C1(new_n882), .C2(new_n883), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(G141gat), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n886), .B2(new_n890), .ZN(G1344gat));
  OAI211_X1 g690(.A(new_n689), .B(new_n872), .C1(new_n882), .C2(new_n883), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n415), .A2(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n690), .A2(new_n269), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n875), .B(new_n569), .C1(new_n879), .C2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n901), .A2(new_n689), .A3(new_n872), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n897), .B1(new_n902), .B2(new_n415), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n892), .A2(KEYINPUT119), .A3(new_n893), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n896), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n869), .A2(new_n415), .A3(new_n689), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1345gat));
  NAND3_X1  g706(.A1(new_n869), .A2(new_n423), .A3(new_n626), .ZN(new_n908));
  OAI21_X1  g707(.A(G155gat), .B1(new_n884), .B2(new_n710), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n884), .B2(new_n663), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n866), .A2(new_n868), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n424), .A3(new_n855), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n574), .A2(new_n692), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n839), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n844), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n269), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT121), .ZN(new_n919));
  INV_X1    g718(.A(new_n572), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n316), .A3(new_n267), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n317), .A3(new_n689), .ZN(new_n924));
  OAI21_X1  g723(.A(G176gat), .B1(new_n917), .B2(new_n711), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  INV_X1    g725(.A(new_n311), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n927), .A3(new_n626), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n917), .B2(new_n710), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g729(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(G1350gat));
  INV_X1    g731(.A(G190gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n921), .A2(new_n933), .A3(new_n723), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n844), .A3(new_n723), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G190gat), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT123), .B1(new_n936), .B2(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n936), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n561), .A2(new_n915), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n901), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(new_n273), .A3(new_n269), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n916), .A2(new_n862), .ZN(new_n946));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n267), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n901), .A2(new_n689), .A3(new_n943), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G204gat), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n946), .A2(KEYINPUT124), .A3(new_n271), .A4(new_n689), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n916), .A2(new_n862), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n689), .A2(new_n271), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n951), .A2(KEYINPUT62), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT62), .B1(new_n951), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n950), .B1(new_n956), .B2(new_n957), .ZN(G1353gat));
  INV_X1    g757(.A(G211gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n946), .A2(new_n959), .A3(new_n626), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n898), .A2(new_n626), .A3(new_n900), .A4(new_n943), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT125), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n960), .B(new_n966), .C1(new_n962), .C2(new_n963), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1354gat));
  INV_X1    g767(.A(G218gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n969), .B1(new_n953), .B2(new_n663), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g771(.A(KEYINPUT126), .B(new_n969), .C1(new_n953), .C2(new_n663), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n944), .B(KEYINPUT127), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n276), .A2(new_n277), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n663), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n975), .B2(new_n977), .ZN(G1355gat));
endmodule


