//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  AOI21_X1  g003(.A(G101), .B1(new_n188), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n190), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n190), .A3(new_n193), .A4(KEYINPUT76), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n199));
  XNOR2_X1  g013(.A(G104), .B(G107), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n188), .A2(G107), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n192), .A2(G104), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT77), .B(G101), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G116), .ZN(new_n211));
  INV_X1    g025(.A(G116), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G116), .B(G119), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(G113), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n196), .A2(new_n197), .B1(new_n202), .B2(new_n205), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT79), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n209), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n209), .A2(KEYINPUT81), .A3(new_n224), .A4(new_n222), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n189), .B(new_n193), .C1(G104), .C2(new_n192), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G101), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n196), .A2(new_n197), .B1(G101), .B2(new_n229), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n231), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n220), .A2(KEYINPUT2), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(new_n217), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n235), .B1(new_n240), .B2(new_n216), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n214), .A2(new_n215), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n217), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT67), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n234), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n227), .A2(new_n228), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G110), .B(G122), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n249), .B(KEYINPUT82), .Z(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n227), .A2(new_n250), .A3(new_n228), .A4(new_n247), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(KEYINPUT6), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT6), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n255), .A3(new_n251), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(new_n262), .ZN(new_n268));
  AND4_X1   g082(.A1(new_n266), .A2(new_n258), .A3(new_n260), .A4(new_n262), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n259), .A2(KEYINPUT1), .A3(G146), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n261), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(new_n258), .A3(new_n260), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n271), .B1(G125), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G224), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G953), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n254), .A2(new_n256), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n221), .A2(KEYINPUT83), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n221), .A2(KEYINPUT83), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n284), .A2(new_n218), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n223), .B1(new_n286), .B2(new_n216), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n207), .A2(new_n222), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n250), .B(KEYINPUT8), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n281), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n271), .A2(KEYINPUT84), .B1(KEYINPUT7), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n292), .A2(new_n279), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n279), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n290), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n295), .B2(new_n253), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n283), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n283), .B2(new_n296), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n270), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n277), .A2(KEYINPUT78), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n277), .A2(KEYINPUT78), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n275), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n223), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT10), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n234), .A2(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT11), .ZN(new_n308));
  INV_X1    g122(.A(G134), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(G137), .ZN(new_n310));
  INV_X1    g124(.A(G137), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT11), .A3(G134), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(G137), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT66), .A4(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n314), .A2(G131), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT66), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT65), .B(G131), .Z(new_n319));
  AND3_X1   g133(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n315), .A2(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n272), .B1(new_n267), .B2(G128), .ZN(new_n322));
  INV_X1    g136(.A(new_n277), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT68), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n261), .A2(new_n274), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n272), .A4(new_n277), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n324), .A2(KEYINPUT10), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n209), .A2(new_n328), .A3(new_n224), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n307), .A2(new_n321), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G110), .B(G140), .ZN(new_n331));
  INV_X1    g145(.A(G953), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n332), .A2(G227), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n322), .A2(new_n323), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n207), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT80), .B1(new_n223), .B2(new_n278), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n305), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n318), .A2(G131), .A3(new_n314), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n320), .A2(new_n319), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n340), .A2(KEYINPUT12), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT12), .B1(new_n340), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n330), .B(new_n335), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n307), .A2(new_n321), .A3(new_n329), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n321), .B1(new_n307), .B2(new_n329), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n334), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G469), .ZN(new_n351));
  INV_X1    g165(.A(G902), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n348), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n330), .A3(new_n335), .ZN(new_n357));
  INV_X1    g171(.A(new_n345), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n340), .A2(KEYINPUT12), .A3(new_n343), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n347), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(G469), .B(new_n357), .C1(new_n360), .C2(new_n335), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n353), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n363));
  INV_X1    g177(.A(G140), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT73), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n257), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT71), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n365), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n364), .A2(KEYINPUT71), .A3(G125), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(G146), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(KEYINPUT85), .A3(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n376), .A2(KEYINPUT85), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT18), .A2(G131), .ZN(new_n379));
  NOR2_X1   g193(.A1(G237), .A2(G953), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(G143), .A3(G214), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G143), .B1(new_n380), .B2(G214), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n259), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(KEYINPUT18), .A3(G131), .A4(new_n381), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n378), .A3(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(G113), .B(G122), .Z(new_n390));
  XOR2_X1   g204(.A(KEYINPUT86), .B(G104), .Z(new_n391));
  XOR2_X1   g205(.A(new_n390), .B(new_n391), .Z(new_n392));
  NAND3_X1  g206(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n375), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n365), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n257), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT72), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n398), .A3(new_n257), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n395), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G146), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n386), .A2(new_n381), .ZN(new_n403));
  INV_X1    g217(.A(new_n319), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n386), .A2(new_n319), .A3(new_n381), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n405), .B1(new_n408), .B2(KEYINPUT17), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n389), .B(new_n392), .C1(new_n402), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT19), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n370), .A2(new_n411), .A3(new_n371), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n374), .A2(KEYINPUT19), .A3(new_n375), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n257), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n401), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n389), .ZN(new_n416));
  INV_X1    g230(.A(new_n392), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT87), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n363), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  AOI211_X1 g237(.A(KEYINPUT20), .B(new_n421), .C1(new_n410), .C2(new_n418), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n389), .B1(new_n402), .B2(new_n409), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n417), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n426), .B2(new_n410), .ZN(new_n427));
  INV_X1    g241(.A(G475), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n423), .A2(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  INV_X1    g244(.A(G217), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n430), .A2(new_n431), .A3(G953), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n212), .A2(G122), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n192), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n192), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(KEYINPUT88), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT88), .ZN(new_n440));
  INV_X1    g254(.A(new_n438), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(new_n436), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G128), .B(G143), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n444), .A2(G134), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(G134), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n274), .A2(G143), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(G134), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n448), .A3(G134), .A4(new_n447), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n443), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n438), .A2(KEYINPUT89), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n434), .A2(new_n435), .A3(new_n454), .A4(new_n192), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n445), .A2(new_n453), .A3(new_n446), .A4(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n212), .A3(G122), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT90), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n192), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n435), .A2(KEYINPUT14), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n461), .A2(KEYINPUT90), .A3(new_n434), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT91), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(KEYINPUT91), .A3(new_n462), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n456), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n432), .B1(new_n452), .B2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n445), .A2(new_n446), .A3(new_n453), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n460), .A2(KEYINPUT91), .A3(new_n462), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT91), .B1(new_n460), .B2(new_n462), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n455), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n443), .A2(new_n450), .A3(new_n451), .ZN(new_n473));
  INV_X1    g287(.A(new_n432), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n468), .A2(KEYINPUT92), .A3(new_n352), .A4(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G478), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT15), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n476), .B(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n332), .A2(G952), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(G234), .B2(G237), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n352), .B(new_n332), .C1(G234), .C2(G237), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT21), .B(G898), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n429), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n362), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n300), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT70), .ZN(new_n489));
  NOR2_X1   g303(.A1(G472), .A2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT32), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n270), .B1(new_n342), .B2(new_n341), .ZN(new_n495));
  INV_X1    g309(.A(G131), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n311), .A2(G134), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(new_n313), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n320), .B2(new_n319), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n278), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n494), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n324), .A2(new_n499), .A3(new_n327), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(KEYINPUT30), .C1(new_n321), .C2(new_n270), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n246), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n503), .B(new_n245), .C1(new_n321), .C2(new_n270), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n380), .A2(G210), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT27), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT26), .B(G101), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT31), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n505), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n505), .B2(new_n511), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n506), .A2(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n343), .A2(new_n301), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n517), .A2(new_n518), .A3(new_n245), .A4(new_n503), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n246), .B1(new_n495), .B2(new_n501), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n510), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT69), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n525));
  NOR4_X1   g339(.A1(new_n522), .A2(new_n513), .A3(new_n514), .A4(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n493), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n503), .A2(KEYINPUT30), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n246), .B1(new_n528), .B2(new_n495), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT30), .B1(new_n517), .B2(new_n500), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n510), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n506), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n520), .A2(new_n535), .A3(new_n521), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n510), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n517), .A2(new_n503), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n246), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n520), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n536), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n527), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n506), .A2(new_n510), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT31), .B1(new_n531), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n505), .A2(new_n511), .A3(new_n512), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n525), .B1(new_n548), .B2(new_n522), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n523), .A2(KEYINPUT69), .A3(new_n546), .A4(new_n547), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT32), .B1(new_n551), .B2(new_n490), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n489), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n490), .B1(new_n524), .B2(new_n526), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n492), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n551), .A2(new_n493), .B1(G472), .B2(new_n542), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(KEYINPUT70), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n332), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n210), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n274), .A2(G119), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G110), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n210), .B2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n274), .A2(KEYINPUT23), .A3(G119), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(G110), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n402), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n564), .A2(new_n565), .ZN(new_n573));
  INV_X1    g387(.A(G110), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n569), .A3(new_n574), .A4(new_n562), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n372), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n257), .B1(new_n393), .B2(new_n395), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n561), .B1(new_n572), .B2(new_n580), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n560), .B(new_n579), .C1(new_n402), .C2(new_n571), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n431), .B1(G234), .B2(new_n352), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G902), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT74), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(KEYINPUT75), .ZN(new_n589));
  INV_X1    g403(.A(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n572), .A2(new_n580), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n560), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n572), .A2(new_n580), .A3(new_n561), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n352), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n583), .A2(KEYINPUT25), .A3(new_n352), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n488), .A2(new_n553), .A3(new_n557), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT93), .B(G101), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G3));
  NAND2_X1  g416(.A1(new_n551), .A2(new_n352), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT94), .A3(G472), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n549), .B2(new_n550), .ZN(new_n606));
  INV_X1    g420(.A(G472), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n610));
  AND4_X1   g424(.A1(new_n554), .A2(new_n599), .A3(new_n362), .A4(new_n486), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT96), .Z(new_n615));
  INV_X1    g429(.A(new_n300), .ZN(new_n616));
  INV_X1    g430(.A(new_n484), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n468), .A2(new_n352), .A3(new_n475), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n477), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n432), .A2(KEYINPUT98), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n452), .B2(new_n467), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n472), .B(new_n473), .C1(KEYINPUT98), .C2(new_n432), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(KEYINPUT33), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n468), .A2(new_n475), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n352), .A2(G478), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n620), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n429), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n618), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n615), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT100), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n429), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n479), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n618), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n615), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n572), .A2(new_n643), .A3(new_n580), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n643), .B1(new_n572), .B2(new_n580), .ZN(new_n646));
  OAI22_X1  g460(.A1(new_n645), .A2(new_n646), .B1(KEYINPUT36), .B2(new_n560), .ZN(new_n647));
  INV_X1    g461(.A(new_n646), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n560), .A2(KEYINPUT36), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n644), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n586), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT25), .B1(new_n583), .B2(new_n352), .ZN(new_n653));
  NOR4_X1   g467(.A1(new_n581), .A2(new_n582), .A3(new_n595), .A4(G902), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n584), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n300), .A2(new_n487), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n491), .B1(new_n549), .B2(new_n550), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n604), .B2(new_n608), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(new_n478), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n476), .B(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n481), .B1(new_n482), .B2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n429), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n362), .A2(new_n486), .A3(new_n670), .A4(new_n656), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n300), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n553), .A3(new_n557), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NOR2_X1   g488(.A1(new_n298), .A2(new_n299), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n669), .B(KEYINPUT39), .Z(new_n677));
  NAND3_X1  g491(.A1(new_n362), .A2(new_n486), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT40), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n429), .A2(new_n187), .A3(new_n479), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT104), .B1(new_n657), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n540), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n352), .B1(new_n683), .B2(new_n533), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n532), .B1(new_n505), .B2(new_n506), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n527), .B(new_n686), .C1(KEYINPUT32), .C2(new_n659), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n657), .A2(new_n681), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n676), .A2(new_n679), .A3(new_n682), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n259), .ZN(G45));
  INV_X1    g506(.A(new_n669), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n429), .A2(new_n629), .A3(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n362), .A2(new_n694), .A3(new_n486), .A4(new_n656), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n300), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n553), .A3(new_n557), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  NAND3_X1  g512(.A1(new_n553), .A2(new_n557), .A3(new_n599), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n700));
  AOI211_X1 g514(.A(G469), .B(G902), .C1(new_n346), .C2(new_n349), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n486), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT105), .ZN(new_n704));
  INV_X1    g518(.A(new_n486), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT105), .A4(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n699), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n632), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND2_X1  g526(.A1(new_n709), .A2(new_n639), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR3_X1   g528(.A1(new_n544), .A2(new_n552), .A3(new_n489), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT70), .B1(new_n555), .B2(new_n556), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n702), .B2(new_n486), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n300), .A3(new_n706), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n485), .A2(new_n656), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n717), .A2(new_n718), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n553), .A2(new_n557), .A3(new_n722), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n616), .A2(new_n704), .A3(new_n707), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  AOI21_X1  g542(.A(new_n510), .B1(new_n520), .B2(new_n540), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n490), .B1(new_n548), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT107), .B(G472), .Z(new_n731));
  OAI211_X1 g545(.A(new_n599), .B(new_n730), .C1(new_n606), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT108), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n720), .A2(new_n706), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n283), .A2(new_n296), .ZN(new_n735));
  INV_X1    g549(.A(new_n297), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n283), .A2(new_n296), .A3(new_n297), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n680), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n733), .A2(new_n617), .A3(new_n734), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  OAI211_X1 g555(.A(new_n656), .B(new_n730), .C1(new_n606), .C2(new_n731), .ZN(new_n742));
  INV_X1    g556(.A(new_n694), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n734), .A2(new_n744), .A3(new_n616), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  NAND2_X1  g560(.A1(new_n362), .A2(new_n486), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n187), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n298), .A2(new_n299), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n362), .A2(KEYINPUT109), .A3(new_n486), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n699), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n743), .A2(KEYINPUT42), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n737), .A2(new_n187), .A3(new_n738), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n748), .B2(new_n747), .ZN(new_n757));
  INV_X1    g571(.A(new_n599), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n555), .B2(new_n556), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n759), .A3(new_n694), .A4(new_n752), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n754), .A2(new_n755), .B1(new_n760), .B2(KEYINPUT42), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  INV_X1    g576(.A(new_n670), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n699), .A2(new_n763), .A3(new_n753), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n309), .ZN(G36));
  INV_X1    g579(.A(new_n629), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n429), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT43), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n656), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n660), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n756), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n357), .B1(new_n360), .B2(new_n335), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n351), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n354), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT46), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n701), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(KEYINPUT46), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n705), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n784), .A2(new_n785), .A3(new_n677), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n785), .B1(new_n784), .B2(new_n677), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n774), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  OR2_X1    g603(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n717), .A2(new_n599), .A3(new_n743), .A4(new_n756), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  XOR2_X1   g609(.A(new_n702), .B(KEYINPUT111), .Z(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT49), .Z(new_n797));
  INV_X1    g611(.A(new_n687), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n705), .A2(new_n750), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n599), .A2(new_n798), .A3(new_n767), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n676), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n802));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n792), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n796), .A2(new_n486), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n790), .A2(KEYINPUT115), .A3(new_n791), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n733), .A2(new_n481), .A3(new_n768), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(new_n751), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n676), .A2(new_n750), .A3(new_n734), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n808), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n708), .A2(new_n756), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n481), .A3(new_n768), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(new_n742), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n599), .A3(new_n481), .A4(new_n798), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n637), .A2(new_n766), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n802), .B1(new_n810), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n790), .A2(new_n791), .A3(new_n805), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n809), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n820), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(KEYINPUT117), .A3(new_n820), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n832), .A2(new_n817), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n832), .B2(new_n817), .ZN(new_n835));
  OAI211_X1 g649(.A(KEYINPUT51), .B(new_n827), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(G952), .B(new_n332), .C1(new_n821), .C2(new_n631), .ZN(new_n837));
  INV_X1    g651(.A(new_n759), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n819), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT48), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n837), .B(new_n840), .C1(new_n721), .C2(new_n808), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n825), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n717), .A2(new_n672), .B1(new_n721), .B2(new_n744), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n598), .A2(new_n651), .A3(new_n669), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n362), .A2(new_n845), .A3(new_n486), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n687), .A2(new_n846), .A3(new_n739), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n717), .B2(new_n696), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n687), .A2(new_n846), .A3(new_n739), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n745), .A2(new_n673), .A3(new_n697), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT112), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n600), .A2(new_n661), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n638), .A2(new_n630), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n618), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n614), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n429), .A2(new_n479), .A3(new_n669), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n362), .A2(new_n486), .A3(new_n656), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n756), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n553), .A3(new_n557), .ZN(new_n864));
  INV_X1    g678(.A(new_n744), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n864), .B1(new_n865), .B2(new_n753), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n764), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n860), .A2(new_n761), .A3(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n710), .A2(new_n727), .A3(new_n713), .A4(new_n740), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT52), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n856), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n860), .A2(new_n761), .A3(new_n867), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n727), .A2(new_n710), .A3(new_n713), .A4(new_n740), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n855), .B1(new_n844), .B2(new_n848), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n854), .B2(new_n855), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n843), .B1(new_n880), .B2(KEYINPUT54), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n843), .B(KEYINPUT54), .C1(new_n873), .C2(new_n879), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n871), .A2(new_n872), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT53), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n842), .A2(new_n881), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n801), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n332), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n352), .B1(new_n883), .B2(new_n885), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT56), .B1(new_n893), .B2(G210), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n254), .A2(new_n256), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n282), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT55), .Z(new_n897));
  OAI21_X1  g711(.A(new_n892), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n894), .B2(new_n897), .ZN(G51));
  INV_X1    g713(.A(new_n350), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT52), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT52), .B1(new_n850), .B2(new_n853), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT53), .B1(new_n903), .B2(new_n876), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT53), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n886), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n354), .B(KEYINPUT57), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g723(.A(G902), .B(new_n779), .C1(new_n904), .C2(new_n905), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n883), .A2(new_n885), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(KEYINPUT119), .A3(G902), .A4(new_n779), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n892), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT120), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n918), .B(new_n892), .C1(new_n909), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n410), .A3(new_n418), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .A4(new_n419), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n892), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n922), .A2(KEYINPUT121), .A3(new_n892), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(G60));
  INV_X1    g742(.A(new_n907), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n624), .A2(new_n626), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n892), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n881), .B2(new_n887), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n627), .ZN(G63));
  NAND2_X1  g750(.A1(new_n647), .A2(new_n650), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n913), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n913), .A2(new_n939), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n892), .B(new_n940), .C1(new_n941), .C2(new_n583), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G66));
  INV_X1    g758(.A(new_n483), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n332), .B1(new_n945), .B2(G224), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n869), .A2(new_n860), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT123), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(new_n332), .ZN(new_n949));
  INV_X1    g763(.A(G898), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n895), .B1(new_n950), .B2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n949), .B(new_n951), .ZN(G69));
  NAND2_X1  g766(.A1(G227), .A2(G900), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n739), .B(new_n759), .C1(new_n786), .C2(new_n787), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n844), .A2(new_n697), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n764), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n761), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n794), .A2(new_n954), .A3(new_n957), .A4(new_n788), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n332), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n668), .A2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT124), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n502), .A2(new_n504), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n412), .A2(new_n413), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n963), .B(new_n964), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(G953), .B(new_n953), .C1(new_n962), .C2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n953), .A2(G953), .ZN(new_n971));
  INV_X1    g785(.A(new_n699), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n756), .A2(new_n678), .A3(new_n858), .ZN(new_n973));
  AOI22_X1  g787(.A1(new_n792), .A2(new_n793), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n955), .A2(new_n691), .A3(KEYINPUT62), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT62), .B1(new_n955), .B2(new_n691), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n974), .A2(new_n788), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n966), .B1(new_n978), .B2(G953), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n970), .A2(new_n971), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n967), .A2(new_n980), .ZN(G72));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n607), .A2(new_n352), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT126), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n948), .B2(new_n977), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n685), .B1(new_n986), .B2(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(KEYINPUT127), .B2(new_n986), .ZN(new_n988));
  INV_X1    g802(.A(new_n984), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n534), .A2(new_n685), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n891), .B1(new_n880), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n985), .B1(new_n948), .B2(new_n958), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n534), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n988), .A2(new_n994), .ZN(G57));
endmodule


