//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT2), .A2(G113), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT2), .A2(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT71), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT2), .A3(G113), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G119), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G146), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(new_n199), .ZN(new_n202));
  NAND3_X1  g016(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT0), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT64), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n198), .B1(new_n202), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n200), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n211), .B1(new_n216), .B2(G143), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(KEYINPUT0), .B2(G128), .ZN(new_n219));
  INV_X1    g033(.A(new_n208), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n203), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n212), .A2(G143), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n216), .B2(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n220), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n210), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT68), .A2(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n231), .A2(KEYINPUT68), .A3(KEYINPUT11), .A4(G134), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(G137), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n232), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT69), .B(G131), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n233), .A2(new_n234), .B1(new_n229), .B2(G137), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n230), .A4(new_n232), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n210), .A2(new_n222), .A3(new_n225), .A4(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n227), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n236), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n229), .A2(G137), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n199), .B1(new_n213), .B2(new_n215), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n217), .B1(new_n254), .B2(new_n206), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n224), .A2(new_n253), .A3(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n197), .B1(new_n245), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n249), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT1), .B1(new_n201), .B2(new_n199), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n202), .B1(G128), .B2(new_n261), .ZN(new_n262));
  NOR4_X1   g076(.A1(new_n252), .A2(KEYINPUT1), .A3(new_n206), .A4(new_n223), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n242), .A2(new_n210), .A3(new_n222), .A4(new_n225), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n197), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n259), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(G237), .A2(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G210), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n188), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n267), .ZN(new_n277));
  INV_X1    g091(.A(new_n269), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n245), .A2(new_n258), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n197), .ZN(new_n280));
  INV_X1    g094(.A(new_n275), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  INV_X1    g098(.A(new_n266), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT30), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n245), .A2(new_n286), .A3(new_n258), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n264), .A2(new_n265), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT30), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n285), .B1(new_n290), .B2(new_n196), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n284), .B1(new_n291), .B2(new_n275), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n197), .B1(new_n287), .B2(new_n289), .ZN(new_n293));
  NOR4_X1   g107(.A1(new_n293), .A2(KEYINPUT31), .A3(new_n285), .A4(new_n281), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n283), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n187), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n275), .A2(KEYINPUT29), .ZN(new_n299));
  AND4_X1   g113(.A1(new_n242), .A2(new_n210), .A3(new_n222), .A4(new_n225), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n196), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n197), .B1(new_n264), .B2(new_n265), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT74), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n266), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT73), .A4(new_n197), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n304), .A2(new_n306), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n268), .B(new_n299), .C1(new_n310), .C2(KEYINPUT28), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT75), .B1(new_n311), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n293), .A2(new_n285), .A3(new_n275), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n270), .A2(new_n281), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(KEYINPUT28), .ZN(new_n317));
  INV_X1    g131(.A(new_n299), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n277), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n312), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G472), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n291), .A2(new_n275), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT31), .ZN(new_n326));
  INV_X1    g140(.A(new_n294), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n276), .A4(new_n282), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n298), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n206), .A2(G119), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G128), .ZN(new_n335));
  MUX2_X1   g149(.A(new_n333), .B(new_n332), .S(new_n335), .Z(new_n336));
  INV_X1    g150(.A(G110), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n331), .A2(new_n335), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT24), .B(G110), .Z(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n342), .B1(new_n348), .B2(new_n216), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n347), .A2(new_n201), .A3(KEYINPUT78), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT16), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n345), .A2(G140), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n343), .B2(G125), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n345), .A2(KEYINPUT76), .A3(G140), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT77), .A3(G146), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT77), .B1(new_n359), .B2(G146), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n341), .B(new_n351), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(G146), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n212), .B(new_n353), .C1(new_n358), .C2(new_n352), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n339), .ZN(new_n367));
  INV_X1    g181(.A(new_n340), .ZN(new_n368));
  OAI221_X1 g182(.A(new_n366), .B1(new_n337), .B2(new_n336), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G953), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(G221), .A3(G234), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT79), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G137), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n363), .A2(new_n369), .A3(new_n375), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n321), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(KEYINPUT25), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(G234), .B2(new_n321), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n380), .A2(KEYINPUT25), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n377), .A2(new_n378), .A3(new_n321), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n383), .A2(G902), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(KEYINPUT81), .Z(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n377), .A2(new_n378), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT82), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n330), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n239), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n271), .A2(G143), .A3(G214), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(G143), .B1(new_n271), .B2(G214), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G237), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n371), .A3(G214), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n199), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n239), .A3(new_n401), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n344), .A2(new_n346), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n216), .B(new_n411), .C1(new_n358), .C2(new_n410), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT77), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n364), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n415), .B2(new_n360), .ZN(new_n416));
  OAI22_X1  g230(.A1(new_n349), .A2(new_n350), .B1(new_n212), .B2(new_n358), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n407), .A2(new_n401), .ZN(new_n418));
  AND2_X1   g232(.A1(KEYINPUT18), .A2(G131), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n399), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n404), .A2(new_n425), .A3(new_n408), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(KEYINPUT17), .A3(new_n400), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n364), .A2(new_n426), .A3(new_n365), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(new_n428), .A3(new_n398), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n395), .B(KEYINPUT20), .C1(new_n423), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(G475), .A2(G902), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n409), .B(new_n412), .C1(new_n361), .C2(new_n362), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n398), .B1(new_n432), .B2(new_n424), .ZN(new_n433));
  INV_X1    g247(.A(new_n429), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n423), .A2(new_n429), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT20), .A3(new_n431), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n430), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n398), .B1(new_n424), .B2(new_n428), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n321), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G475), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(KEYINPUT91), .A3(new_n436), .ZN(new_n444));
  INV_X1    g258(.A(new_n431), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n394), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G214), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT3), .B1(new_n397), .B2(G107), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n451));
  INV_X1    g265(.A(G107), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(G104), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n397), .A2(G107), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G101), .ZN(new_n456));
  INV_X1    g270(.A(G101), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n450), .A2(new_n453), .A3(new_n457), .A4(new_n454), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(KEYINPUT4), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n460), .A3(G101), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n196), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n194), .A2(new_n195), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT5), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n334), .A3(G116), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(G113), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n397), .A2(G107), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n452), .A2(G104), .ZN(new_n469));
  OAI21_X1  g283(.A(G101), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n458), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n458), .B2(new_n470), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n463), .B(new_n467), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n462), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(G110), .A2(G122), .ZN(new_n476));
  NAND2_X1  g290(.A1(G110), .A2(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT87), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n462), .A2(new_n474), .A3(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n345), .B1(new_n262), .B2(new_n263), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n210), .A2(new_n222), .A3(new_n225), .A4(G125), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G224), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G953), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n491), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n475), .A2(new_n496), .A3(new_n483), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n486), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n458), .A2(new_n470), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n467), .A2(new_n463), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT88), .B(KEYINPUT8), .Z(new_n503));
  AND3_X1   g317(.A1(new_n479), .A2(new_n481), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n479), .B2(new_n481), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n467), .B(new_n463), .C1(new_n499), .C2(KEYINPUT89), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT90), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n492), .A2(KEYINPUT7), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n487), .A2(new_n513), .A3(new_n488), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n489), .A2(KEYINPUT7), .A3(new_n492), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n512), .A2(new_n514), .A3(new_n485), .A4(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n498), .A2(new_n516), .A3(new_n321), .ZN(new_n517));
  OAI21_X1  g331(.A(G210), .B1(G237), .B2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n498), .A2(new_n516), .A3(new_n321), .A4(new_n518), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n449), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT20), .B1(new_n438), .B2(new_n431), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n436), .B(new_n445), .C1(new_n423), .C2(new_n429), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n444), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n430), .A2(new_n431), .B1(G475), .B2(new_n442), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT92), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n371), .A2(G952), .ZN(new_n528));
  NAND2_X1  g342(.A1(G234), .A2(G237), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT95), .Z(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT21), .B(G898), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(G902), .A3(G953), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n447), .A2(new_n522), .A3(new_n527), .A4(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G469), .ZN(new_n536));
  OAI21_X1  g350(.A(G128), .B1(new_n200), .B2(new_n253), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n252), .B2(new_n223), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT83), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(KEYINPUT83), .C1(new_n252), .C2(new_n223), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n256), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n499), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT10), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n459), .A2(new_n461), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n226), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n257), .B(KEYINPUT10), .C1(new_n473), .C2(new_n472), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n242), .B(KEYINPUT85), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n546), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT86), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(KEYINPUT86), .A2(KEYINPUT12), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n262), .A2(new_n543), .A3(new_n263), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n543), .B2(new_n542), .ZN(new_n557));
  INV_X1    g371(.A(new_n242), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n554), .B(new_n555), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G140), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n371), .A2(G227), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n560), .B(new_n561), .Z(new_n562));
  OAI21_X1  g376(.A(new_n544), .B1(new_n257), .B2(new_n543), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(new_n552), .A3(new_n553), .A4(new_n242), .ZN(new_n564));
  AND4_X1   g378(.A1(new_n551), .A2(new_n559), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n242), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n567), .B2(new_n551), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n536), .B(new_n321), .C1(new_n565), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(G469), .A2(G902), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n559), .A2(new_n551), .A3(new_n564), .ZN(new_n571));
  INV_X1    g385(.A(new_n562), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n551), .A2(new_n562), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n567), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(G469), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n570), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT9), .B(G234), .Z(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G221), .B1(new_n579), .B2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT94), .ZN(new_n582));
  XNOR2_X1  g396(.A(G116), .B(G122), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT93), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n452), .ZN(new_n585));
  XNOR2_X1  g399(.A(G128), .B(G143), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n229), .ZN(new_n587));
  INV_X1    g401(.A(G116), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(KEYINPUT14), .A3(G122), .ZN(new_n589));
  INV_X1    g403(.A(new_n583), .ZN(new_n590));
  OAI211_X1 g404(.A(G107), .B(new_n589), .C1(new_n590), .C2(KEYINPUT14), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n585), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n229), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n586), .A2(KEYINPUT13), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n199), .A2(G128), .ZN(new_n596));
  OAI21_X1  g410(.A(G134), .B1(new_n596), .B2(KEYINPUT13), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n594), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n583), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G107), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n598), .B1(new_n601), .B2(new_n585), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n579), .A2(new_n382), .A3(G953), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OR3_X1    g418(.A1(new_n593), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n593), .B2(new_n602), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G478), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(KEYINPUT15), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n321), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n607), .B2(new_n321), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n582), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(KEYINPUT94), .A3(new_n611), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n535), .A2(new_n581), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n393), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n328), .B2(new_n321), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n295), .A2(new_n297), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n581), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n392), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n522), .A2(new_n534), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n605), .A2(KEYINPUT33), .A3(new_n606), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT33), .B1(new_n605), .B2(new_n606), .ZN(new_n629));
  OAI21_X1  g443(.A(G478), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n607), .A2(new_n608), .A3(new_n321), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n608), .A2(new_n321), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n440), .A2(new_n446), .A3(new_n394), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT92), .B1(new_n525), .B2(new_n526), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n626), .A2(new_n627), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT34), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  XOR2_X1   g455(.A(new_n534), .B(KEYINPUT96), .Z(new_n642));
  NAND2_X1  g456(.A1(new_n522), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n523), .A2(new_n524), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n614), .A2(new_n616), .A3(new_n443), .A4(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n626), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT35), .B(G107), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n370), .A2(KEYINPUT97), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n376), .A2(KEYINPUT36), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n363), .A2(new_n369), .A3(new_n651), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n650), .B1(new_n649), .B2(new_n652), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n389), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n386), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n618), .A2(new_n624), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n529), .A2(new_n660), .A3(G902), .A4(G953), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n531), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT99), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n645), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n577), .A2(new_n580), .A3(new_n522), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n330), .A2(new_n665), .A3(new_n656), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XOR2_X1   g482(.A(new_n664), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n625), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT40), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n447), .A2(new_n527), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(new_n617), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n291), .A2(new_n281), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n321), .B1(new_n310), .B2(new_n275), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n298), .A2(new_n329), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n298), .A2(KEYINPUT101), .A3(new_n329), .A4(new_n676), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n520), .A2(new_n521), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  OR3_X1    g498(.A1(new_n684), .A2(new_n449), .A3(new_n656), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n671), .A2(new_n673), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  AOI211_X1 g502(.A(new_n664), .B(new_n634), .C1(new_n447), .C2(new_n527), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n330), .A2(new_n656), .A3(new_n666), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  AND2_X1   g505(.A1(new_n559), .A2(new_n564), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n567), .A2(new_n551), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n692), .A2(new_n574), .B1(new_n693), .B2(new_n572), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n694), .B2(G902), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n580), .A3(new_n569), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n638), .A2(new_n696), .A3(new_n627), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n330), .A2(new_n697), .A3(new_n392), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n695), .A2(new_n522), .A3(new_n580), .A4(new_n569), .ZN(new_n701));
  INV_X1    g515(.A(new_n642), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n701), .A2(new_n702), .A3(new_n645), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n330), .A2(new_n392), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  NOR3_X1   g519(.A1(new_n535), .A2(new_n696), .A3(new_n617), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n330), .A2(new_n656), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  XOR2_X1   g522(.A(new_n296), .B(KEYINPUT102), .Z(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n305), .B(new_n303), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n308), .A2(new_n309), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n267), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n711), .B1(new_n714), .B2(new_n268), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n317), .A2(KEYINPUT103), .A3(new_n277), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n281), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n292), .A2(new_n294), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n710), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n328), .A2(new_n321), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT104), .B(G472), .Z(new_n721));
  AOI21_X1  g535(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n701), .A2(new_n702), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n386), .A2(new_n391), .A3(KEYINPUT105), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT105), .B1(new_n386), .B2(new_n391), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n673), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  INV_X1    g542(.A(new_n721), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n328), .B2(new_n321), .ZN(new_n730));
  INV_X1    g544(.A(new_n656), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n730), .A2(new_n719), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n701), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n689), .A3(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT106), .B(G125), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G27));
  NAND2_X1  g550(.A1(new_n330), .A2(new_n726), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n682), .A2(new_n449), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n577), .A3(new_n580), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(new_n689), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n330), .A3(new_n392), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n738), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NAND3_X1  g561(.A1(new_n393), .A2(new_n665), .A3(new_n741), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  INV_X1    g563(.A(new_n672), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n635), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n672), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n755), .A2(KEYINPUT43), .A3(new_n635), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n751), .A2(new_n759), .A3(new_n752), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n754), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n624), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(KEYINPUT44), .A3(new_n762), .A4(new_n656), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n764), .A3(new_n740), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n763), .B2(new_n740), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n762), .A3(new_n656), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n573), .A2(new_n575), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT45), .ZN(new_n773));
  OAI21_X1  g587(.A(G469), .B1(new_n773), .B2(G902), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n569), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n580), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n669), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n689), .A3(new_n740), .A4(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n330), .A3(new_n392), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n343), .ZN(G42));
  NAND2_X1  g602(.A1(new_n695), .A2(new_n569), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT49), .Z(new_n790));
  AND4_X1   g604(.A1(new_n580), .A2(new_n790), .A3(new_n684), .A4(new_n726), .ZN(new_n791));
  INV_X1    g605(.A(new_n681), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n755), .A2(new_n635), .A3(new_n757), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n448), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n612), .A2(new_n613), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n672), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n643), .B1(new_n797), .B2(new_n638), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n624), .A3(new_n392), .A4(new_n625), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n619), .A2(new_n657), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n698), .A2(new_n707), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n704), .A2(new_n727), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT110), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n698), .A2(new_n704), .A3(new_n707), .A4(new_n727), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n800), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n742), .A2(KEYINPUT111), .A3(new_n732), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT111), .B1(new_n742), .B2(new_n732), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n664), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n796), .A2(new_n443), .A3(new_n644), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n330), .A2(new_n812), .A3(new_n656), .A4(new_n741), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n746), .A2(new_n810), .A3(new_n748), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n795), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n739), .A2(new_n742), .B1(new_n744), .B2(new_n738), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n813), .B1(new_n808), .B2(new_n809), .ZN(new_n817));
  INV_X1    g631(.A(new_n748), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n804), .B(new_n805), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT112), .A4(new_n800), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n734), .A2(new_n667), .A3(new_n690), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n656), .A2(new_n664), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n681), .A2(new_n666), .A3(new_n673), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n823), .A2(new_n825), .A3(new_n822), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n823), .A2(new_n825), .A3(new_n822), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT52), .B1(new_n831), .B2(new_n826), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n815), .A2(new_n821), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n828), .B1(new_n823), .B2(new_n825), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n831), .A2(new_n826), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n835), .B1(new_n836), .B2(new_n828), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n815), .A4(new_n821), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n833), .A2(new_n838), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n804), .A2(new_n838), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n837), .A2(new_n800), .A3(new_n819), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n834), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n839), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT115), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n842), .A2(new_n851), .A3(new_n847), .A4(new_n848), .ZN(new_n852));
  INV_X1    g666(.A(new_n531), .ZN(new_n853));
  INV_X1    g667(.A(new_n740), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n696), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n792), .A2(new_n392), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(new_n672), .A3(new_n635), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n789), .A2(new_n580), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n784), .B2(new_n785), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n854), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n761), .A2(new_n853), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n722), .A2(new_n726), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n857), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n684), .A3(new_n862), .ZN(new_n865));
  NAND2_X1  g679(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n866));
  INV_X1    g680(.A(new_n696), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n867), .B(new_n449), .C1(KEYINPUT116), .C2(KEYINPUT50), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n866), .B1(new_n865), .B2(new_n868), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n861), .A2(KEYINPUT117), .A3(new_n855), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT117), .B1(new_n861), .B2(new_n855), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n732), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n864), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n871), .A2(new_n864), .A3(KEYINPUT51), .A4(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n863), .A2(new_n733), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n528), .A4(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n330), .B(new_n726), .C1(new_n872), .C2(new_n873), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT48), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n856), .A2(new_n638), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n850), .A2(new_n852), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n794), .B1(new_n885), .B2(new_n886), .ZN(G75));
  AOI21_X1  g701(.A(new_n321), .B1(new_n843), .B2(new_n846), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(G210), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT56), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n486), .A2(new_n497), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(new_n495), .Z(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n889), .B2(new_n890), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n371), .A2(G952), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G51));
  NAND2_X1  g711(.A1(new_n843), .A2(new_n846), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n847), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n570), .B(KEYINPUT57), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT118), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT118), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n694), .B(KEYINPUT119), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n888), .A2(G469), .A3(new_n773), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n896), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(new_n438), .Z(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n896), .ZN(G60));
  NOR2_X1   g727(.A1(new_n628), .A2(new_n629), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n632), .B(KEYINPUT59), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n900), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n896), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n850), .A2(new_n852), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n915), .ZN(new_n920));
  INV_X1    g734(.A(new_n914), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n843), .B2(new_n846), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n653), .B2(new_n654), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n377), .A2(new_n378), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n926), .B(new_n917), .C1(new_n927), .C2(new_n925), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g743(.A(G953), .B1(new_n532), .B2(new_n490), .ZN(new_n930));
  INV_X1    g744(.A(new_n807), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(G953), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  INV_X1    g747(.A(G898), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n891), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  NAND2_X1  g750(.A1(new_n687), .A2(new_n823), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n787), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n687), .A2(new_n823), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n797), .A2(new_n638), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n393), .A2(new_n669), .A3(new_n741), .A4(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(new_n781), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n371), .ZN(new_n945));
  MUX2_X1   g759(.A(new_n347), .B(new_n358), .S(KEYINPUT19), .Z(new_n946));
  XOR2_X1   g760(.A(new_n290), .B(new_n946), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n371), .B1(G227), .B2(G900), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n660), .A2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT122), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n673), .A2(new_n522), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n737), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n780), .B1(new_n771), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n746), .A2(new_n748), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n787), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n957), .A3(new_n823), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n952), .B1(new_n958), .B2(new_n371), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n948), .B(new_n950), .C1(new_n947), .C2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT123), .B1(new_n959), .B2(new_n947), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  INV_X1    g776(.A(new_n947), .ZN(new_n963));
  INV_X1    g777(.A(new_n823), .ZN(new_n964));
  INV_X1    g778(.A(new_n954), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n763), .A2(new_n740), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n765), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n965), .B1(new_n968), .B2(new_n770), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(new_n969), .B2(new_n780), .ZN(new_n970));
  AOI21_X1  g784(.A(G953), .B1(new_n970), .B2(new_n957), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n962), .B(new_n963), .C1(new_n971), .C2(new_n952), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n961), .A2(new_n972), .A3(new_n948), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n973), .A2(KEYINPUT124), .A3(new_n949), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT124), .B1(new_n973), .B2(new_n949), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n960), .B1(new_n974), .B2(new_n975), .ZN(G72));
  XNOR2_X1  g790(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n621), .A2(new_n321), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n977), .B(new_n978), .Z(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n958), .B2(new_n807), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n314), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n980), .B1(new_n944), .B2(new_n807), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n896), .B1(new_n984), .B2(new_n674), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n674), .A2(new_n314), .A3(new_n979), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT127), .Z(new_n987));
  NAND3_X1  g801(.A1(new_n834), .A2(new_n839), .A3(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(G57));
endmodule


