//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT64), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n202), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n252), .A2(new_n213), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G1), .B2(new_n207), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n254), .B2(new_n202), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT65), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(new_n207), .A3(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n252), .A2(new_n213), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n255), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G169), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1698), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G222), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT3), .B(G33), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(G1698), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n271), .B1(new_n272), .B2(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n278), .A3(G274), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n285), .B1(G226), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n264), .B1(new_n265), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n280), .A2(new_n292), .A3(new_n289), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(G200), .ZN(new_n295));
  XOR2_X1   g0095(.A(new_n295), .B(KEYINPUT66), .Z(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n264), .A2(KEYINPUT9), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(KEYINPUT9), .B2(new_n264), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n298), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n295), .B(KEYINPUT66), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT10), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n294), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n284), .B1(new_n220), .B2(new_n287), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT67), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n284), .B(KEYINPUT67), .C1(new_n220), .C2(new_n287), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G97), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n226), .A2(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(G226), .B2(G1698), .ZN(new_n313));
  AND2_X1   g0113(.A1(KEYINPUT3), .A2(G33), .ZN(new_n314));
  NOR2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n311), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n309), .A2(new_n310), .B1(new_n317), .B2(new_n279), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n319));
  XNOR2_X1  g0119(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G200), .ZN(new_n321));
  INV_X1    g0121(.A(new_n260), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n322), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n207), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n272), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n263), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT11), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT12), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n250), .B2(new_n219), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n249), .A2(KEYINPUT12), .A3(G68), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n254), .A2(new_n219), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n318), .A2(new_n319), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n335), .B(G190), .C1(new_n336), .C2(new_n318), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n321), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n335), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n318), .A2(new_n319), .ZN(new_n340));
  OAI21_X1  g0140(.A(G169), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n335), .B(G179), .C1(new_n336), .C2(new_n318), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n320), .A2(new_n344), .A3(G169), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n334), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n338), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n288), .A2(G244), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n270), .A2(G232), .ZN(new_n350));
  INV_X1    g0150(.A(G107), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n350), .B1(new_n351), .B2(new_n273), .C1(new_n220), .C2(new_n275), .ZN(new_n352));
  AOI211_X1 g0152(.A(new_n285), .B(new_n349), .C1(new_n352), .C2(new_n279), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G20), .A2(G77), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n356), .B1(new_n256), .B2(new_n322), .C1(new_n324), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n263), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n250), .A2(new_n272), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n272), .C2(new_n254), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n353), .B2(G190), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n353), .A2(new_n292), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n361), .B1(new_n353), .B2(G169), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n306), .A2(new_n348), .A3(new_n363), .A4(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n284), .B1(new_n226), .B2(new_n287), .ZN(new_n370));
  INV_X1    g0170(.A(G1698), .ZN(new_n371));
  OAI211_X1 g0171(.A(G223), .B(new_n371), .C1(new_n314), .C2(new_n315), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT71), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n273), .A2(new_n374), .A3(G223), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n273), .A2(G226), .A3(G1698), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n370), .B1(new_n378), .B2(new_n279), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n265), .ZN(new_n380));
  AOI211_X1 g0180(.A(new_n292), .B(new_n370), .C1(new_n378), .C2(new_n279), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n369), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n258), .A2(new_n254), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n250), .B2(new_n258), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n225), .A2(new_n219), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n201), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n260), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NOR4_X1   g0191(.A1(new_n314), .A2(new_n315), .A3(new_n391), .A4(G20), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT69), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n314), .B2(new_n315), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n268), .A2(KEYINPUT69), .A3(new_n269), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(new_n207), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n396), .B2(new_n391), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n390), .B1(new_n397), .B2(new_n219), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n263), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n391), .B1(new_n273), .B2(G20), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT70), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT70), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n316), .A2(new_n403), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(G68), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n388), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT16), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n384), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n378), .A2(new_n279), .ZN(new_n409));
  INV_X1    g0209(.A(new_n370), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(G179), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(KEYINPUT72), .C1(new_n265), .C2(new_n379), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n382), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n354), .B1(new_n409), .B2(new_n410), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n299), .B(new_n370), .C1(new_n378), .C2(new_n279), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n409), .A2(G190), .A3(new_n410), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(KEYINPUT73), .C1(new_n354), .C2(new_n379), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n384), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n396), .A2(new_n391), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n401), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G68), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n253), .B1(new_n426), .B2(new_n390), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n405), .A2(new_n406), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n389), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n423), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n408), .B1(new_n419), .B2(new_n421), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT17), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n415), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  OR3_X1    g0236(.A1(new_n368), .A2(KEYINPUT74), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT74), .B1(new_n368), .B2(new_n436), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OR3_X1    g0239(.A1(new_n249), .A2(KEYINPUT25), .A3(G107), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT25), .B1(new_n249), .B2(G107), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n206), .A2(G33), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n249), .A2(new_n442), .A3(new_n213), .A4(new_n252), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n440), .B(new_n441), .C1(new_n351), .C2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT76), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n273), .A2(new_n207), .A3(G87), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT22), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT22), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n273), .A2(new_n448), .A3(new_n207), .A4(G87), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G116), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G20), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT23), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n207), .B2(G107), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n351), .A2(KEYINPUT23), .A3(G20), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT24), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n456), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n447), .B2(new_n449), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n263), .B1(new_n461), .B2(KEYINPUT24), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n445), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n282), .A2(G1), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n278), .A2(G274), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n279), .B1(new_n465), .B2(new_n464), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(G264), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n273), .A2(G257), .ZN(new_n471));
  INV_X1    g0271(.A(G294), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n471), .A2(new_n371), .B1(new_n267), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT77), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n270), .A2(new_n474), .A3(G250), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n273), .A2(new_n371), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT77), .B1(new_n476), .B2(new_n222), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n470), .B1(new_n478), .B2(new_n278), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n265), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n470), .B(new_n292), .C1(new_n478), .C2(new_n278), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n463), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n477), .A2(new_n475), .ZN(new_n483));
  INV_X1    g0283(.A(new_n473), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n278), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n470), .ZN(new_n486));
  OAI21_X1  g0286(.A(G200), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n457), .A2(new_n458), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n263), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n470), .B(G190), .C1(new_n478), .C2(new_n278), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n487), .A2(new_n490), .A3(new_n445), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n482), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n482), .A2(new_n492), .A3(KEYINPUT78), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n468), .B1(G270), .B2(new_n469), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n273), .A2(G264), .A3(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n316), .A2(G303), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n471), .C2(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n279), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n498), .A2(new_n502), .A3(G179), .ZN(new_n503));
  INV_X1    g0303(.A(new_n443), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G116), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n250), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(new_n207), .C1(G33), .C2(new_n227), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n509), .B(new_n263), .C1(new_n207), .C2(G116), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT20), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n505), .B(new_n507), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n503), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n498), .A2(new_n502), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(new_n514), .A3(KEYINPUT21), .A4(G169), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n514), .A3(G169), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n514), .B1(new_n516), .B2(G200), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n299), .B2(new_n516), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n518), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G244), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n525));
  OAI211_X1 g0325(.A(G238), .B(new_n371), .C1(new_n314), .C2(new_n315), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(new_n451), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n279), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n278), .A2(G274), .A3(new_n465), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n206), .A2(G45), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n278), .A2(G250), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n265), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n279), .B2(new_n527), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n292), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n207), .B1(new_n311), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n221), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n207), .B(G68), .C1(new_n314), .C2(new_n315), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n538), .B1(new_n324), .B2(new_n227), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n263), .B1(new_n250), .B2(new_n357), .ZN(new_n546));
  INV_X1    g0346(.A(new_n357), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n504), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n535), .A2(new_n537), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n536), .A2(new_n354), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n249), .A2(new_n442), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT75), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(G87), .A4(new_n253), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT75), .B1(new_n443), .B2(new_n221), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n546), .B(new_n556), .C1(new_n534), .C2(new_n299), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n550), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n402), .A2(G107), .A3(new_n404), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n351), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n227), .A2(new_n351), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(new_n540), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n563), .B2(KEYINPUT6), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n253), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n250), .A2(new_n227), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n443), .B2(new_n227), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G250), .B(G1698), .C1(new_n314), .C2(new_n315), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(new_n371), .C1(new_n314), .C2(new_n315), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n508), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT4), .B1(new_n270), .B2(G244), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n279), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n468), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n469), .A2(G257), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n578), .A2(new_n354), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(G190), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n569), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n265), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n575), .A2(new_n292), .A3(new_n577), .A4(new_n576), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n566), .C2(new_n568), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n559), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n524), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n439), .A2(new_n497), .A3(new_n586), .ZN(G372));
  OAI21_X1  g0387(.A(new_n411), .B1(new_n265), .B2(new_n379), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n408), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT18), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n338), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n366), .B1(new_n347), .B2(new_n346), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n433), .A2(new_n435), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n302), .A2(new_n305), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n294), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n439), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n532), .A2(KEYINPUT80), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT80), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n529), .A2(new_n531), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT79), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n527), .A2(new_n604), .A3(new_n279), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n265), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n537), .A2(new_n549), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(G200), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n528), .A2(new_n533), .A3(G190), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n546), .A2(new_n556), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n608), .A2(new_n607), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n583), .B1(new_n566), .B2(new_n568), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n578), .A2(new_n265), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT26), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g0418(.A(KEYINPUT82), .B(KEYINPUT26), .Z(new_n619));
  NOR3_X1   g0419(.A1(new_n584), .A2(new_n558), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n609), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(KEYINPUT83), .B(new_n609), .C1(new_n618), .C2(new_n620), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n518), .A2(new_n482), .A3(new_n521), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n614), .A2(new_n581), .A3(new_n492), .A4(new_n584), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT81), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n623), .A2(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n597), .B1(new_n598), .B2(new_n630), .ZN(G369));
  NAND3_X1  g0431(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n514), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT84), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n524), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n518), .A2(new_n521), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n639), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G330), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n637), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n482), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n463), .A2(new_n637), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n497), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n641), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n637), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n497), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n637), .B(KEYINPUT85), .Z(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n482), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n210), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n540), .A2(new_n221), .A3(new_n506), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n666), .B(KEYINPUT86), .Z(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n217), .B2(new_n665), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT31), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n485), .A2(new_n486), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n575), .A2(new_n577), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n673), .A2(new_n503), .A3(new_n675), .A4(new_n536), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT87), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(G179), .B1(new_n498), .B2(new_n502), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n479), .A2(new_n681), .A3(new_n578), .A4(new_n606), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n676), .B2(new_n678), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n677), .B1(new_n676), .B2(new_n678), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n672), .B1(new_n685), .B2(new_n648), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n497), .A2(new_n586), .A3(new_n658), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n470), .B(new_n536), .C1(new_n478), .C2(new_n278), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n498), .A2(new_n502), .A3(G179), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n688), .A2(new_n689), .A3(new_n674), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(KEYINPUT30), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT31), .B(new_n659), .C1(new_n683), .C2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n686), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n623), .A2(new_n624), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n628), .A2(new_n629), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n659), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT88), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT88), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n630), .B2(new_n659), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n625), .A2(new_n626), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n608), .B2(new_n607), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n614), .A2(new_n617), .A3(KEYINPUT26), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n619), .B1(new_n584), .B2(new_n558), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n637), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n695), .B1(new_n703), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n671), .B1(new_n711), .B2(G1), .ZN(G364));
  AND2_X1   g0512(.A1(new_n207), .A2(G13), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n206), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n664), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n644), .A2(new_n645), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n647), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n213), .B1(G20), .B2(new_n265), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n210), .A2(new_n273), .ZN(new_n725));
  INV_X1    g0525(.A(G355), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n725), .A2(new_n726), .B1(G116), .B2(new_n210), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT89), .Z(new_n728));
  NAND2_X1  g0528(.A1(new_n394), .A2(new_n395), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n663), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G45), .B2(new_n217), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(G45), .B2(new_n247), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n724), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n716), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n207), .A2(new_n292), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G190), .A3(G200), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(KEYINPUT91), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(KEYINPUT91), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G326), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n207), .A2(new_n299), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n292), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n207), .A2(G190), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G322), .A2(new_n745), .B1(new_n749), .B2(G329), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n354), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n743), .A2(new_n746), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G303), .A2(new_n753), .B1(new_n755), .B2(G311), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n207), .B1(new_n747), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n746), .A2(new_n751), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n316), .B1(new_n757), .B2(new_n472), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n735), .A2(new_n299), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(KEYINPUT33), .B(G317), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n741), .A2(new_n750), .A3(new_n756), .A4(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n273), .B1(new_n759), .B2(new_n351), .C1(new_n221), .C2(new_n752), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n761), .A2(new_n219), .B1(new_n757), .B2(new_n227), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n740), .C2(G50), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G58), .A2(new_n745), .B1(new_n755), .B2(G77), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT32), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n771), .B1(new_n748), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n749), .A2(KEYINPUT32), .A3(G159), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n770), .A2(KEYINPUT90), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n769), .B(new_n775), .C1(KEYINPUT90), .C2(new_n770), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n765), .A2(KEYINPUT92), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n766), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n734), .B1(new_n778), .B2(new_n723), .ZN(new_n779));
  INV_X1    g0579(.A(new_n722), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n643), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n719), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT93), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(G396));
  NAND2_X1  g0584(.A1(new_n361), .A2(new_n637), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n363), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n367), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n366), .A2(new_n648), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n699), .A2(new_n702), .A3(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n789), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n698), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(new_n695), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n717), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n790), .A2(new_n792), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n794), .A2(KEYINPUT97), .B1(new_n694), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(KEYINPUT97), .B2(new_n794), .ZN(new_n797));
  INV_X1    g0597(.A(new_n723), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G143), .A2(new_n745), .B1(new_n755), .B2(G159), .ZN(new_n799));
  INV_X1    g0599(.A(G150), .ZN(new_n800));
  INV_X1    g0600(.A(G137), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n799), .B1(new_n800), .B2(new_n761), .C1(new_n739), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT94), .B(KEYINPUT34), .Z(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n729), .B1(new_n806), .B2(new_n748), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT95), .Z(new_n808));
  INV_X1    g0608(.A(new_n759), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G68), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n202), .B2(new_n752), .C1(new_n225), .C2(new_n757), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n805), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n803), .B2(new_n804), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n740), .A2(G303), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n752), .A2(new_n351), .B1(new_n754), .B2(new_n506), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n744), .A2(new_n472), .B1(new_n748), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n762), .A2(G283), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n316), .B1(new_n759), .B2(new_n221), .ZN(new_n820));
  INV_X1    g0620(.A(new_n757), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(G97), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n814), .A2(new_n818), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n798), .B1(new_n813), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n723), .A2(new_n720), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n717), .B(new_n824), .C1(new_n272), .C2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT96), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n721), .B2(new_n791), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n797), .A2(new_n828), .ZN(G384));
  AOI211_X1 g0629(.A(new_n506), .B(new_n215), .C1(new_n564), .C2(KEYINPUT35), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(KEYINPUT35), .B2(new_n564), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT36), .Z(new_n832));
  OR3_X1    g0632(.A1(new_n217), .A2(new_n272), .A3(new_n385), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n202), .A2(G68), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n206), .B(G13), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT16), .B1(new_n426), .B2(new_n406), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n384), .B1(new_n837), .B2(new_n399), .ZN(new_n838));
  INV_X1    g0638(.A(new_n635), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n422), .A2(new_n430), .B1(new_n838), .B2(new_n588), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT98), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n380), .A2(new_n381), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n397), .A2(new_n219), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n389), .B1(new_n845), .B2(new_n388), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n427), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n844), .B1(new_n847), .B2(new_n384), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n434), .A2(new_n848), .A3(KEYINPUT98), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT37), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n434), .A2(KEYINPUT37), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT100), .B1(new_n430), .B2(new_n635), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT100), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n408), .A2(new_n853), .A3(new_n839), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n413), .A2(KEYINPUT99), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT99), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n382), .A2(new_n408), .A3(new_n412), .A4(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n851), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n850), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n840), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n436), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT101), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n408), .A2(new_n853), .A3(new_n839), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n853), .B1(new_n408), .B2(new_n839), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n431), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n856), .A2(new_n858), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n430), .A2(new_n844), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n434), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n865), .B1(new_n872), .B2(new_n855), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n864), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n866), .A2(new_n867), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n431), .A2(new_n589), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n859), .A3(KEYINPUT101), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n875), .B1(new_n594), .B2(new_n590), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n874), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n863), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n690), .A2(KEYINPUT30), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n886), .B(new_n682), .C1(new_n691), .C2(new_n677), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT31), .B(new_n637), .C1(new_n887), .C2(new_n680), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n686), .A2(new_n687), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n345), .A2(new_n343), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n344), .B1(new_n320), .B2(G169), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n347), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n347), .A2(new_n637), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n592), .A3(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n347), .B(new_n637), .C1(new_n346), .C2(new_n338), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n789), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT103), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT103), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n889), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n898), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n889), .A2(new_n896), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT98), .B1(new_n434), .B2(new_n848), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n838), .A2(new_n588), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n431), .A2(new_n842), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n906), .A3(new_n840), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n870), .B1(KEYINPUT37), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n433), .A2(new_n435), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n840), .B1(new_n909), .B2(new_n415), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n908), .A2(new_n882), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n860), .B2(new_n862), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n902), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n439), .A2(new_n889), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n645), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n792), .A2(new_n788), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n882), .B1(new_n908), .B2(new_n910), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n863), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n894), .A2(new_n895), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n590), .A2(new_n635), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n346), .A2(new_n347), .A3(new_n648), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n883), .B2(new_n884), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n922), .A2(KEYINPUT39), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n926), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n439), .A2(new_n703), .A3(new_n710), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n934), .A2(new_n597), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n919), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n206), .B2(new_n713), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n919), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n836), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT104), .ZN(G367));
  INV_X1    g0741(.A(new_n730), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n724), .B1(new_n210), .B2(new_n357), .C1(new_n942), .C2(new_n239), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n943), .A2(new_n716), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n612), .A2(new_n637), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n614), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n609), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n757), .A2(new_n219), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n273), .B1(new_n752), .B2(new_n225), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(G159), .C2(new_n762), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n744), .A2(new_n800), .B1(new_n759), .B2(new_n272), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n754), .A2(new_n202), .B1(new_n748), .B2(new_n801), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(G143), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n950), .B(new_n953), .C1(new_n954), .C2(new_n739), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n753), .A2(G116), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT46), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n956), .A2(new_n957), .B1(new_n761), .B2(new_n472), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n729), .B(new_n958), .C1(G107), .C2(new_n821), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n816), .B2(new_n739), .ZN(new_n960));
  INV_X1    g0760(.A(G317), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n754), .A2(new_n758), .B1(new_n748), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n809), .A2(G97), .ZN(new_n963));
  INV_X1    g0763(.A(G303), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n964), .B2(new_n744), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT109), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n956), .A2(new_n957), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n962), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n955), .B1(new_n960), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT47), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n944), .B1(new_n947), .B2(new_n780), .C1(new_n971), .C2(new_n798), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n581), .B(new_n584), .C1(new_n569), .C2(new_n658), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n617), .A2(new_n659), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n661), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT45), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n661), .A2(new_n975), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n653), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n651), .B1(new_n654), .B2(new_n637), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(KEYINPUT107), .A3(new_n656), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(KEYINPUT107), .B2(new_n982), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n647), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n711), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n711), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n664), .B(KEYINPUT41), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n715), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n657), .A2(new_n975), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(KEYINPUT42), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n584), .B1(new_n973), .B2(new_n482), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n994), .A2(KEYINPUT42), .B1(new_n658), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT105), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n998), .B2(new_n997), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT106), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1000), .B(new_n1002), .C1(KEYINPUT43), .C2(new_n947), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n652), .A2(new_n975), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1009), .B(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n972), .B1(new_n993), .B2(new_n1012), .ZN(G387));
  INV_X1    g0813(.A(new_n724), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n668), .A2(new_n725), .B1(G107), .B2(new_n210), .ZN(new_n1015));
  AOI211_X1 g0815(.A(G45), .B(new_n667), .C1(G68), .C2(G77), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n256), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n942), .B1(new_n236), .B2(G45), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G77), .A2(new_n753), .B1(new_n755), .B2(G68), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n258), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n202), .B2(new_n744), .C1(new_n1025), .C2(new_n761), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n739), .A2(new_n772), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n757), .A2(new_n357), .ZN(new_n1028));
  XOR2_X1   g0828(.A(KEYINPUT111), .B(G150), .Z(new_n1029));
  OAI211_X1 g0829(.A(new_n963), .B(new_n729), .C1(new_n748), .C2(new_n1029), .ZN(new_n1030));
  NOR4_X1   g0830(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n745), .B1(new_n755), .B2(G303), .ZN(new_n1032));
  INV_X1    g0832(.A(G322), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n816), .B2(new_n761), .C1(new_n739), .C2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n753), .A2(G294), .B1(new_n821), .B2(G283), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(G326), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n759), .A2(new_n506), .B1(new_n748), .B2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1041), .A2(new_n729), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1031), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n716), .B1(new_n1014), .B2(new_n1023), .C1(new_n1046), .C2(new_n798), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n651), .B2(new_n722), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n985), .B2(new_n715), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n986), .A2(new_n664), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n985), .A2(new_n711), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G393));
  OR2_X1    g0852(.A1(new_n988), .A2(new_n989), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n981), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n665), .B1(new_n1054), .B2(new_n986), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G68), .A2(new_n753), .B1(new_n809), .B2(G87), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n729), .C1(new_n954), .C2(new_n748), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT112), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n739), .A2(new_n800), .B1(new_n772), .B2(new_n744), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n757), .A2(new_n272), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n754), .A2(new_n256), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G50), .C2(new_n762), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1059), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n739), .A2(new_n961), .B1(new_n816), .B2(new_n744), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n316), .B1(new_n759), .B2(new_n351), .C1(new_n761), .C2(new_n964), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G283), .A2(new_n753), .B1(new_n755), .B2(G294), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1033), .B2(new_n748), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(G116), .C2(new_n821), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n798), .B1(new_n1065), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n942), .A2(new_n243), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1014), .B(new_n1074), .C1(G97), .C2(new_n663), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n717), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n975), .B2(new_n780), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1054), .B2(new_n714), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1056), .A2(new_n1078), .ZN(G390));
  OAI221_X1 g0879(.A(new_n810), .B1(new_n506), .B2(new_n744), .C1(new_n472), .C2(new_n748), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n316), .B1(new_n752), .B2(new_n221), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1080), .A2(new_n1062), .A3(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n762), .A2(G107), .B1(new_n755), .B2(G97), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n740), .A2(G283), .B1(KEYINPUT117), .B2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(KEYINPUT117), .C2(new_n1083), .ZN(new_n1085));
  INV_X1    g0885(.A(G128), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n739), .A2(new_n1086), .B1(new_n806), .B2(new_n744), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT116), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT54), .B(G143), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n761), .A2(new_n801), .B1(new_n754), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT115), .ZN(new_n1091));
  INV_X1    g0891(.A(G125), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n273), .B1(new_n748), .B2(new_n1092), .C1(new_n202), .C2(new_n759), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G159), .B2(new_n821), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1029), .A2(new_n752), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1085), .B1(new_n1088), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n798), .B1(new_n1098), .B2(KEYINPUT118), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(KEYINPUT118), .B2(new_n1098), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n717), .B1(new_n1025), .B2(new_n825), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n932), .C2(new_n721), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n788), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n698), .B2(new_n791), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n923), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n927), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n930), .A2(new_n931), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n709), .A2(new_n787), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n788), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n928), .B1(new_n1109), .B2(new_n923), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n885), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n693), .A2(G330), .A3(new_n791), .A4(new_n923), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1107), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n889), .A2(G330), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n896), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1102), .B1(new_n1118), .B2(new_n714), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT114), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n889), .A2(G330), .A3(new_n791), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1105), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1103), .B1(new_n709), .B2(new_n787), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1112), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n693), .A2(G330), .A3(new_n791), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1114), .A2(new_n896), .B1(new_n1126), .B2(new_n1105), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1127), .B2(new_n1104), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n439), .A2(new_n1114), .ZN(new_n1129));
  AND4_X1   g0929(.A1(new_n597), .A2(new_n1128), .A3(new_n934), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT113), .B1(new_n1117), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1115), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1107), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1134), .A2(new_n1130), .A3(KEYINPUT113), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1121), .B(new_n664), .C1(new_n1131), .C2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1117), .A2(new_n1130), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT113), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n665), .B1(new_n1144), .B2(new_n1136), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n1121), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1120), .B1(new_n1141), .B2(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(new_n825), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n716), .B1(G50), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n394), .A2(new_n395), .A3(new_n281), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n744), .A2(new_n351), .B1(new_n759), .B2(new_n225), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n547), .C2(new_n755), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n752), .A2(new_n272), .B1(new_n748), .B2(new_n758), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n948), .B(new_n1153), .C1(G97), .C2(new_n762), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n506), .C2(new_n739), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G50), .B1(new_n267), .B2(new_n281), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1155), .A2(new_n1156), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1086), .A2(new_n744), .B1(new_n752), .B2(new_n1089), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G137), .B2(new_n755), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n762), .A2(G132), .B1(new_n821), .B2(G150), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n1092), .C2(new_n739), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n267), .B(new_n281), .C1(new_n759), .C2(new_n772), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G124), .B2(new_n749), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1158), .B1(new_n1156), .B2(new_n1155), .C1(new_n1163), .C2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1149), .B1(new_n1168), .B2(new_n723), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n264), .A2(new_n635), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT55), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n306), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n306), .A2(new_n1172), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OR3_X1    g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1169), .B1(new_n1179), .B2(new_n721), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT120), .Z(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n645), .B1(new_n913), .B2(new_n914), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1179), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n880), .A2(new_n882), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT102), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n911), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n898), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1183), .B(new_n1184), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1184), .B1(new_n902), .B2(new_n1183), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n933), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n924), .A2(new_n925), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1195), .A2(new_n929), .B1(KEYINPUT39), .B2(new_n922), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1196), .B2(new_n927), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1189), .B1(new_n1195), .B2(new_n863), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n915), .A2(G330), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1179), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1197), .A2(new_n1200), .A3(new_n1190), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1193), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1197), .A2(new_n1200), .A3(KEYINPUT121), .A4(new_n1190), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1182), .B1(new_n1205), .B2(new_n714), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n935), .A2(new_n1129), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1208), .B1(new_n1144), .B2(new_n1136), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT122), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1193), .A2(new_n1201), .A3(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(KEYINPUT122), .B(new_n933), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n664), .B1(new_n1213), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1207), .B1(new_n1212), .B2(new_n1218), .ZN(G375));
  INV_X1    g1019(.A(new_n1128), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1208), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1130), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n992), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1105), .A2(new_n720), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n716), .B1(G68), .B2(new_n1148), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n273), .B(new_n1028), .C1(G77), .C2(new_n809), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n227), .A2(new_n752), .B1(new_n744), .B2(new_n758), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G303), .B2(new_n749), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n762), .A2(G116), .B1(new_n755), .B2(G107), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1226), .B(new_n1228), .C1(KEYINPUT123), .C2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT123), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n472), .B2(new_n739), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n739), .A2(new_n806), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n744), .A2(new_n801), .B1(new_n754), .B2(new_n800), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G159), .B2(new_n753), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G58), .A2(new_n809), .B1(new_n749), .B2(G128), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1089), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n762), .A2(new_n1237), .B1(new_n821), .B2(G50), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n729), .A3(new_n1236), .A4(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1230), .A2(new_n1232), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1225), .B1(new_n1240), .B2(new_n723), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1128), .A2(new_n715), .B1(new_n1224), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1223), .A2(new_n1242), .ZN(G381));
  OR2_X1    g1043(.A1(new_n993), .A2(new_n1012), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1056), .A2(new_n1078), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n972), .ZN(new_n1246));
  OR3_X1    g1046(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1246), .A2(G381), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1139), .B1(new_n1145), .B2(new_n1121), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n664), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT114), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1119), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1216), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n665), .B1(new_n1253), .B2(new_n1210), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT57), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1213), .B2(new_n1205), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1206), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1248), .A2(new_n1252), .A3(new_n1257), .ZN(G407));
  INV_X1    g1058(.A(G213), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(G343), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1252), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G407), .A2(G213), .A3(new_n1261), .ZN(G409));
  NAND2_X1  g1062(.A1(G390), .A2(G387), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(G393), .B(new_n783), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1246), .A3(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1263), .A2(new_n1246), .A3(new_n1270), .A4(new_n1266), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT125), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1221), .B1(new_n1276), .B2(new_n1130), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1208), .A2(KEYINPUT60), .A3(new_n1220), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n664), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1279), .A3(new_n1242), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G384), .A2(new_n1281), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1275), .A2(new_n1279), .A3(new_n1242), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1260), .A2(G2897), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1285), .B(new_n1286), .Z(new_n1287));
  NAND3_X1  g1087(.A1(new_n1215), .A2(new_n715), .A3(new_n1216), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1180), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1213), .A2(new_n1205), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(new_n992), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(G378), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT124), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(G375), .B2(new_n1252), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(G378), .A2(new_n1295), .A3(KEYINPUT124), .A4(new_n1207), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1292), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1287), .B1(new_n1297), .B2(new_n1260), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1285), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1297), .A2(new_n1260), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1273), .B(new_n1298), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1292), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1260), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n1285), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1272), .B1(new_n1302), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1272), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1300), .A2(KEYINPUT63), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1311), .A2(new_n1273), .A3(new_n1312), .A4(new_n1298), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(G405));
  AND3_X1   g1114(.A1(new_n1269), .A2(new_n1285), .A3(new_n1271), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1285), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G375), .A2(new_n1252), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1303), .A2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(KEYINPUT127), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1317), .B(new_n1320), .ZN(G402));
endmodule


