//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT83), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT3), .B1(new_n197), .B2(G107), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G104), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(G107), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n198), .A2(new_n201), .A3(new_n202), .A4(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n197), .A2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n200), .A2(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(G101), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT10), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(G128), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n216), .B2(new_n212), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n215), .B2(G143), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n211), .A2(KEYINPUT65), .A3(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(new_n211), .B2(G146), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n215), .A3(G143), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n221), .A2(new_n222), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n210), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT0), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(new_n225), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n221), .A2(new_n231), .A3(new_n222), .A4(new_n224), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n222), .A2(new_n224), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n235), .A2(KEYINPUT66), .A3(new_n231), .A4(new_n221), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n216), .A2(new_n212), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n198), .A2(new_n201), .A3(new_n203), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G101), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n246), .A3(G101), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n229), .B1(new_n242), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n211), .A2(KEYINPUT65), .A3(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT65), .B1(new_n211), .B2(G146), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n222), .B(new_n224), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n214), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(KEYINPUT84), .A3(new_n214), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n227), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n204), .A2(new_n207), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n251), .B(KEYINPUT10), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n215), .A2(G143), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n225), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n235), .B2(new_n221), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n227), .B1(new_n264), .B2(KEYINPUT84), .ZN(new_n265));
  INV_X1    g079(.A(new_n258), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT85), .B1(new_n267), .B2(new_n209), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n250), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT87), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G137), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT11), .A3(G134), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G137), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(G134), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT11), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g094(.A(KEYINPUT67), .B(KEYINPUT11), .C1(new_n272), .C2(G134), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G131), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n273), .A2(new_n275), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n279), .B1(new_n274), .B2(G137), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(new_n277), .A3(new_n279), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G131), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT87), .B(new_n250), .C1(new_n261), .C2(new_n268), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n271), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n291), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(new_n250), .C1(new_n261), .C2(new_n268), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n196), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n228), .A2(new_n260), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n267), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n291), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT12), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n297), .B1(new_n259), .B2(new_n260), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n294), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n294), .B1(new_n267), .B2(new_n298), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT86), .B1(new_n305), .B2(KEYINPUT12), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n295), .A2(new_n196), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n190), .B(new_n191), .C1(new_n296), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n308), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n295), .B1(new_n304), .B2(new_n306), .ZN(new_n312));
  INV_X1    g126(.A(new_n196), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n293), .A2(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G469), .B1(new_n314), .B2(G902), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n189), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G125), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n329), .B2(new_n318), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n322), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n215), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n322), .A2(G146), .A3(new_n324), .A4(new_n330), .ZN(new_n333));
  NOR2_X1   g147(.A1(G237), .A2(G953), .ZN(new_n334));
  AOI21_X1  g148(.A(G143), .B1(new_n334), .B2(G214), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(G143), .A3(G214), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT17), .A3(G131), .ZN(new_n339));
  INV_X1    g153(.A(new_n337), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n340), .B2(new_n335), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n289), .A3(new_n337), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT17), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n332), .A2(new_n333), .A3(new_n339), .A4(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G113), .B(G122), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n197), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n338), .A2(KEYINPUT18), .A3(G131), .ZN(new_n348));
  NAND2_X1  g162(.A1(KEYINPUT18), .A2(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n336), .A2(new_n337), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n329), .A2(G146), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n323), .A2(new_n215), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n345), .A2(new_n347), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n341), .A2(new_n342), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n215), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n333), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n354), .ZN(new_n361));
  INV_X1    g175(.A(new_n347), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(G475), .A2(G902), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n317), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  AOI211_X1 g181(.A(KEYINPUT20), .B(new_n367), .C1(new_n355), .C2(new_n363), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G475), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n345), .A2(new_n354), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n362), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT92), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n355), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n347), .B1(new_n345), .B2(new_n354), .ZN(new_n375));
  AOI21_X1  g189(.A(G902), .B1(new_n375), .B2(KEYINPUT92), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n370), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT69), .B(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G122), .ZN(new_n381));
  INV_X1    g195(.A(G116), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n382), .A2(G122), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n200), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G128), .B(G143), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n274), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n381), .A2(new_n387), .A3(new_n383), .ZN(new_n388));
  OAI21_X1  g202(.A(G107), .B1(new_n381), .B2(new_n387), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n384), .B(new_n386), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n225), .A2(G143), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n274), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n385), .ZN(new_n394));
  INV_X1    g208(.A(new_n384), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n200), .B1(new_n381), .B2(new_n383), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G217), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n187), .A2(new_n398), .A3(G953), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n390), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n390), .B2(new_n397), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n191), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n379), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n194), .A2(G952), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(G234), .B2(G237), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n191), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT21), .B(G898), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G214), .B1(G237), .B2(G902), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G122), .ZN(new_n415));
  INV_X1    g229(.A(G119), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G116), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n418), .B1(new_n380), .B2(G119), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT2), .B(G113), .Z(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n382), .A2(KEYINPUT69), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(G116), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n424), .A3(G119), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n417), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT2), .B(G113), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n247), .A3(new_n245), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(KEYINPUT5), .A3(new_n417), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n417), .A2(KEYINPUT5), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(G113), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n421), .A3(new_n260), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n415), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT6), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n426), .A2(new_n427), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n420), .B1(new_n417), .B2(new_n425), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n434), .B(new_n415), .C1(new_n248), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT88), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n430), .A2(new_n443), .A3(new_n434), .A4(new_n415), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n437), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n436), .B1(new_n445), .B2(new_n435), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n242), .A2(new_n447), .A3(G125), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n240), .B1(new_n234), .B2(new_n236), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT89), .B1(new_n449), .B2(new_n327), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n217), .A2(new_n227), .A3(new_n327), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT90), .B(G224), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n194), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n194), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n448), .A2(new_n450), .A3(new_n455), .A4(new_n451), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n442), .A2(new_n444), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT7), .B1(new_n455), .B2(KEYINPUT91), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(KEYINPUT91), .B2(new_n455), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n448), .A2(new_n450), .A3(new_n451), .A4(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n451), .B1(new_n449), .B2(new_n327), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n464));
  OAI21_X1  g278(.A(G113), .B1(new_n417), .B2(KEYINPUT5), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n419), .B2(KEYINPUT5), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n208), .B1(new_n466), .B2(new_n438), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n434), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n415), .B(KEYINPUT8), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n463), .A2(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n459), .A2(new_n462), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n471), .A2(new_n191), .ZN(new_n472));
  OAI21_X1  g286(.A(G210), .B1(G237), .B2(G902), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n458), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n458), .B2(new_n472), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n414), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n316), .A2(new_n413), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n334), .A2(G210), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT27), .Z(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G101), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n481), .B(new_n482), .Z(new_n483));
  AOI21_X1  g297(.A(new_n289), .B1(new_n278), .B2(new_n275), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n288), .B2(new_n289), .ZN(new_n485));
  AOI221_X4 g299(.A(new_n429), .B1(new_n485), .B2(new_n228), .C1(new_n449), .C2(new_n291), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT68), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(KEYINPUT68), .A2(KEYINPUT30), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n291), .A2(new_n237), .A3(new_n241), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n485), .A2(new_n228), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  AND4_X1   g307(.A1(new_n487), .A2(new_n491), .A3(new_n488), .A4(new_n492), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n429), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n486), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n491), .A2(new_n492), .ZN(new_n498));
  INV_X1    g312(.A(new_n489), .ZN(new_n499));
  INV_X1    g313(.A(new_n490), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n491), .A2(new_n487), .A3(new_n488), .A4(new_n492), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT70), .A3(new_n429), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n483), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n440), .B1(new_n491), .B2(new_n492), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT28), .B1(new_n486), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(KEYINPUT28), .C1(new_n486), .C2(new_n506), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n486), .A2(KEYINPUT28), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n508), .A2(new_n483), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n479), .B1(new_n505), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n483), .ZN(new_n516));
  INV_X1    g330(.A(new_n486), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n440), .B1(new_n501), .B2(new_n502), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(KEYINPUT70), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n496), .B(new_n440), .C1(new_n501), .C2(new_n502), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n521), .A2(KEYINPUT72), .A3(new_n513), .A4(new_n512), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n511), .A2(new_n507), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n516), .A2(new_n513), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n515), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G472), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n495), .A2(new_n496), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n528), .A2(new_n483), .A3(new_n517), .A4(new_n504), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT31), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n516), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n497), .A2(new_n533), .A3(new_n483), .A4(new_n504), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT32), .ZN(new_n536));
  NOR2_X1   g350(.A1(G472), .A2(G902), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n527), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT82), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT81), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT22), .B(G137), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n225), .A2(G119), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n416), .A2(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT78), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT74), .ZN(new_n558));
  NAND2_X1  g372(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n225), .B2(G119), .ZN(new_n560));
  NOR2_X1   g374(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n416), .A2(G128), .B1(KEYINPUT73), .B2(KEYINPUT23), .ZN(new_n563));
  INV_X1    g377(.A(new_n561), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT74), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n557), .B1(new_n566), .B2(new_n548), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT77), .B(G110), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n556), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n333), .A2(new_n352), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n547), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n560), .A2(new_n558), .A3(new_n561), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT74), .B1(new_n563), .B2(new_n564), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n548), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n557), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n568), .ZN(new_n576));
  INV_X1    g390(.A(new_n556), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n333), .A2(new_n352), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n550), .A2(new_n551), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n332), .B2(new_n333), .ZN(new_n583));
  INV_X1    g397(.A(G110), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n567), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n546), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n569), .A2(new_n547), .A3(new_n570), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT79), .B1(new_n578), .B2(new_n579), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT80), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n581), .A2(new_n591), .A3(new_n585), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n586), .B1(new_n593), .B2(new_n546), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n542), .B1(new_n594), .B2(G902), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n581), .A2(new_n591), .A3(new_n585), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n591), .B1(new_n581), .B2(new_n585), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n546), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n586), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(KEYINPUT25), .A3(new_n191), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n398), .B1(G234), .B2(new_n191), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n602), .A2(new_n603), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n540), .A2(new_n541), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n541), .B1(new_n540), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n478), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NAND2_X1  g423(.A1(new_n535), .A2(new_n191), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n535), .A2(new_n537), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n605), .A3(new_n316), .A4(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n476), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(KEYINPUT93), .B(new_n414), .C1(new_n474), .C2(new_n475), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n412), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n404), .A2(G902), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT33), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n390), .A2(new_n397), .ZN(new_n624));
  INV_X1    g438(.A(new_n399), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n623), .B1(new_n626), .B2(new_n400), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n621), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT94), .B1(new_n403), .B2(new_n404), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT33), .B1(new_n401), .B2(new_n402), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n623), .A3(new_n400), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT94), .A3(new_n621), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n630), .B(new_n634), .C1(new_n369), .C2(new_n377), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n620), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n614), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  NOR2_X1   g453(.A1(new_n378), .A2(new_n406), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n620), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n614), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT96), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NAND3_X1  g461(.A1(new_n611), .A2(new_n612), .A3(new_n316), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT25), .B1(new_n600), .B2(new_n191), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n542), .B(G902), .C1(new_n598), .C2(new_n599), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n603), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n546), .A2(KEYINPUT36), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n593), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n593), .A2(new_n653), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n604), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n413), .A3(new_n477), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT37), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n310), .A2(new_n315), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n188), .ZN(new_n664));
  INV_X1    g478(.A(new_n603), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n595), .B2(new_n601), .ZN(new_n666));
  INV_X1    g480(.A(new_n657), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n410), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n409), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n640), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n616), .B2(new_n617), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n669), .A2(new_n540), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n225), .ZN(G30));
  OR2_X1    g491(.A1(new_n379), .A2(new_n406), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n668), .A2(new_n414), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT97), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n673), .B(KEYINPUT39), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n316), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT40), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n519), .A2(new_n520), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n516), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n486), .A2(new_n506), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n191), .B1(new_n689), .B2(new_n483), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n538), .B2(new_n539), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n458), .A2(new_n472), .ZN(new_n695));
  INV_X1    g509(.A(new_n473), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n458), .A2(new_n472), .A3(new_n473), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT38), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n684), .A2(new_n685), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n682), .A2(new_n694), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  INV_X1    g517(.A(new_n673), .ZN(new_n704));
  AOI211_X1 g518(.A(new_n635), .B(new_n704), .C1(new_n616), .C2(new_n617), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n669), .A2(new_n705), .A3(new_n540), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  INV_X1    g521(.A(new_n605), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n612), .A2(KEYINPUT32), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n708), .B1(new_n711), .B2(new_n527), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT84), .B1(new_n254), .B2(new_n214), .ZN(new_n713));
  INV_X1    g527(.A(new_n227), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n208), .B1(new_n715), .B2(new_n258), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n251), .B1(new_n716), .B2(KEYINPUT10), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n267), .A2(KEYINPUT85), .A3(new_n209), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n249), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n291), .B1(new_n719), .B2(KEYINPUT87), .ZN(new_n720));
  INV_X1    g534(.A(new_n292), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n295), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n309), .B1(new_n722), .B2(new_n313), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n723), .B2(G902), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n188), .A3(new_n310), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT98), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT98), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n724), .A2(new_n727), .A3(new_n188), .A4(new_n310), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n712), .A2(new_n729), .A3(new_n636), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND3_X1  g546(.A1(new_n712), .A2(new_n729), .A3(new_n642), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  INV_X1    g548(.A(KEYINPUT99), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT93), .B1(new_n699), .B2(new_n414), .ZN(new_n736));
  INV_X1    g550(.A(new_n617), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n735), .B1(new_n738), .B2(new_n725), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n724), .A2(new_n188), .A3(new_n310), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(KEYINPUT99), .A3(new_n618), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n709), .A2(new_n710), .B1(G472), .B2(new_n526), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n658), .A2(new_n413), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  AOI21_X1  g561(.A(new_n412), .B1(new_n616), .B2(new_n617), .ZN(new_n748));
  AND4_X1   g562(.A1(new_n748), .A2(new_n726), .A3(new_n679), .A4(new_n728), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n530), .B(new_n534), .C1(new_n483), .C2(new_n523), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n537), .B(KEYINPUT100), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n610), .A2(G472), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(new_n605), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  INV_X1    g569(.A(KEYINPUT102), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n635), .B2(new_n704), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT94), .ZN(new_n758));
  INV_X1    g572(.A(new_n621), .ZN(new_n759));
  AOI211_X1 g573(.A(new_n758), .B(new_n759), .C1(new_n631), .C2(new_n632), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n628), .B2(new_n629), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n378), .A2(new_n761), .A3(KEYINPUT102), .A4(new_n673), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n739), .B2(new_n741), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n750), .A2(new_n751), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n611), .A2(new_n658), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT101), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n752), .A2(KEYINPUT101), .A3(new_n658), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  NAND2_X1  g587(.A1(new_n540), .A2(new_n605), .ZN(new_n774));
  INV_X1    g588(.A(new_n414), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n699), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n316), .A2(new_n763), .A3(KEYINPUT42), .A4(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT103), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n777), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT103), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n780), .A3(new_n540), .A4(new_n605), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  INV_X1    g596(.A(new_n776), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n664), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n540), .A3(new_n605), .A4(new_n763), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n778), .A2(new_n781), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(KEYINPUT104), .B(G131), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G33));
  INV_X1    g602(.A(new_n674), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n784), .A2(new_n540), .A3(new_n605), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  NAND2_X1  g605(.A1(new_n611), .A2(new_n612), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n630), .A2(new_n634), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n378), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT43), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(KEYINPUT44), .A3(new_n658), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n776), .ZN(new_n797));
  INV_X1    g611(.A(new_n310), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n314), .A2(KEYINPUT45), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n314), .A2(KEYINPUT45), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(G469), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(G469), .A2(G902), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n798), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n801), .A2(KEYINPUT46), .A3(new_n802), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n189), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n792), .A2(new_n658), .A3(new_n795), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n797), .A2(new_n683), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT105), .B(G137), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G39));
  NOR2_X1   g627(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g629(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n816));
  AOI211_X1 g630(.A(new_n189), .B(new_n816), .C1(new_n805), .C2(new_n806), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n783), .A2(new_n635), .A3(new_n704), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n743), .A2(new_n708), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(new_n319), .ZN(G42));
  NOR2_X1   g635(.A1(G952), .A2(G953), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT115), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT110), .B1(new_n740), .B2(new_n776), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n672), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n740), .A2(KEYINPUT110), .A3(new_n776), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n605), .A2(new_n826), .A3(new_n693), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n379), .A3(new_n793), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n795), .A2(new_n409), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n753), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT109), .ZN(new_n834));
  OR3_X1    g648(.A1(new_n700), .A2(new_n725), .A3(new_n414), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n832), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n833), .A2(KEYINPUT109), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n834), .B(new_n837), .C1(new_n832), .C2(new_n835), .ZN(new_n838));
  INV_X1    g652(.A(new_n771), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n826), .A2(new_n795), .A3(new_n827), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n836), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n824), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n836), .A2(new_n838), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n840), .A2(new_n839), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(KEYINPUT111), .A3(new_n829), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n832), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n815), .A2(new_n817), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n724), .A2(new_n310), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n188), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n776), .B(new_n846), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n842), .A2(KEYINPUT51), .A3(new_n845), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  INV_X1    g666(.A(new_n850), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n843), .A2(new_n829), .A3(new_n844), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n846), .A2(new_n742), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT113), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n408), .B(KEYINPUT112), .Z(new_n858));
  INV_X1    g672(.A(new_n635), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n858), .B1(new_n828), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n840), .A2(new_n774), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT48), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n851), .A2(new_n855), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT114), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n851), .A2(new_n867), .A3(new_n855), .A4(new_n864), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n678), .B1(new_n616), .B2(new_n617), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n666), .A2(new_n667), .A3(new_n704), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n692), .A2(new_n316), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n706), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n676), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n772), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n676), .B1(new_n765), .B2(new_n771), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n706), .A2(new_n872), .A3(KEYINPUT52), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT108), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT108), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n785), .A2(new_n782), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n780), .B1(new_n712), .B2(new_n779), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n743), .A2(new_n777), .A3(KEYINPUT103), .A4(new_n708), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n784), .A2(new_n763), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n769), .B2(new_n770), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n783), .A2(new_n407), .A3(new_n704), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n669), .A2(new_n889), .A3(new_n540), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n790), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n641), .A2(new_n635), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n619), .A3(new_n477), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n613), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n749), .B2(new_n753), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n660), .B1(new_n742), .B2(new_n745), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n712), .B(new_n729), .C1(new_n642), .C2(new_n636), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n608), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n893), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n882), .A2(new_n902), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n608), .A2(new_n897), .A3(new_n898), .A4(new_n899), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n764), .A2(new_n664), .A3(new_n783), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n752), .A2(KEYINPUT101), .A3(new_n658), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT101), .B1(new_n752), .B2(new_n658), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n790), .A3(new_n890), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n786), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n875), .A2(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n903), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n911), .A2(new_n912), .A3(new_n901), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(KEYINPUT107), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n893), .A2(new_n900), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT107), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n920), .A3(new_n882), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n921), .B2(new_n901), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n915), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n823), .B1(new_n869), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n794), .A2(new_n188), .A3(new_n414), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n925), .B(new_n700), .C1(KEYINPUT49), .C2(new_n848), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n848), .A2(KEYINPUT49), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n926), .A2(new_n605), .A3(new_n693), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n924), .A2(new_n928), .ZN(G75));
  NOR2_X1   g743(.A1(new_n194), .A2(G952), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n903), .A2(new_n913), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G902), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT56), .B1(new_n934), .B2(G210), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n446), .B(new_n457), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n931), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  AOI211_X1 g753(.A(KEYINPUT56), .B(new_n937), .C1(new_n934), .C2(G210), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(new_n802), .B(KEYINPUT116), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT57), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n903), .A2(new_n913), .A3(new_n914), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n914), .B1(new_n903), .B2(new_n913), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT117), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT117), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n723), .B(KEYINPUT118), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n933), .A2(new_n801), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n930), .B1(new_n951), .B2(new_n952), .ZN(G54));
  NAND2_X1  g767(.A1(KEYINPUT58), .A2(G475), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT119), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n355), .B(new_n363), .C1(new_n933), .C2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n932), .A2(G902), .A3(new_n364), .A4(new_n955), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n931), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n957), .A2(KEYINPUT120), .A3(new_n931), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n633), .B1(new_n923), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n633), .A2(new_n965), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT52), .B1(new_n878), .B2(new_n873), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n878), .A2(new_n879), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT108), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT108), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n904), .A2(new_n910), .A3(KEYINPUT53), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n877), .A2(new_n969), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT53), .B1(new_n976), .B2(new_n918), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT54), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n967), .B1(new_n978), .B2(new_n915), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT121), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n930), .ZN(new_n981));
  INV_X1    g795(.A(new_n967), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n944), .B2(new_n945), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT121), .B1(new_n983), .B2(new_n931), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n966), .A2(new_n981), .A3(new_n984), .ZN(G63));
  NOR2_X1   g799(.A1(new_n975), .A2(new_n977), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n655), .A2(new_n656), .ZN(new_n987));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  OR3_X1    g803(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n594), .B1(new_n986), .B2(new_n989), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n931), .A3(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n990), .A2(KEYINPUT61), .A3(new_n931), .A4(new_n991), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(G66));
  INV_X1    g810(.A(new_n411), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n194), .B1(new_n997), .B2(new_n453), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT122), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n904), .B2(G953), .ZN(new_n1000));
  INV_X1    g814(.A(new_n446), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(G898), .B2(new_n194), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1000), .B(new_n1002), .ZN(G69));
  NAND2_X1  g817(.A1(G900), .A2(G953), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n807), .A2(new_n712), .A3(new_n683), .A4(new_n870), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n811), .A2(new_n790), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(new_n820), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1007), .A2(new_n706), .A3(new_n886), .A4(new_n878), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1004), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n503), .B(KEYINPUT123), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n357), .A2(new_n358), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1010), .B(new_n1011), .Z(new_n1012));
  INV_X1    g826(.A(KEYINPUT62), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n702), .A2(new_n1013), .A3(new_n706), .A4(new_n878), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1014), .A2(KEYINPUT124), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n894), .A2(new_n776), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n684), .B(new_n1016), .C1(new_n606), .C2(new_n607), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n811), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT125), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT125), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n811), .A2(new_n1020), .A3(new_n1017), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n702), .A2(new_n706), .A3(new_n878), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n820), .B1(new_n1023), .B2(KEYINPUT62), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1014), .A2(KEYINPUT124), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1015), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1012), .A2(G953), .ZN(new_n1027));
  AOI22_X1  g841(.A1(new_n1009), .A2(new_n1012), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1028), .B(new_n1029), .ZN(G72));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  OAI21_X1  g846(.A(new_n1032), .B1(new_n1008), .B2(new_n900), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n687), .A2(new_n516), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n930), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n688), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1036), .B1(new_n922), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1032), .B1(new_n1026), .B2(new_n900), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n688), .B1(new_n1040), .B2(KEYINPUT126), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT126), .ZN(new_n1042));
  AND2_X1   g856(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n1043), .A2(new_n904), .A3(new_n1025), .A4(new_n1015), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1042), .B1(new_n1044), .B2(new_n1032), .ZN(new_n1045));
  OAI21_X1  g859(.A(KEYINPUT127), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1044), .A2(new_n1042), .A3(new_n1032), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1040), .A2(KEYINPUT126), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT127), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n688), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n1039), .B1(new_n1046), .B2(new_n1050), .ZN(G57));
endmodule


