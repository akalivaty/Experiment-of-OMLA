

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XOR2_X1 U324 ( .A(n453), .B(n452), .Z(n292) );
  XOR2_X1 U325 ( .A(G176GAT), .B(G120GAT), .Z(n293) );
  INV_X1 U326 ( .A(n554), .ZN(n395) );
  OR2_X1 U327 ( .A1(n563), .A2(n395), .ZN(n396) );
  XNOR2_X1 U328 ( .A(n372), .B(n293), .ZN(n373) );
  NOR2_X1 U329 ( .A1(n462), .A2(n568), .ZN(n449) );
  XNOR2_X1 U330 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U331 ( .A(n462), .B(KEYINPUT28), .Z(n528) );
  XOR2_X1 U332 ( .A(G99GAT), .B(G85GAT), .Z(n372) );
  XOR2_X1 U333 ( .A(G36GAT), .B(G218GAT), .Z(n410) );
  XOR2_X1 U334 ( .A(n372), .B(n410), .Z(n295) );
  XOR2_X1 U335 ( .A(G43GAT), .B(G134GAT), .Z(n311) );
  XOR2_X1 U336 ( .A(G50GAT), .B(G162GAT), .Z(n328) );
  XNOR2_X1 U337 ( .A(n311), .B(n328), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n300) );
  XNOR2_X1 U339 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n296), .B(KEYINPUT7), .ZN(n354) );
  XOR2_X1 U341 ( .A(n354), .B(KEYINPUT9), .Z(n298) );
  NAND2_X1 U342 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U344 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n302) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U348 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n304) );
  XNOR2_X1 U349 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n554) );
  XOR2_X1 U353 ( .A(KEYINPUT20), .B(KEYINPUT66), .Z(n310) );
  XNOR2_X1 U354 ( .A(G183GAT), .B(G71GAT), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n315) );
  XOR2_X1 U356 ( .A(KEYINPUT81), .B(G99GAT), .Z(n313) );
  XOR2_X1 U357 ( .A(G15GAT), .B(G127GAT), .Z(n392) );
  XNOR2_X1 U358 ( .A(n311), .B(n392), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U360 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U361 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U363 ( .A(n318), .B(KEYINPUT80), .Z(n321) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n319) );
  XNOR2_X1 U365 ( .A(n319), .B(G120GAT), .ZN(n441) );
  XNOR2_X1 U366 ( .A(n441), .B(KEYINPUT82), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U368 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n323) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(G176GAT), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n325) );
  XOR2_X1 U371 ( .A(G190GAT), .B(KEYINPUT19), .Z(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n415) );
  XOR2_X2 U373 ( .A(n326), .B(n415), .Z(n526) );
  INV_X1 U374 ( .A(n526), .ZN(n451) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(G78GAT), .ZN(n327) );
  XNOR2_X1 U376 ( .A(n327), .B(G148GAT), .ZN(n369) );
  XOR2_X1 U377 ( .A(n369), .B(n328), .Z(n330) );
  NAND2_X1 U378 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U380 ( .A(n331), .B(G204GAT), .Z(n333) );
  XOR2_X1 U381 ( .A(G22GAT), .B(G155GAT), .Z(n384) );
  XNOR2_X1 U382 ( .A(G218GAT), .B(n384), .ZN(n332) );
  XNOR2_X1 U383 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U384 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n335) );
  XNOR2_X1 U385 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U387 ( .A(n337), .B(n336), .Z(n342) );
  XOR2_X1 U388 ( .A(G211GAT), .B(KEYINPUT21), .Z(n339) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n338) );
  XNOR2_X1 U390 ( .A(n339), .B(n338), .ZN(n416) );
  XNOR2_X1 U391 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n340), .B(KEYINPUT2), .ZN(n434) );
  XNOR2_X1 U393 ( .A(n416), .B(n434), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n462) );
  XOR2_X1 U395 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n421) );
  XNOR2_X1 U396 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n399) );
  XOR2_X1 U397 ( .A(G141GAT), .B(G197GAT), .Z(n344) );
  XNOR2_X1 U398 ( .A(G15GAT), .B(G113GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n348) );
  XOR2_X1 U400 ( .A(KEYINPUT69), .B(G8GAT), .Z(n346) );
  XNOR2_X1 U401 ( .A(G22GAT), .B(G1GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U403 ( .A(n348), .B(n347), .Z(n353) );
  XOR2_X1 U404 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n350) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U407 ( .A(KEYINPUT68), .B(n351), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U409 ( .A(G50GAT), .B(G43GAT), .Z(n356) );
  XNOR2_X1 U410 ( .A(n354), .B(G36GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U413 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n360) );
  XNOR2_X1 U414 ( .A(KEYINPUT70), .B(KEYINPUT67), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U416 ( .A(G169GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n569) );
  XNOR2_X1 U418 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n376) );
  XNOR2_X1 U419 ( .A(G71GAT), .B(G57GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n364), .B(KEYINPUT13), .ZN(n380) );
  XOR2_X1 U421 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n366) );
  NAND2_X1 U422 ( .A1(G230GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U424 ( .A(n367), .B(KEYINPUT31), .Z(n371) );
  XNOR2_X1 U425 ( .A(G204GAT), .B(G92GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n368), .B(G64GAT), .ZN(n413) );
  XNOR2_X1 U427 ( .A(n369), .B(n413), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n374) );
  XOR2_X1 U429 ( .A(n380), .B(n375), .Z(n575) );
  XOR2_X1 U430 ( .A(n376), .B(n575), .Z(n559) );
  NOR2_X1 U431 ( .A1(n569), .A2(n559), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n377), .B(KEYINPUT46), .ZN(n397) );
  XOR2_X1 U433 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n383) );
  XOR2_X1 U434 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n379) );
  XNOR2_X1 U435 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U439 ( .A(G8GAT), .B(G183GAT), .Z(n407) );
  XOR2_X1 U440 ( .A(n407), .B(n384), .Z(n386) );
  NAND2_X1 U441 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U443 ( .A(n388), .B(n387), .Z(n394) );
  XOR2_X1 U444 ( .A(G64GAT), .B(G78GAT), .Z(n390) );
  XNOR2_X1 U445 ( .A(G1GAT), .B(G211GAT), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n551) );
  XNOR2_X1 U449 ( .A(KEYINPUT108), .B(n551), .ZN(n563) );
  NOR2_X1 U450 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n404) );
  XOR2_X1 U452 ( .A(n554), .B(KEYINPUT36), .Z(n583) );
  NAND2_X1 U453 ( .A1(n551), .A2(n583), .ZN(n400) );
  XNOR2_X1 U454 ( .A(KEYINPUT45), .B(n400), .ZN(n402) );
  NAND2_X1 U455 ( .A1(n575), .A2(n569), .ZN(n401) );
  NOR2_X1 U456 ( .A1(n402), .A2(n401), .ZN(n403) );
  NOR2_X1 U457 ( .A1(n404), .A2(n403), .ZN(n406) );
  INV_X1 U458 ( .A(KEYINPUT48), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n525) );
  XNOR2_X1 U460 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U462 ( .A(n410), .B(n409), .Z(n412) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U465 ( .A(n414), .B(n413), .Z(n419) );
  INV_X1 U466 ( .A(n415), .ZN(n417) );
  XNOR2_X1 U467 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U468 ( .A(n419), .B(n418), .ZN(n458) );
  NAND2_X1 U469 ( .A1(n525), .A2(n458), .ZN(n420) );
  XNOR2_X1 U470 ( .A(n421), .B(n420), .ZN(n446) );
  XOR2_X1 U471 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n423) );
  XNOR2_X1 U472 ( .A(G155GAT), .B(G148GAT), .ZN(n422) );
  XNOR2_X1 U473 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U474 ( .A(KEYINPUT75), .B(G85GAT), .Z(n425) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(G127GAT), .ZN(n424) );
  XNOR2_X1 U476 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U477 ( .A(n427), .B(n426), .ZN(n445) );
  XOR2_X1 U478 ( .A(KEYINPUT89), .B(G57GAT), .Z(n429) );
  XNOR2_X1 U479 ( .A(KEYINPUT4), .B(KEYINPUT88), .ZN(n428) );
  XNOR2_X1 U480 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U481 ( .A(KEYINPUT87), .B(KEYINPUT5), .Z(n431) );
  XNOR2_X1 U482 ( .A(KEYINPUT6), .B(KEYINPUT86), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U484 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U485 ( .A(G162GAT), .B(n434), .Z(n436) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U488 ( .A(G134GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U489 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U490 ( .A(n440), .B(KEYINPUT1), .Z(n443) );
  XNOR2_X1 U491 ( .A(G1GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U492 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n445), .B(n444), .ZN(n512) );
  NAND2_X1 U494 ( .A1(n446), .A2(n512), .ZN(n447) );
  XOR2_X1 U495 ( .A(n447), .B(KEYINPUT65), .Z(n568) );
  XNOR2_X1 U496 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n448) );
  XNOR2_X1 U497 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U498 ( .A1(n451), .A2(n450), .ZN(n562) );
  NOR2_X1 U499 ( .A1(n554), .A2(n562), .ZN(n454) );
  XOR2_X1 U500 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n453) );
  XNOR2_X1 U501 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n454), .B(n292), .ZN(G1351GAT) );
  INV_X1 U503 ( .A(n569), .ZN(n499) );
  AND2_X1 U504 ( .A1(n499), .A2(n575), .ZN(n486) );
  XOR2_X1 U505 ( .A(n458), .B(KEYINPUT27), .Z(n465) );
  NOR2_X1 U506 ( .A1(n512), .A2(n465), .ZN(n524) );
  NAND2_X1 U507 ( .A1(n528), .A2(n524), .ZN(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT83), .B(n526), .ZN(n455) );
  NOR2_X1 U509 ( .A1(n456), .A2(n455), .ZN(n471) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(KEYINPUT96), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT95), .ZN(n461) );
  INV_X1 U512 ( .A(n458), .ZN(n514) );
  NOR2_X1 U513 ( .A1(n526), .A2(n514), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n462), .A2(n459), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n461), .B(n460), .ZN(n467) );
  XOR2_X1 U516 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n464) );
  NAND2_X1 U517 ( .A1(n462), .A2(n526), .ZN(n463) );
  XOR2_X1 U518 ( .A(n464), .B(n463), .Z(n567) );
  NOR2_X1 U519 ( .A1(n567), .A2(n465), .ZN(n466) );
  NOR2_X1 U520 ( .A1(n467), .A2(n466), .ZN(n469) );
  INV_X1 U521 ( .A(n512), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U523 ( .A1(n471), .A2(n470), .ZN(n483) );
  XOR2_X1 U524 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n473) );
  NAND2_X1 U525 ( .A1(n551), .A2(n554), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n473), .B(n472), .ZN(n474) );
  NOR2_X1 U527 ( .A1(n483), .A2(n474), .ZN(n501) );
  NAND2_X1 U528 ( .A1(n486), .A2(n501), .ZN(n481) );
  NOR2_X1 U529 ( .A1(n512), .A2(n481), .ZN(n476) );
  XNOR2_X1 U530 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U531 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U533 ( .A1(n514), .A2(n481), .ZN(n478) );
  XOR2_X1 U534 ( .A(G8GAT), .B(n478), .Z(G1325GAT) );
  NOR2_X1 U535 ( .A1(n526), .A2(n481), .ZN(n480) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NOR2_X1 U538 ( .A1(n528), .A2(n481), .ZN(n482) );
  XOR2_X1 U539 ( .A(G22GAT), .B(n482), .Z(G1327GAT) );
  XNOR2_X1 U540 ( .A(KEYINPUT39), .B(KEYINPUT98), .ZN(n489) );
  NOR2_X1 U541 ( .A1(n551), .A2(n483), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n583), .A2(n484), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n485), .ZN(n511) );
  NAND2_X1 U544 ( .A1(n511), .A2(n486), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT38), .B(n487), .ZN(n494) );
  NOR2_X1 U546 ( .A1(n512), .A2(n494), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(G29GAT), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n494), .A2(n514), .ZN(n491) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n491), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n494), .A2(n526), .ZN(n492) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(n492), .Z(n493) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  XNOR2_X1 U554 ( .A(G50GAT), .B(KEYINPUT99), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n528), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n498) );
  XNOR2_X1 U558 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n503) );
  NOR2_X1 U560 ( .A1(n499), .A2(n559), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT101), .B(n500), .Z(n510) );
  NAND2_X1 U562 ( .A1(n510), .A2(n501), .ZN(n507) );
  NOR2_X1 U563 ( .A1(n512), .A2(n507), .ZN(n502) );
  XOR2_X1 U564 ( .A(n503), .B(n502), .Z(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT100), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n507), .ZN(n505) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n526), .A2(n507), .ZN(n506) );
  XOR2_X1 U569 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U570 ( .A1(n528), .A2(n507), .ZN(n509) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n510), .ZN(n520) );
  NOR2_X1 U574 ( .A1(n512), .A2(n520), .ZN(n513) );
  XOR2_X1 U575 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U576 ( .A1(n514), .A2(n520), .ZN(n515) );
  XOR2_X1 U577 ( .A(KEYINPUT104), .B(n515), .Z(n516) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U579 ( .A1(n526), .A2(n520), .ZN(n518) );
  XNOR2_X1 U580 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n528), .A2(n520), .ZN(n522) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n543) );
  NOR2_X1 U588 ( .A1(n526), .A2(n543), .ZN(n527) );
  XNOR2_X1 U589 ( .A(KEYINPUT110), .B(n527), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n539) );
  NOR2_X1 U591 ( .A1(n569), .A2(n539), .ZN(n530) );
  XOR2_X1 U592 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  NOR2_X1 U593 ( .A1(n539), .A2(n559), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n532) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT112), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n537) );
  INV_X1 U599 ( .A(n539), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n535), .A2(n563), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  NOR2_X1 U603 ( .A1(n554), .A2(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(KEYINPUT114), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  OR2_X1 U607 ( .A1(n567), .A2(n543), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n569), .A2(n553), .ZN(n545) );
  XNOR2_X1 U609 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  NOR2_X1 U612 ( .A1(n553), .A2(n559), .ZN(n550) );
  XOR2_X1 U613 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n548) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  INV_X1 U617 ( .A(n551), .ZN(n579) );
  NOR2_X1 U618 ( .A1(n579), .A2(n553), .ZN(n552) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NOR2_X1 U622 ( .A1(n569), .A2(n562), .ZN(n556) );
  XOR2_X1 U623 ( .A(G169GAT), .B(n556), .Z(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n561) );
  NOR2_X1 U627 ( .A1(n562), .A2(n559), .ZN(n560) );
  XOR2_X1 U628 ( .A(n561), .B(n560), .Z(G1349GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT121), .Z(n566) );
  INV_X1 U630 ( .A(n562), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n584) );
  INV_X1 U634 ( .A(n584), .ZN(n578) );
  NOR2_X1 U635 ( .A1(n569), .A2(n578), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(KEYINPUT59), .B(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n578), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

