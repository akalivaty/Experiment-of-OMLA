

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X2 U552 ( .A(n534), .B(KEYINPUT65), .ZN(G160) );
  NOR2_X2 U553 ( .A1(n779), .A2(n675), .ZN(n704) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n780) );
  NOR2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XNOR2_X2 U556 ( .A(KEYINPUT66), .B(n551), .ZN(n573) );
  AND2_X1 U557 ( .A1(n823), .A2(n816), .ZN(n517) );
  AND2_X1 U558 ( .A1(n751), .A2(n750), .ZN(n518) );
  NOR2_X1 U559 ( .A1(n1022), .A2(n679), .ZN(n682) );
  INV_X1 U560 ( .A(KEYINPUT96), .ZN(n680) );
  XNOR2_X1 U561 ( .A(n681), .B(n680), .ZN(n689) );
  AND2_X1 U562 ( .A1(n736), .A2(n711), .ZN(n713) );
  INV_X1 U563 ( .A(KEYINPUT90), .ZN(n708) );
  XNOR2_X1 U564 ( .A(n709), .B(n708), .ZN(n736) );
  XNOR2_X1 U565 ( .A(KEYINPUT29), .B(KEYINPUT98), .ZN(n701) );
  XNOR2_X1 U566 ( .A(n731), .B(KEYINPUT32), .ZN(n754) );
  INV_X1 U567 ( .A(n704), .ZN(n720) );
  NAND2_X1 U568 ( .A1(G160), .A2(G40), .ZN(n779) );
  NAND2_X1 U569 ( .A1(n517), .A2(n813), .ZN(n814) );
  OR2_X1 U570 ( .A1(n815), .A2(n814), .ZN(n831) );
  XOR2_X1 U571 ( .A(KEYINPUT70), .B(n571), .Z(n1022) );
  XOR2_X2 U572 ( .A(KEYINPUT17), .B(n519), .Z(n1011) );
  NAND2_X1 U573 ( .A1(n1011), .A2(G138), .ZN(n526) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n1006) );
  NAND2_X1 U575 ( .A1(G114), .A2(n1006), .ZN(n521) );
  INV_X1 U576 ( .A(G2104), .ZN(n522) );
  AND2_X1 U577 ( .A1(n522), .A2(G2105), .ZN(n1007) );
  NAND2_X1 U578 ( .A1(G126), .A2(n1007), .ZN(n520) );
  AND2_X1 U579 ( .A1(n521), .A2(n520), .ZN(n524) );
  NOR2_X1 U580 ( .A1(G2105), .A2(n522), .ZN(n1010) );
  BUF_X1 U581 ( .A(n1010), .Z(n893) );
  NAND2_X1 U582 ( .A1(G102), .A2(n893), .ZN(n523) );
  AND2_X1 U583 ( .A1(n524), .A2(n523), .ZN(n525) );
  AND2_X1 U584 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U585 ( .A1(G137), .A2(n1011), .ZN(n533) );
  NAND2_X1 U586 ( .A1(G101), .A2(n1010), .ZN(n527) );
  XNOR2_X1 U587 ( .A(KEYINPUT23), .B(n527), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G113), .A2(n1006), .ZN(n529) );
  NAND2_X1 U589 ( .A1(G125), .A2(n1007), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U592 ( .A1(G111), .A2(n1006), .ZN(n536) );
  NAND2_X1 U593 ( .A1(G135), .A2(n1011), .ZN(n535) );
  NAND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n1007), .A2(G123), .ZN(n537) );
  XOR2_X1 U596 ( .A(KEYINPUT18), .B(n537), .Z(n538) );
  NOR2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n893), .A2(G99), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n998) );
  XNOR2_X1 U600 ( .A(G2096), .B(n998), .ZN(n542) );
  OR2_X1 U601 ( .A1(G2100), .A2(n542), .ZN(G156) );
  INV_X1 U602 ( .A(G120), .ZN(G236) );
  INV_X1 U603 ( .A(G69), .ZN(G235) );
  INV_X1 U604 ( .A(G108), .ZN(G238) );
  XOR2_X1 U605 ( .A(G543), .B(KEYINPUT0), .Z(n629) );
  NOR2_X1 U606 ( .A1(G651), .A2(n629), .ZN(n612) );
  NAND2_X1 U607 ( .A1(n612), .A2(G51), .ZN(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT75), .B(n543), .ZN(n547) );
  INV_X1 U609 ( .A(G651), .ZN(n550) );
  NOR2_X1 U610 ( .A1(G543), .A2(n550), .ZN(n544) );
  XOR2_X1 U611 ( .A(KEYINPUT1), .B(n544), .Z(n584) );
  BUF_X1 U612 ( .A(n584), .Z(n641) );
  NAND2_X1 U613 ( .A1(n641), .A2(G63), .ZN(n545) );
  XOR2_X1 U614 ( .A(KEYINPUT74), .B(n545), .Z(n546) );
  NOR2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT6), .ZN(n556) );
  NOR2_X2 U617 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U618 ( .A1(n638), .A2(G89), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n549), .B(KEYINPUT4), .ZN(n553) );
  NOR2_X1 U620 ( .A1(n629), .A2(n550), .ZN(n551) );
  NAND2_X1 U621 ( .A1(G76), .A2(n573), .ZN(n552) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(KEYINPUT5), .B(n554), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G94), .A2(G452), .ZN(n558) );
  XNOR2_X1 U628 ( .A(n558), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n559) );
  XOR2_X1 U630 ( .A(n559), .B(KEYINPUT10), .Z(n842) );
  INV_X1 U631 ( .A(n842), .ZN(G223) );
  INV_X1 U632 ( .A(G567), .ZN(n669) );
  NOR2_X1 U633 ( .A1(G223), .A2(n669), .ZN(n560) );
  XOR2_X1 U634 ( .A(KEYINPUT11), .B(n560), .Z(n561) );
  XNOR2_X1 U635 ( .A(KEYINPUT69), .B(n561), .ZN(G234) );
  INV_X1 U636 ( .A(G860), .ZN(n602) );
  NAND2_X1 U637 ( .A1(n638), .A2(G81), .ZN(n562) );
  XNOR2_X1 U638 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U639 ( .A1(G68), .A2(n573), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U641 ( .A(n565), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U642 ( .A1(G43), .A2(n612), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n584), .A2(G56), .ZN(n566) );
  XNOR2_X1 U644 ( .A(KEYINPUT14), .B(n566), .ZN(n567) );
  AND2_X1 U645 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U646 ( .A1(n570), .A2(n569), .ZN(n571) );
  OR2_X1 U647 ( .A1(n602), .A2(n1022), .ZN(n572) );
  XOR2_X1 U648 ( .A(KEYINPUT71), .B(n572), .Z(G153) );
  NAND2_X1 U649 ( .A1(G90), .A2(n638), .ZN(n575) );
  NAND2_X1 U650 ( .A1(G77), .A2(n573), .ZN(n574) );
  NAND2_X1 U651 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U652 ( .A(KEYINPUT9), .B(n576), .ZN(n580) );
  NAND2_X1 U653 ( .A1(G52), .A2(n612), .ZN(n578) );
  NAND2_X1 U654 ( .A1(G64), .A2(n641), .ZN(n577) );
  AND2_X1 U655 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n580), .A2(n579), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U658 ( .A1(n612), .A2(G54), .ZN(n582) );
  NAND2_X1 U659 ( .A1(G79), .A2(n573), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U661 ( .A(n583), .B(KEYINPUT73), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G92), .A2(n638), .ZN(n586) );
  NAND2_X1 U663 ( .A1(G66), .A2(n584), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U665 ( .A(KEYINPUT72), .B(n587), .Z(n588) );
  NAND2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U667 ( .A(n590), .B(KEYINPUT15), .ZN(n1023) );
  OR2_X1 U668 ( .A1(n1023), .A2(G868), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U670 ( .A1(G91), .A2(n638), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G53), .A2(n612), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n573), .A2(G78), .ZN(n595) );
  XOR2_X1 U674 ( .A(KEYINPUT68), .B(n595), .Z(n596) );
  NOR2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n641), .A2(G65), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(G299) );
  INV_X1 U678 ( .A(G868), .ZN(n654) );
  NOR2_X1 U679 ( .A1(G286), .A2(n654), .ZN(n601) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n603), .A2(n1023), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(n1022), .A2(G868), .ZN(n607) );
  NAND2_X1 U686 ( .A1(G868), .A2(n1023), .ZN(n605) );
  NOR2_X1 U687 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G559), .A2(n1023), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n608), .B(n1022), .ZN(n651) );
  NOR2_X1 U691 ( .A1(G860), .A2(n651), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G93), .A2(n638), .ZN(n610) );
  NAND2_X1 U693 ( .A1(G80), .A2(n573), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U695 ( .A(KEYINPUT76), .B(n611), .Z(n614) );
  NAND2_X1 U696 ( .A1(n612), .A2(G55), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U698 ( .A1(G67), .A2(n641), .ZN(n615) );
  XNOR2_X1 U699 ( .A(KEYINPUT77), .B(n615), .ZN(n616) );
  OR2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n653) );
  XOR2_X1 U701 ( .A(n618), .B(n653), .Z(G145) );
  NAND2_X1 U702 ( .A1(G86), .A2(n638), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G48), .A2(n612), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n573), .A2(G73), .ZN(n621) );
  XOR2_X1 U706 ( .A(KEYINPUT2), .B(n621), .Z(n622) );
  NOR2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n641), .A2(G61), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G49), .A2(n612), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U713 ( .A1(n641), .A2(n628), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(G288) );
  AND2_X1 U716 ( .A1(G72), .A2(n573), .ZN(n635) );
  NAND2_X1 U717 ( .A1(G85), .A2(n638), .ZN(n633) );
  NAND2_X1 U718 ( .A1(G47), .A2(n612), .ZN(n632) );
  NAND2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U720 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n641), .A2(G60), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(G290) );
  NAND2_X1 U723 ( .A1(G88), .A2(n638), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G75), .A2(n573), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n645) );
  NAND2_X1 U726 ( .A1(G50), .A2(n612), .ZN(n643) );
  NAND2_X1 U727 ( .A1(G62), .A2(n641), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(G166) );
  INV_X1 U730 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(G305), .ZN(n646) );
  XNOR2_X1 U732 ( .A(n646), .B(G288), .ZN(n647) );
  XOR2_X1 U733 ( .A(n653), .B(n647), .Z(n649) );
  XOR2_X1 U734 ( .A(G290), .B(G303), .Z(n648) );
  XNOR2_X1 U735 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U736 ( .A(G299), .B(n650), .Z(n1026) );
  XNOR2_X1 U737 ( .A(n1026), .B(n651), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n652), .A2(G868), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U740 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U745 ( .A1(n660), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U747 ( .A1(G132), .A2(G82), .ZN(n661) );
  XNOR2_X1 U748 ( .A(n661), .B(KEYINPUT78), .ZN(n662) );
  XNOR2_X1 U749 ( .A(n662), .B(KEYINPUT22), .ZN(n663) );
  NOR2_X1 U750 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U751 ( .A1(G96), .A2(n664), .ZN(n968) );
  NAND2_X1 U752 ( .A1(G2106), .A2(n968), .ZN(n665) );
  XNOR2_X1 U753 ( .A(n665), .B(KEYINPUT79), .ZN(n671) );
  NOR2_X1 U754 ( .A1(G235), .A2(G236), .ZN(n666) );
  XNOR2_X1 U755 ( .A(KEYINPUT80), .B(n666), .ZN(n667) );
  NAND2_X1 U756 ( .A1(n667), .A2(G57), .ZN(n668) );
  NOR2_X1 U757 ( .A1(G238), .A2(n668), .ZN(n970) );
  NOR2_X1 U758 ( .A1(n669), .A2(n970), .ZN(n670) );
  NOR2_X1 U759 ( .A1(n671), .A2(n670), .ZN(G319) );
  INV_X1 U760 ( .A(G319), .ZN(n673) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n672) );
  NOR2_X1 U762 ( .A1(n673), .A2(n672), .ZN(n845) );
  NAND2_X1 U763 ( .A1(n845), .A2(G36), .ZN(G176) );
  INV_X1 U764 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U765 ( .A(G1996), .B(KEYINPUT94), .ZN(n919) );
  INV_X1 U766 ( .A(n780), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n919), .A2(n704), .ZN(n676) );
  XNOR2_X1 U768 ( .A(n676), .B(KEYINPUT26), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n720), .A2(G1341), .ZN(n677) );
  NAND2_X1 U770 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U771 ( .A1(n682), .A2(n1023), .ZN(n681) );
  NAND2_X1 U772 ( .A1(n682), .A2(n1023), .ZN(n687) );
  AND2_X1 U773 ( .A1(n704), .A2(G2067), .ZN(n683) );
  XNOR2_X1 U774 ( .A(n683), .B(KEYINPUT95), .ZN(n685) );
  NAND2_X1 U775 ( .A1(n720), .A2(G1348), .ZN(n684) );
  NAND2_X1 U776 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U777 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n720), .A2(G1956), .ZN(n692) );
  NAND2_X1 U780 ( .A1(n704), .A2(G2072), .ZN(n690) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(n690), .Z(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U783 ( .A(n693), .B(KEYINPUT93), .Z(n697) );
  OR2_X1 U784 ( .A1(G299), .A2(n697), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U786 ( .A(KEYINPUT97), .B(n696), .ZN(n700) );
  NAND2_X1 U787 ( .A1(G299), .A2(n697), .ZN(n698) );
  XOR2_X1 U788 ( .A(KEYINPUT28), .B(n698), .Z(n699) );
  NOR2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U790 ( .A(n702), .B(n701), .ZN(n735) );
  INV_X1 U791 ( .A(G1961), .ZN(n985) );
  NAND2_X1 U792 ( .A1(n720), .A2(n985), .ZN(n706) );
  XOR2_X1 U793 ( .A(G2078), .B(KEYINPUT91), .Z(n703) );
  XNOR2_X1 U794 ( .A(KEYINPUT25), .B(n703), .ZN(n924) );
  NAND2_X1 U795 ( .A1(n704), .A2(n924), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n715) );
  AND2_X1 U797 ( .A1(n715), .A2(G171), .ZN(n707) );
  XOR2_X1 U798 ( .A(KEYINPUT92), .B(n707), .Z(n733) );
  NAND2_X1 U799 ( .A1(n735), .A2(n733), .ZN(n725) );
  NAND2_X2 U800 ( .A1(G8), .A2(n720), .ZN(n775) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n775), .ZN(n709) );
  INV_X1 U802 ( .A(G8), .ZN(n710) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n720), .ZN(n732) );
  NOR2_X1 U804 ( .A1(n710), .A2(n732), .ZN(n711) );
  XNOR2_X1 U805 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n712) );
  XNOR2_X1 U806 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U807 ( .A1(G168), .A2(n714), .ZN(n717) );
  NOR2_X1 U808 ( .A1(G171), .A2(n715), .ZN(n716) );
  NOR2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n719) );
  XOR2_X1 U810 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n718) );
  XNOR2_X1 U811 ( .A(n719), .B(n718), .ZN(n737) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n775), .ZN(n722) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U815 ( .A1(G303), .A2(n723), .ZN(n726) );
  AND2_X1 U816 ( .A1(n737), .A2(n726), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n730) );
  INV_X1 U818 ( .A(n726), .ZN(n727) );
  OR2_X1 U819 ( .A1(n727), .A2(G286), .ZN(n728) );
  AND2_X1 U820 ( .A1(n728), .A2(G8), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U822 ( .A1(G8), .A2(n732), .ZN(n740) );
  AND2_X1 U823 ( .A1(n733), .A2(n736), .ZN(n734) );
  NAND2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n750) );
  INV_X1 U825 ( .A(n736), .ZN(n738) );
  OR2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n749) );
  NAND2_X1 U827 ( .A1(n750), .A2(n749), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U829 ( .A1(n741), .A2(n775), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n754), .A2(n742), .ZN(n747) );
  INV_X1 U831 ( .A(n775), .ZN(n752) );
  NOR2_X1 U832 ( .A1(G2090), .A2(G303), .ZN(n743) );
  XOR2_X1 U833 ( .A(KEYINPUT101), .B(n743), .Z(n744) );
  NAND2_X1 U834 ( .A1(G8), .A2(n744), .ZN(n745) );
  OR2_X1 U835 ( .A1(n752), .A2(n745), .ZN(n746) );
  AND2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U837 ( .A(n748), .B(KEYINPUT102), .ZN(n771) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n863) );
  AND2_X1 U839 ( .A1(n749), .A2(n863), .ZN(n751) );
  AND2_X1 U840 ( .A1(n518), .A2(n752), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n759) );
  INV_X1 U842 ( .A(n863), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n764) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n764), .A2(n755), .ZN(n864) );
  OR2_X1 U846 ( .A1(n756), .A2(n864), .ZN(n757) );
  OR2_X1 U847 ( .A1(n775), .A2(n757), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n761) );
  INV_X1 U849 ( .A(KEYINPUT64), .ZN(n760) );
  XNOR2_X1 U850 ( .A(n761), .B(n760), .ZN(n763) );
  INV_X1 U851 ( .A(KEYINPUT33), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n769) );
  NAND2_X1 U853 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U854 ( .A1(n765), .A2(n775), .ZN(n767) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n853) );
  INV_X1 U856 ( .A(n853), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U860 ( .A(KEYINPUT103), .B(n772), .Z(n778) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n773) );
  XNOR2_X1 U862 ( .A(n773), .B(KEYINPUT89), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT24), .ZN(n776) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n815) );
  NOR2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n828) );
  NAND2_X1 U867 ( .A1(G104), .A2(n893), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G140), .A2(n1011), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U870 ( .A(KEYINPUT34), .B(n783), .ZN(n790) );
  XNOR2_X1 U871 ( .A(KEYINPUT35), .B(KEYINPUT82), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n1006), .A2(G116), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n1007), .A2(G128), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT81), .B(n784), .Z(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U876 ( .A(n788), .B(n787), .Z(n789) );
  NOR2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U878 ( .A(n791), .B(KEYINPUT36), .Z(n792) );
  XNOR2_X1 U879 ( .A(KEYINPUT83), .B(n792), .ZN(n1003) );
  XNOR2_X1 U880 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NOR2_X1 U881 ( .A1(n1003), .A2(n825), .ZN(n886) );
  NAND2_X1 U882 ( .A1(n828), .A2(n886), .ZN(n793) );
  XNOR2_X1 U883 ( .A(KEYINPUT84), .B(n793), .ZN(n823) );
  XOR2_X1 U884 ( .A(KEYINPUT86), .B(KEYINPUT38), .Z(n795) );
  NAND2_X1 U885 ( .A1(G105), .A2(n893), .ZN(n794) );
  XNOR2_X1 U886 ( .A(n795), .B(n794), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G117), .A2(n1006), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G129), .A2(n1007), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U891 ( .A(KEYINPUT87), .B(n800), .Z(n802) );
  NAND2_X1 U892 ( .A1(n1011), .A2(G141), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n1017) );
  NAND2_X1 U894 ( .A1(G1996), .A2(n1017), .ZN(n811) );
  NAND2_X1 U895 ( .A1(G119), .A2(n1007), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G131), .A2(n1011), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G95), .A2(n893), .ZN(n805) );
  XNOR2_X1 U899 ( .A(KEYINPUT85), .B(n805), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n1006), .A2(G107), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n997) );
  NAND2_X1 U903 ( .A1(G1991), .A2(n997), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U905 ( .A(KEYINPUT88), .B(n812), .ZN(n887) );
  NAND2_X1 U906 ( .A1(n887), .A2(n828), .ZN(n816) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n871) );
  NAND2_X1 U908 ( .A1(n871), .A2(n828), .ZN(n813) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n1017), .ZN(n878) );
  INV_X1 U910 ( .A(n816), .ZN(n819) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n997), .ZN(n882) );
  NOR2_X1 U913 ( .A1(n817), .A2(n882), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n820), .B(KEYINPUT104), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n878), .A2(n821), .ZN(n822) );
  XNOR2_X1 U917 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n1003), .A2(n825), .ZN(n891) );
  NAND2_X1 U920 ( .A1(n826), .A2(n891), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U922 ( .A(KEYINPUT105), .B(n829), .Z(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U924 ( .A(KEYINPUT40), .B(n832), .ZN(G329) );
  XNOR2_X1 U925 ( .A(G1341), .B(G2454), .ZN(n833) );
  XNOR2_X1 U926 ( .A(n833), .B(G2430), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(G1348), .ZN(n840) );
  XOR2_X1 U928 ( .A(G2443), .B(G2427), .Z(n836) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n835) );
  XNOR2_X1 U930 ( .A(n836), .B(n835), .ZN(n838) );
  XOR2_X1 U931 ( .A(G2451), .B(G2435), .Z(n837) );
  XNOR2_X1 U932 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U933 ( .A(n840), .B(n839), .ZN(n841) );
  NAND2_X1 U934 ( .A1(n841), .A2(G14), .ZN(n1031) );
  XOR2_X1 U935 ( .A(KEYINPUT106), .B(n1031), .Z(G401) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G188) );
  NAND2_X1 U942 ( .A1(G124), .A2(n1007), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U944 ( .A1(n1006), .A2(G112), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n852) );
  NAND2_X1 U946 ( .A1(G100), .A2(n893), .ZN(n850) );
  NAND2_X1 U947 ( .A1(G136), .A2(n1011), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U949 ( .A1(n852), .A2(n851), .ZN(G162) );
  INV_X1 U950 ( .A(G16), .ZN(n962) );
  XOR2_X1 U951 ( .A(n962), .B(KEYINPUT56), .Z(n875) );
  XNOR2_X1 U952 ( .A(G1348), .B(n1023), .ZN(n857) );
  XNOR2_X1 U953 ( .A(G1966), .B(G168), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n855), .B(KEYINPUT57), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n860) );
  XNOR2_X1 U957 ( .A(G1341), .B(n1022), .ZN(n858) );
  XNOR2_X1 U958 ( .A(KEYINPUT122), .B(n858), .ZN(n859) );
  NOR2_X1 U959 ( .A1(n860), .A2(n859), .ZN(n873) );
  XOR2_X1 U960 ( .A(G171), .B(G1961), .Z(n862) );
  XNOR2_X1 U961 ( .A(G299), .B(G1956), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n869) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n866) );
  INV_X1 U964 ( .A(G1971), .ZN(n986) );
  NOR2_X1 U965 ( .A1(G166), .A2(n986), .ZN(n865) );
  NOR2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(KEYINPUT121), .B(n867), .Z(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n874) );
  NAND2_X1 U971 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U972 ( .A(n876), .B(KEYINPUT123), .ZN(n911) );
  INV_X1 U973 ( .A(G29), .ZN(n912) );
  XOR2_X1 U974 ( .A(G2090), .B(G162), .Z(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U976 ( .A(KEYINPUT51), .B(n879), .Z(n884) );
  XNOR2_X1 U977 ( .A(G160), .B(G2084), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n880), .A2(n998), .ZN(n881) );
  NOR2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n889) );
  INV_X1 U982 ( .A(n887), .ZN(n888) );
  NAND2_X1 U983 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U984 ( .A(n890), .B(KEYINPUT115), .ZN(n892) );
  NAND2_X1 U985 ( .A1(n892), .A2(n891), .ZN(n906) );
  NAND2_X1 U986 ( .A1(G103), .A2(n893), .ZN(n895) );
  NAND2_X1 U987 ( .A1(G139), .A2(n1011), .ZN(n894) );
  NAND2_X1 U988 ( .A1(n895), .A2(n894), .ZN(n901) );
  NAND2_X1 U989 ( .A1(G115), .A2(n1006), .ZN(n897) );
  NAND2_X1 U990 ( .A1(G127), .A2(n1007), .ZN(n896) );
  NAND2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U992 ( .A(KEYINPUT113), .B(n898), .ZN(n899) );
  XNOR2_X1 U993 ( .A(KEYINPUT47), .B(n899), .ZN(n900) );
  NOR2_X1 U994 ( .A1(n901), .A2(n900), .ZN(n1002) );
  XOR2_X1 U995 ( .A(G2072), .B(n1002), .Z(n903) );
  XOR2_X1 U996 ( .A(G164), .B(G2078), .Z(n902) );
  NOR2_X1 U997 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U998 ( .A(KEYINPUT50), .B(n904), .Z(n905) );
  NOR2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1000 ( .A(KEYINPUT52), .B(n907), .Z(n908) );
  NOR2_X1 U1001 ( .A1(KEYINPUT55), .A2(n908), .ZN(n909) );
  NOR2_X1 U1002 ( .A1(n912), .A2(n909), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(n911), .A2(n910), .ZN(n938) );
  XNOR2_X1 U1004 ( .A(n912), .B(KEYINPUT120), .ZN(n936) );
  XOR2_X1 U1005 ( .A(KEYINPUT119), .B(G34), .Z(n914) );
  XNOR2_X1 U1006 ( .A(G2084), .B(KEYINPUT54), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(n914), .B(n913), .ZN(n933) );
  XNOR2_X1 U1008 ( .A(G2090), .B(G35), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(KEYINPUT116), .ZN(n930) );
  XNOR2_X1 U1010 ( .A(G2067), .B(G26), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(G33), .B(G2072), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n923) );
  XOR2_X1 U1013 ( .A(G1991), .B(G25), .Z(n918) );
  NAND2_X1 U1014 ( .A1(n918), .A2(G28), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G32), .B(n919), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(n926) );
  XOR2_X1 U1018 ( .A(G27), .B(n924), .Z(n925) );
  NOR2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1020 ( .A(n927), .B(KEYINPUT117), .Z(n928) );
  XNOR2_X1 U1021 ( .A(KEYINPUT53), .B(n928), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1023 ( .A(KEYINPUT118), .B(n931), .Z(n932) );
  NOR2_X1 U1024 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1025 ( .A(n934), .B(KEYINPUT55), .ZN(n935) );
  NAND2_X1 U1026 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1027 ( .A1(n938), .A2(n937), .ZN(n966) );
  XOR2_X1 U1028 ( .A(G5), .B(G1961), .Z(n958) );
  XOR2_X1 U1029 ( .A(G1986), .B(KEYINPUT126), .Z(n939) );
  XNOR2_X1 U1030 ( .A(G24), .B(n939), .ZN(n943) );
  XNOR2_X1 U1031 ( .A(G1976), .B(G23), .ZN(n941) );
  XOR2_X1 U1032 ( .A(n986), .B(G22), .Z(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1035 ( .A(n944), .B(KEYINPUT58), .ZN(n956) );
  XNOR2_X1 U1036 ( .A(G1956), .B(G20), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n945), .B(KEYINPUT124), .ZN(n950) );
  XNOR2_X1 U1038 ( .A(G1981), .B(G6), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G1341), .B(G19), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(n948), .B(KEYINPUT125), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT59), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n951), .B(G4), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(KEYINPUT60), .B(n954), .ZN(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(G21), .B(G1966), .ZN(n959) );
  NOR2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(KEYINPUT61), .B(n961), .ZN(n963) );
  NAND2_X1 U1052 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1053 ( .A1(n964), .A2(G11), .ZN(n965) );
  NOR2_X1 U1054 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1055 ( .A(n967), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1056 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1057 ( .A(n968), .ZN(n969) );
  NAND2_X1 U1058 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1059 ( .A(KEYINPUT107), .B(n971), .ZN(G325) );
  XOR2_X1 U1060 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U1061 ( .A(G132), .ZN(G219) );
  INV_X1 U1062 ( .A(G82), .ZN(G220) );
  INV_X1 U1063 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1064 ( .A(G2678), .B(G2078), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G2067), .B(G2084), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n974) );
  XOR2_X1 U1067 ( .A(n974), .B(KEYINPUT109), .Z(n976) );
  XNOR2_X1 U1068 ( .A(G2072), .B(KEYINPUT42), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n976), .B(n975), .ZN(n980) );
  XOR2_X1 U1070 ( .A(G2100), .B(G2096), .Z(n978) );
  XNOR2_X1 U1071 ( .A(G2090), .B(KEYINPUT43), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n978), .B(n977), .ZN(n979) );
  XOR2_X1 U1073 ( .A(n980), .B(n979), .Z(G227) );
  XOR2_X1 U1074 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n982) );
  XNOR2_X1 U1075 ( .A(G1976), .B(G1956), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n982), .B(n981), .ZN(n994) );
  XOR2_X1 U1077 ( .A(KEYINPUT112), .B(G2474), .Z(n984) );
  XNOR2_X1 U1078 ( .A(G1996), .B(G1986), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n984), .B(n983), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(n985), .B(G1966), .ZN(n988) );
  XOR2_X1 U1081 ( .A(G1991), .B(n986), .Z(n987) );
  XNOR2_X1 U1082 ( .A(n988), .B(n987), .ZN(n989) );
  XOR2_X1 U1083 ( .A(n990), .B(n989), .Z(n992) );
  XNOR2_X1 U1084 ( .A(G1981), .B(KEYINPUT110), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n992), .B(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n994), .B(n993), .ZN(G229) );
  XOR2_X1 U1087 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n996) );
  XNOR2_X1 U1088 ( .A(G164), .B(G160), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n996), .B(n995), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G162), .B(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n999), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n1001), .B(n1000), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(n1003), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(n1005), .B(n1004), .ZN(n1020) );
  NAND2_X1 U1095 ( .A1(G118), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(G130), .A2(n1007), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1016) );
  NAND2_X1 U1098 ( .A1(G106), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(G142), .A2(n1011), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(n1014), .B(KEYINPUT45), .Z(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(n1018), .B(n1017), .ZN(n1019) );
  XNOR2_X1 U1104 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(G37), .A2(n1021), .ZN(G395) );
  XOR2_X1 U1106 ( .A(G286), .B(n1022), .Z(n1025) );
  XOR2_X1 U1107 ( .A(G301), .B(n1023), .Z(n1024) );
  XNOR2_X1 U1108 ( .A(n1025), .B(n1024), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(n1027), .B(n1026), .ZN(n1028) );
  NOR2_X1 U1110 ( .A1(G37), .A2(n1028), .ZN(G397) );
  NOR2_X1 U1111 ( .A1(G227), .A2(G229), .ZN(n1030) );
  XNOR2_X1 U1112 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1030), .B(n1029), .ZN(n1033) );
  NAND2_X1 U1114 ( .A1(G319), .A2(n1031), .ZN(n1032) );
  NOR2_X1 U1115 ( .A1(n1033), .A2(n1032), .ZN(n1035) );
  NOR2_X1 U1116 ( .A1(G395), .A2(G397), .ZN(n1034) );
  NAND2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(G225) );
  INV_X1 U1118 ( .A(G225), .ZN(G308) );
  INV_X1 U1119 ( .A(G96), .ZN(G221) );
endmodule

