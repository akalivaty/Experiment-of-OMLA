//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT64), .Z(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT27), .B(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n206), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n208), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT27), .B1(new_n208), .B2(KEYINPUT66), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT67), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  INV_X1    g014(.A(G176gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n216), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(KEYINPUT26), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n207), .B(new_n212), .C1(new_n214), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT25), .B1(new_n217), .B2(KEYINPUT65), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(KEYINPUT65), .B2(new_n217), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(new_n227), .C1(new_n208), .C2(new_n205), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n226), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n225), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT25), .B1(new_n230), .B2(new_n218), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n221), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT69), .ZN(new_n234));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G134gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT68), .B1(new_n238), .B2(G127gat), .ZN(new_n239));
  INV_X1    g038(.A(G120gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G113gat), .ZN(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G120gat), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n237), .A2(new_n239), .B1(KEYINPUT1), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT1), .B1(new_n241), .B2(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n235), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n221), .B(new_n249), .C1(new_n231), .C2(new_n232), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n248), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n203), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n203), .A3(new_n253), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT32), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT33), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G71gat), .B(G99gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(G15gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G43gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(new_n259), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n256), .B(KEYINPUT32), .C1(new_n258), .C2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT34), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n254), .B2(KEYINPUT71), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n266), .B2(new_n268), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n255), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n268), .ZN(new_n274));
  INV_X1    g073(.A(new_n270), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n255), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT86), .ZN(new_n281));
  INV_X1    g080(.A(G22gat), .ZN(new_n282));
  XOR2_X1   g081(.A(G141gat), .B(G148gat), .Z(new_n283));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G155gat), .B(G162gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT73), .B1(new_n289), .B2(KEYINPUT2), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n289), .A2(KEYINPUT73), .A3(KEYINPUT2), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n283), .B(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT22), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G218gat), .ZN(new_n295));
  INV_X1    g094(.A(G211gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G211gat), .B(G218gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT29), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n304), .A2(KEYINPUT80), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n304), .B2(KEYINPUT80), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n293), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G228gat), .ZN(new_n309));
  INV_X1    g108(.A(G233gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n303), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n293), .B2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n283), .A2(new_n286), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n291), .A2(new_n290), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(new_n285), .B2(new_n287), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n306), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT81), .A3(new_n313), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n316), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n317), .B1(new_n316), .B2(new_n322), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n308), .B(new_n311), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n312), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n314), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n293), .A2(KEYINPUT3), .ZN(new_n328));
  INV_X1    g127(.A(new_n304), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n327), .B(new_n328), .C1(new_n320), .C2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n309), .B2(new_n310), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n282), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n325), .A2(new_n282), .A3(new_n331), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT79), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT31), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(G50gat), .Z(new_n339));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n333), .A2(new_n340), .A3(new_n334), .A4(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n280), .A2(new_n281), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT35), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n248), .B2(new_n293), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n320), .A2(new_n245), .A3(new_n247), .A4(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n245), .A2(new_n355), .A3(new_n247), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n245), .B2(new_n247), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n321), .B(new_n328), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n353), .A2(new_n354), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n252), .A2(new_n320), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n350), .ZN(new_n362));
  INV_X1    g161(.A(new_n359), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n248), .A2(new_n293), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n365), .A3(new_n358), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n354), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n369), .B(new_n293), .C1(new_n356), .C2(new_n357), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n361), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n248), .A2(KEYINPUT74), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n245), .A2(new_n355), .A3(new_n247), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n369), .B1(new_n374), .B2(new_n293), .ZN(new_n375));
  OAI211_X1 g174(.A(KEYINPUT78), .B(new_n363), .C1(new_n371), .C2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n362), .A2(new_n365), .A3(new_n358), .A4(KEYINPUT76), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n368), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n363), .B1(new_n371), .B2(new_n375), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT78), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n360), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT0), .ZN(new_n384));
  XNOR2_X1  g183(.A(G57gat), .B(G85gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT6), .ZN(new_n388));
  INV_X1    g187(.A(new_n386), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n360), .C1(new_n378), .C2(new_n381), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n386), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G226gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n310), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n233), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n233), .B2(new_n313), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n397), .A2(new_n398), .A3(new_n326), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n326), .B1(new_n397), .B2(new_n398), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(new_n401), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n399), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT30), .A4(new_n404), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n280), .A2(new_n393), .A3(new_n344), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n347), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n346), .A3(new_n345), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n390), .A2(new_n388), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n379), .A2(new_n380), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n376), .A3(new_n377), .A4(new_n368), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n389), .B1(new_n421), .B2(new_n360), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n392), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n413), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n344), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n273), .A2(new_n279), .A3(KEYINPUT36), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT36), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n280), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT84), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(new_n430), .A3(new_n433), .A4(new_n428), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT37), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n400), .A2(new_n401), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT37), .B1(new_n409), .B2(new_n399), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n408), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n438), .A2(KEYINPUT38), .ZN(new_n439));
  INV_X1    g238(.A(new_n405), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n438), .B2(KEYINPUT38), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n391), .A2(new_n439), .A3(new_n392), .A4(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n353), .A2(new_n358), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n363), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n293), .B1(new_n356), .B2(new_n357), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT77), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(new_n361), .A3(new_n359), .A4(new_n370), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(KEYINPUT39), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n359), .B1(new_n353), .B2(new_n358), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT39), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n386), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT40), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(new_n422), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n443), .B1(new_n457), .B2(new_n412), .ZN(new_n458));
  INV_X1    g257(.A(new_n455), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n453), .ZN(new_n460));
  AND4_X1   g259(.A1(new_n443), .A2(new_n412), .A3(new_n460), .A4(new_n387), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n344), .B(new_n442), .C1(new_n458), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n432), .A2(new_n434), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n418), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G113gat), .B(G141gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(G197gat), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT11), .B(G169gat), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n468), .B(KEYINPUT12), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G29gat), .ZN(new_n471));
  INV_X1    g270(.A(G36gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT14), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT14), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G29gat), .B2(G36gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n476), .A2(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(KEYINPUT87), .B2(new_n476), .ZN(new_n478));
  XOR2_X1   g277(.A(G43gat), .B(G50gat), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(KEYINPUT15), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n482), .A2(new_n471), .A3(new_n472), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n476), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n480), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT15), .B1(new_n479), .B2(KEYINPUT88), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n282), .A2(G15gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n262), .A2(G22gat), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT90), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT90), .B1(new_n492), .B2(new_n493), .ZN(new_n495));
  OR3_X1    g294(.A1(new_n494), .A2(new_n495), .A3(G1gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT16), .ZN(new_n497));
  INV_X1    g296(.A(G1gat), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(KEYINPUT91), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(KEYINPUT91), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n494), .B2(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G8gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n501), .B2(KEYINPUT92), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n496), .B(new_n501), .C1(KEYINPUT92), .C2(new_n503), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT93), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT93), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n491), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n481), .A2(new_n510), .A3(new_n490), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n481), .B2(new_n490), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n506), .B(new_n505), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT18), .B1(new_n515), .B2(KEYINPUT94), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(KEYINPUT94), .A3(KEYINPUT18), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n514), .B(KEYINPUT13), .Z(new_n520));
  INV_X1    g319(.A(new_n509), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n507), .A2(new_n508), .A3(new_n491), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n470), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n518), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n523), .B(new_n470), .C1(new_n525), .C2(new_n516), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n464), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(G71gat), .A2(G78gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G57gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G64gat), .ZN(new_n538));
  INV_X1    g337(.A(G64gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G57gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n535), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n536), .A2(new_n544), .A3(KEYINPUT95), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G127gat), .B(G155gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT20), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n553), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G183gat), .B(G211gat), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n549), .A2(new_n550), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n507), .A2(new_n508), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  OR2_X1    g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  INV_X1    g368(.A(G85gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(G92gat), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G92gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT8), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(KEYINPUT97), .A2(G99gat), .A3(G106gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n573), .A2(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(KEYINPUT98), .A3(new_n577), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584));
  AND2_X1   g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n568), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n583), .A2(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n572), .A2(G92gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n575), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(KEYINPUT8), .A3(new_n580), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n596), .A3(KEYINPUT99), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n588), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n589), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n589), .A2(new_n597), .A3(KEYINPUT100), .A4(new_n598), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n491), .ZN(new_n604));
  NAND3_X1  g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n511), .A2(new_n512), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n603), .ZN(new_n607));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608));
  OR2_X1    g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n608), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n609), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n609), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n536), .B(new_n544), .C1(new_n590), .C2(new_n596), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n581), .A2(new_n588), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT101), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n536), .A2(new_n544), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n590), .A2(new_n596), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n598), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n599), .A2(new_n549), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n549), .A2(new_n626), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n601), .A3(new_n602), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT103), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n620), .A2(new_n624), .B1(new_n549), .B2(new_n599), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n636), .A2(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G120gat), .B(G148gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT102), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n631), .A2(new_n632), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(new_n637), .A3(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n567), .A2(new_n617), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n530), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n393), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G1gat), .ZN(G1324gat));
  INV_X1    g452(.A(new_n650), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n413), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT42), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(KEYINPUT42), .A3(new_n656), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n659), .B(new_n660), .C1(new_n503), .C2(new_n655), .ZN(G1325gat));
  NAND2_X1  g460(.A1(new_n430), .A2(new_n428), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G15gat), .B1(new_n654), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n650), .A2(new_n262), .A3(new_n280), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(G1326gat));
  OAI21_X1  g465(.A(KEYINPUT104), .B1(new_n654), .B2(new_n344), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n650), .A2(new_n668), .A3(new_n426), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n670), .B(new_n672), .ZN(G1327gat));
  NOR3_X1   g472(.A1(new_n567), .A2(new_n617), .A3(new_n647), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n530), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n471), .A3(new_n651), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n617), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n464), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n462), .A2(new_n427), .A3(new_n428), .A4(new_n430), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n416), .A2(new_n683), .A3(new_n417), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n616), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n680), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n566), .B(KEYINPUT105), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(new_n528), .A3(new_n647), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(G29gat), .B1(new_n689), .B2(new_n393), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n677), .A2(new_n678), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n679), .A2(new_n690), .A3(new_n691), .ZN(G1328gat));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n472), .A3(new_n412), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT46), .ZN(new_n694));
  OAI21_X1  g493(.A(G36gat), .B1(new_n689), .B2(new_n413), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(KEYINPUT46), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(G1329gat));
  OAI21_X1  g496(.A(G43gat), .B1(new_n689), .B2(new_n663), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n676), .A2(new_n264), .A3(new_n280), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1330gat));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n682), .A2(new_n686), .A3(new_n426), .A4(new_n688), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G50gat), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(KEYINPUT107), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n344), .A2(G50gat), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n704), .A2(G50gat), .B1(new_n676), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n706), .B(new_n708), .ZN(G1331gat));
  NOR4_X1   g508(.A1(new_n529), .A2(new_n566), .A3(new_n616), .A4(new_n648), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n684), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n684), .A2(KEYINPUT108), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n393), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(new_n537), .ZN(G1332gat));
  INV_X1    g516(.A(new_n715), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n413), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n718), .B(new_n719), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n724), .B(new_n726), .ZN(G1333gat));
  NAND3_X1  g526(.A1(new_n718), .A2(G71gat), .A3(new_n662), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  INV_X1    g528(.A(new_n280), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n715), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(G71gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n715), .A2(new_n729), .A3(new_n730), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n728), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT50), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n737), .B(new_n728), .C1(new_n733), .C2(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n718), .A2(new_n426), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n567), .A2(new_n529), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n647), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n682), .A2(new_n686), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n393), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n684), .A2(new_n616), .A3(new_n742), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n684), .A2(KEYINPUT51), .A3(new_n616), .A4(new_n742), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n651), .A2(new_n570), .A3(new_n647), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(G1336gat));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n750), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n754), .A2(new_n574), .A3(new_n412), .A4(new_n647), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n745), .A2(new_n413), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(new_n574), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT52), .ZN(G1337gat));
  NOR2_X1   g557(.A1(new_n745), .A2(new_n663), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT112), .B(G99gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n280), .A2(new_n647), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT113), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n759), .A2(new_n760), .B1(new_n751), .B2(new_n762), .ZN(G1338gat));
  NAND4_X1  g562(.A1(new_n682), .A2(new_n686), .A3(new_n426), .A4(new_n744), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n764), .A2(G106gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n344), .A2(G106gat), .A3(new_n648), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT53), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT114), .B1(new_n751), .B2(new_n767), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n772), .A3(new_n766), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n764), .B2(G106gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n770), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n772), .B1(new_n754), .B2(new_n766), .ZN(new_n778));
  AOI211_X1 g577(.A(KEYINPUT114), .B(new_n767), .C1(new_n749), .C2(new_n750), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n776), .B(new_n770), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n769), .B1(new_n777), .B2(new_n781), .ZN(G1339gat));
  INV_X1    g581(.A(new_n687), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n643), .B1(new_n635), .B2(KEYINPUT54), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n628), .A2(new_n630), .A3(new_n633), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n603), .A2(new_n629), .B1(new_n636), .B2(new_n626), .ZN(new_n786));
  INV_X1    g585(.A(new_n632), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT54), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n631), .B2(new_n632), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(KEYINPUT117), .A3(new_n785), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n784), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT118), .B1(new_n794), .B2(KEYINPUT55), .ZN(new_n795));
  INV_X1    g594(.A(new_n646), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n794), .B2(KEYINPUT55), .ZN(new_n797));
  INV_X1    g596(.A(new_n784), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n792), .A2(KEYINPUT117), .A3(new_n785), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT117), .B1(new_n792), .B2(new_n785), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n795), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n797), .A2(new_n795), .A3(new_n804), .A4(KEYINPUT119), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n529), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n521), .A2(new_n522), .A3(new_n520), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n514), .B1(new_n509), .B2(new_n513), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n468), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n526), .A2(new_n647), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n616), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n616), .A2(new_n526), .A3(new_n812), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n807), .A2(new_n815), .A3(new_n808), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n783), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n649), .A2(new_n529), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n426), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n821), .A2(new_n651), .A3(new_n413), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n280), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n823), .A2(new_n242), .A3(new_n528), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n393), .B1(new_n818), .B2(new_n820), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n730), .A2(new_n426), .A3(new_n412), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n529), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n824), .A2(new_n829), .ZN(G1340gat));
  AOI21_X1  g629(.A(G120gat), .B1(new_n828), .B2(new_n647), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n730), .A2(new_n240), .A3(new_n648), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n822), .B2(new_n832), .ZN(G1341gat));
  OAI21_X1  g632(.A(G127gat), .B1(new_n823), .B2(new_n783), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n566), .A2(G127gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n834), .B1(new_n827), .B2(new_n835), .ZN(G1342gat));
  NOR2_X1   g635(.A1(new_n617), .A2(G134gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n828), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT120), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n828), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n823), .B2(new_n617), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n839), .A2(KEYINPUT56), .A3(new_n841), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  NOR3_X1   g646(.A1(new_n662), .A2(new_n393), .A3(new_n412), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n818), .A2(new_n820), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n849), .B2(new_n426), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n426), .A2(KEYINPUT57), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n526), .A2(new_n852), .A3(new_n647), .A4(new_n812), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n813), .A2(KEYINPUT121), .ZN(new_n854));
  XOR2_X1   g653(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n855));
  OAI22_X1  g654(.A1(new_n524), .A2(new_n527), .B1(new_n794), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n797), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n853), .B(new_n854), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n617), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n567), .B1(new_n859), .B2(new_n816), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT123), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n819), .B1(new_n860), .B2(KEYINPUT123), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n851), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n848), .B1(new_n850), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G141gat), .B1(new_n864), .B2(new_n528), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n662), .A2(new_n344), .A3(new_n412), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n825), .A2(new_n866), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n867), .A2(G141gat), .A3(new_n528), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n868), .B2(KEYINPUT124), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n865), .B(new_n868), .C1(KEYINPUT124), .C2(new_n870), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1344gat));
  AOI21_X1  g673(.A(new_n851), .B1(new_n818), .B2(new_n820), .ZN(new_n875));
  INV_X1    g674(.A(new_n805), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n858), .A2(new_n617), .B1(new_n815), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n820), .B1(new_n877), .B2(new_n567), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n878), .B2(new_n426), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n647), .B(new_n848), .C1(new_n875), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G148gat), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n647), .B(new_n848), .C1(new_n850), .C2(new_n863), .ZN(new_n882));
  INV_X1    g681(.A(G148gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(KEYINPUT59), .ZN(new_n884));
  AOI22_X1  g683(.A1(KEYINPUT59), .A2(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n867), .A2(G148gat), .A3(new_n648), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT125), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888));
  INV_X1    g687(.A(new_n886), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n882), .A2(new_n884), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n880), .B2(G148gat), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n888), .B(new_n889), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n887), .A2(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(G155gat), .B1(new_n864), .B2(new_n783), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n566), .A2(G155gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n867), .B2(new_n896), .ZN(G1346gat));
  INV_X1    g696(.A(G162gat), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n864), .A2(new_n898), .A3(new_n617), .ZN(new_n899));
  INV_X1    g698(.A(new_n867), .ZN(new_n900));
  AOI21_X1  g699(.A(G162gat), .B1(new_n900), .B2(new_n616), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(G1347gat));
  NOR3_X1   g701(.A1(new_n730), .A2(new_n651), .A3(new_n413), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n821), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n215), .A3(new_n528), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n651), .B1(new_n818), .B2(new_n820), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n730), .A2(new_n426), .A3(new_n413), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n529), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n215), .B2(new_n910), .ZN(G1348gat));
  NOR3_X1   g710(.A1(new_n904), .A2(new_n216), .A3(new_n648), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n647), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n216), .B2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(G183gat), .B1(new_n904), .B2(new_n783), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n567), .A2(new_n204), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n908), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n821), .A2(new_n616), .A3(new_n903), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(G190gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT126), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(KEYINPUT126), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(KEYINPUT61), .A3(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n908), .A2(G190gat), .A3(new_n617), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(G1351gat));
  NOR3_X1   g727(.A1(new_n662), .A2(new_n344), .A3(new_n413), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n906), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT127), .B(G197gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n529), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n875), .A2(new_n879), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n663), .A2(new_n393), .A3(new_n412), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n529), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n933), .B1(new_n938), .B2(new_n932), .ZN(G1352gat));
  OR3_X1    g738(.A1(new_n930), .A2(G204gat), .A3(new_n648), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n647), .B1(new_n875), .B2(new_n879), .ZN(new_n942));
  OAI21_X1  g741(.A(G204gat), .B1(new_n942), .B2(new_n935), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(G1353gat));
  NAND3_X1  g744(.A1(new_n931), .A2(new_n296), .A3(new_n567), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n936), .A2(new_n567), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  AOI21_X1  g749(.A(G218gat), .B1(new_n931), .B2(new_n616), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n617), .A2(new_n295), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n936), .B2(new_n952), .ZN(G1355gat));
endmodule


