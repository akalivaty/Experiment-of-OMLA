//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT15), .B1(new_n209), .B2(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(G50gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G43gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(new_n211), .B2(G43gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(G43gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n209), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n214), .A2(KEYINPUT88), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n208), .A2(new_n213), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n214), .A2(new_n221), .B1(new_n223), .B2(KEYINPUT88), .ZN(new_n224));
  INV_X1    g023(.A(G8gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(G1gat), .ZN(new_n227));
  INV_X1    g026(.A(G1gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT16), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n225), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n227), .A2(new_n225), .A3(new_n230), .ZN(new_n232));
  OAI22_X1  g031(.A1(new_n222), .A2(new_n224), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n222), .B2(new_n224), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n232), .A2(new_n231), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n214), .A2(KEYINPUT88), .A3(new_n221), .ZN(new_n239));
  INV_X1    g038(.A(new_n213), .ZN(new_n240));
  INV_X1    g039(.A(new_n208), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n221), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT88), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(new_n208), .B2(new_n213), .ZN(new_n244));
  OAI211_X1 g043(.A(KEYINPUT17), .B(new_n239), .C1(new_n242), .C2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n238), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT89), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n237), .A2(new_n248), .A3(new_n245), .A4(new_n238), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n235), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n251));
  INV_X1    g050(.A(new_n224), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n238), .A2(new_n252), .A3(new_n239), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n233), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n234), .B(KEYINPUT13), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G169gat), .B(G197gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n251), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n249), .ZN(new_n264));
  INV_X1    g063(.A(new_n235), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT90), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT18), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT90), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n263), .B1(new_n271), .B2(KEYINPUT91), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT91), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n267), .A2(new_n273), .A3(new_n268), .A4(new_n270), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n268), .B1(new_n250), .B2(new_n269), .ZN(new_n275));
  AOI211_X1 g074(.A(KEYINPUT90), .B(new_n235), .C1(new_n247), .C2(new_n249), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n256), .B(new_n251), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n262), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n272), .A2(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G127gat), .B(G134gat), .Z(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT1), .ZN(new_n281));
  INV_X1    g080(.A(G120gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G113gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT67), .B(G113gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(new_n282), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n283), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n282), .A2(G113gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n280), .B1(new_n289), .B2(KEYINPUT1), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G155gat), .B(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  INV_X1    g095(.A(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(KEYINPUT75), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G148gat), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G141gat), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n302), .A2(new_n304), .B1(KEYINPUT2), .B2(new_n299), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n295), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n305), .A2(new_n293), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n306), .B2(new_n307), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n292), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n312), .B2(new_n311), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(new_n292), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT80), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT4), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(KEYINPUT80), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n314), .B(new_n317), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n318), .B1(new_n320), .B2(new_n316), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n314), .B(new_n326), .C1(new_n320), .C2(new_n318), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n310), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n291), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n318), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n331), .B2(new_n316), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(KEYINPUT77), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT77), .B1(new_n327), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n325), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(KEYINPUT79), .ZN(new_n338));
  XOR2_X1   g137(.A(G57gat), .B(G85gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  OAI21_X1  g141(.A(KEYINPUT81), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n335), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n333), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346));
  INV_X1    g145(.A(new_n342), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n325), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n336), .A2(new_n342), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT6), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n343), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT6), .A3(new_n342), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(G183gat), .A3(G190gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT24), .ZN(new_n361));
  NOR2_X1   g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  OAI221_X1 g161(.A(new_n358), .B1(new_n359), .B2(KEYINPUT23), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(KEYINPUT23), .ZN(new_n364));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n356), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT64), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n366), .A2(KEYINPUT65), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(new_n363), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n356), .B1(new_n366), .B2(KEYINPUT65), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n365), .ZN(new_n374));
  OR3_X1    g173(.A1(new_n374), .A2(new_n359), .A3(KEYINPUT26), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n359), .A2(KEYINPUT26), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n360), .A3(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n377), .B(KEYINPUT66), .Z(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT27), .B(G183gat), .ZN(new_n379));
  INV_X1    g178(.A(G190gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT28), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n355), .B1(new_n384), .B2(KEYINPUT29), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n355), .B2(new_n384), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT73), .B(G218gat), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT22), .B1(new_n387), .B2(G211gat), .ZN(new_n388));
  XOR2_X1   g187(.A(G197gat), .B(G204gat), .Z(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G211gat), .B(G218gat), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n385), .B(new_n394), .C1(new_n355), .C2(new_n384), .ZN(new_n397));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G64gat), .ZN(new_n399));
  INV_X1    g198(.A(G92gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT74), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT74), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n396), .A2(new_n404), .A3(new_n397), .A4(new_n401), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT30), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n396), .A2(new_n397), .ZN(new_n407));
  INV_X1    g206(.A(new_n401), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n402), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n353), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n394), .A2(KEYINPUT82), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n392), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n312), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n329), .ZN(new_n419));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n415), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT83), .A3(new_n395), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n395), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n419), .A2(new_n420), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n394), .B2(new_n415), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n423), .B1(new_n311), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(G228gat), .A3(G233gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT31), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G22gat), .B(G50gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n432), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n413), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n384), .A2(new_n291), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n292), .B1(new_n373), .B2(new_n383), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n444), .A2(G227gat), .A3(G233gat), .A4(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(KEYINPUT32), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT69), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n449));
  AND3_X1   g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n446), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n443), .A2(new_n449), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(KEYINPUT32), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT70), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT70), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n446), .A2(new_n456), .A3(KEYINPUT32), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n445), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT72), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT34), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n460), .A2(KEYINPUT72), .A3(new_n461), .A4(new_n462), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n459), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n465), .A2(new_n468), .A3(new_n467), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n458), .B2(new_n452), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT36), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT71), .A3(new_n469), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(KEYINPUT71), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(new_n458), .A3(new_n452), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n403), .A2(new_n405), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n408), .B1(new_n407), .B2(KEYINPUT37), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n396), .B2(new_n397), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT38), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(KEYINPUT85), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n408), .C1(new_n407), .C2(KEYINPUT37), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n480), .B(new_n484), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n438), .B1(new_n488), .B2(new_n353), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n314), .B1(new_n323), .B2(new_n324), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n316), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n319), .A2(new_n321), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n322), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n315), .B1(new_n495), .B2(new_n314), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT39), .B1(new_n331), .B2(new_n316), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n492), .B(new_n347), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT40), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n496), .A2(new_n497), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n504), .A2(KEYINPUT40), .A3(new_n492), .A4(new_n347), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n505), .B(new_n349), .C1(new_n406), .C2(new_n411), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n440), .B(new_n479), .C1(new_n489), .C2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n470), .A2(new_n472), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n509), .A2(new_n353), .A3(new_n412), .A4(new_n438), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n411), .B(new_n406), .C1(new_n351), .C2(new_n352), .ZN(new_n512));
  AND4_X1   g311(.A1(KEYINPUT35), .A2(new_n475), .A3(new_n438), .A4(new_n477), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n279), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  INV_X1    g315(.A(G57gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G64gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(G64gat), .ZN(new_n519));
  INV_X1    g318(.A(G64gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT92), .A3(G57gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  OR2_X1    g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT9), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n523), .ZN(new_n528));
  NOR2_X1   g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G127gat), .B(G155gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT20), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n537), .B(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n238), .B1(new_n534), .B2(new_n533), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G183gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n540), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G211gat), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n543), .A2(new_n545), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G85gat), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT7), .B1(new_n549), .B2(new_n400), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(G85gat), .A3(G92gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(KEYINPUT8), .A2(new_n554), .B1(new_n549), .B2(new_n400), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G99gat), .B(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(new_n557), .A3(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n252), .B2(new_n239), .ZN(new_n562));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(KEYINPUT41), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n237), .A2(new_n245), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n568), .B2(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n548), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT94), .B1(new_n553), .B2(new_n555), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n560), .B(new_n559), .C1(new_n533), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n517), .A2(G64gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n520), .A2(G57gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT9), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n530), .A2(new_n583), .B1(new_n522), .B2(new_n526), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n556), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n560), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n557), .B1(new_n553), .B2(new_n555), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n584), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n580), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(KEYINPUT10), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(new_n561), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n578), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n578), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n580), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT95), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n577), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n515), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n353), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n228), .ZN(G1324gat));
  NOR2_X1   g413(.A1(new_n609), .A2(new_n412), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT16), .B(G8gat), .Z(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT42), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT42), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  OAI221_X1 g420(.A(new_n617), .B1(new_n225), .B2(new_n615), .C1(new_n620), .C2(new_n621), .ZN(G1325gat));
  INV_X1    g421(.A(new_n609), .ZN(new_n623));
  INV_X1    g422(.A(new_n479), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n623), .A2(G15gat), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(G15gat), .B1(new_n623), .B2(new_n509), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n626), .A2(KEYINPUT98), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(KEYINPUT98), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(G1326gat));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n438), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT43), .B(G22gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT99), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n630), .B(new_n632), .ZN(G1327gat));
  NAND3_X1  g432(.A1(new_n548), .A2(new_n576), .A3(new_n606), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n515), .A2(new_n202), .A3(new_n611), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT45), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n508), .A2(new_n514), .ZN(new_n638));
  OR2_X1    g437(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n639));
  NAND2_X1  g438(.A1(KEYINPUT100), .A2(KEYINPUT44), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n638), .A2(new_n576), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n576), .ZN(new_n642));
  INV_X1    g441(.A(new_n640), .ZN(new_n643));
  AOI211_X1 g442(.A(new_n642), .B(new_n643), .C1(new_n508), .C2(new_n514), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n548), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n646), .A2(new_n279), .A3(new_n605), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n611), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n637), .B1(new_n649), .B2(new_n202), .ZN(G1328gat));
  INV_X1    g449(.A(new_n412), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n651), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G36gat), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n515), .A2(new_n203), .A3(new_n651), .A4(new_n635), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT46), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(KEYINPUT101), .A3(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(G1329gat));
  OAI211_X1 g459(.A(new_n624), .B(new_n647), .C1(new_n641), .C2(new_n644), .ZN(new_n661));
  INV_X1    g460(.A(new_n509), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(new_n634), .A3(G43gat), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n661), .A2(G43gat), .B1(new_n515), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g464(.A(new_n439), .B(new_n647), .C1(new_n641), .C2(new_n644), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(G50gat), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n515), .A2(new_n211), .A3(new_n439), .A4(new_n635), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n667), .A2(new_n668), .B1(KEYINPUT102), .B2(KEYINPUT48), .ZN(new_n669));
  NOR2_X1   g468(.A1(KEYINPUT102), .A2(KEYINPUT48), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1331gat));
  AND3_X1   g470(.A1(new_n577), .A2(new_n279), .A3(new_n605), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n638), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n612), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n517), .ZN(G1332gat));
  INV_X1    g474(.A(new_n673), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n412), .B(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT104), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1333gat));
  INV_X1    g482(.A(G71gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n676), .B2(new_n624), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n673), .A2(G71gat), .A3(new_n662), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT105), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT105), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n687), .A2(KEYINPUT50), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT50), .B1(new_n687), .B2(new_n688), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(G1334gat));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n439), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G78gat), .ZN(G1335gat));
  INV_X1    g492(.A(new_n279), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n646), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n638), .A2(new_n576), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT51), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n642), .B1(new_n508), .B2(new_n514), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n695), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n606), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n549), .A3(new_n611), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n694), .A2(new_n646), .A3(new_n606), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n645), .A2(new_n611), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n702), .B1(new_n705), .B2(new_n549), .ZN(G1336gat));
  OAI211_X1 g505(.A(new_n651), .B(new_n703), .C1(new_n641), .C2(new_n644), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G92gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n605), .A2(new_n400), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT106), .B1(new_n678), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n412), .B(KEYINPUT103), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n711), .A2(new_n712), .A3(new_n400), .A4(new_n605), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n697), .A2(KEYINPUT108), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n699), .A2(new_n695), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n699), .B2(new_n695), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n708), .A2(KEYINPUT52), .A3(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n711), .B(new_n703), .C1(new_n641), .C2(new_n644), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G92gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n698), .A2(new_n700), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n714), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT52), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT109), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n708), .A2(KEYINPUT52), .A3(new_n720), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  AOI22_X1  g528(.A1(G92gat), .A2(new_n722), .B1(new_n724), .B2(new_n714), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(KEYINPUT52), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(G1337gat));
  INV_X1    g531(.A(G99gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n701), .A2(new_n733), .A3(new_n509), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n645), .A2(new_n624), .A3(new_n703), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(new_n733), .ZN(G1338gat));
  OAI211_X1 g536(.A(new_n439), .B(new_n703), .C1(new_n641), .C2(new_n644), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G106gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n438), .A2(G106gat), .A3(new_n606), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT110), .Z(new_n742));
  INV_X1    g541(.A(new_n700), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n699), .B2(new_n695), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n739), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n742), .B(KEYINPUT111), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n718), .B2(new_n719), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n740), .B1(new_n739), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT112), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n739), .A2(new_n740), .A3(new_n745), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n718), .A2(new_n719), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n753), .A2(new_n747), .B1(new_n738), .B2(G106gat), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n751), .B(new_n752), .C1(new_n754), .C2(new_n740), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n750), .A2(new_n755), .ZN(G1339gat));
  NOR2_X1   g555(.A1(new_n607), .A2(new_n694), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT91), .B1(new_n275), .B2(new_n276), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n251), .A2(new_n256), .A3(new_n262), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n274), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n254), .A2(new_n255), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT114), .Z(new_n763));
  AOI21_X1  g562(.A(new_n234), .B1(new_n264), .B2(new_n233), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n261), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n761), .A2(new_n605), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n580), .A2(new_n589), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT10), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n592), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n594), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n771), .A2(KEYINPUT54), .A3(new_n593), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(new_n578), .C1(new_n590), .C2(new_n592), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n772), .A2(KEYINPUT55), .A3(new_n601), .A4(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n774), .A2(new_n601), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(KEYINPUT113), .A3(new_n772), .A4(KEYINPUT55), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT55), .B1(new_n778), .B2(new_n772), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n602), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n277), .A2(new_n278), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n761), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT115), .B1(new_n766), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n761), .A2(new_n605), .A3(new_n765), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n787), .B(new_n788), .C1(new_n279), .C2(new_n783), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n789), .A3(new_n642), .ZN(new_n790));
  INV_X1    g589(.A(new_n783), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(new_n761), .A3(new_n576), .A4(new_n765), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT116), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n548), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT116), .B1(new_n790), .B2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n758), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n611), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n509), .A2(new_n438), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n797), .A2(new_n798), .A3(new_n711), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G113gat), .B1(new_n800), .B2(new_n279), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n475), .A2(new_n477), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n438), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n797), .A2(new_n803), .A3(new_n711), .ZN(new_n804));
  INV_X1    g603(.A(new_n284), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n805), .A3(new_n694), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(G1340gat));
  AOI21_X1  g606(.A(G120gat), .B1(new_n804), .B2(new_n605), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n606), .A2(new_n282), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n799), .B2(new_n809), .ZN(G1341gat));
  OAI21_X1  g609(.A(G127gat), .B1(new_n800), .B2(new_n548), .ZN(new_n811));
  INV_X1    g610(.A(G127gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n804), .A2(new_n812), .A3(new_n646), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1342gat));
  OAI21_X1  g613(.A(G134gat), .B1(new_n800), .B2(new_n642), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n790), .A2(new_n792), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n548), .A3(new_n793), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n612), .B1(new_n819), .B2(new_n758), .ZN(new_n820));
  INV_X1    g619(.A(G134gat), .ZN(new_n821));
  INV_X1    g620(.A(new_n803), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n651), .A2(new_n642), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n815), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  NAND3_X1  g626(.A1(new_n796), .A2(KEYINPUT119), .A3(new_n611), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n624), .A2(new_n438), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT119), .B1(new_n796), .B2(new_n611), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n279), .A2(G141gat), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n830), .A2(new_n831), .A3(new_n711), .A4(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT58), .B1(new_n834), .B2(KEYINPUT118), .ZN(new_n835));
  INV_X1    g634(.A(new_n829), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n820), .B2(KEYINPUT119), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n797), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n837), .A2(new_n678), .A3(new_n839), .A4(new_n832), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n796), .A2(new_n842), .A3(new_n439), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n611), .A2(new_n479), .A3(new_n678), .ZN(new_n844));
  INV_X1    g643(.A(new_n792), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n642), .B1(new_n766), .B2(new_n785), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT117), .B(new_n642), .C1(new_n766), .C2(new_n785), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n646), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n439), .B1(new_n850), .B2(new_n757), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n844), .B1(new_n851), .B2(KEYINPUT57), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n843), .A2(new_n852), .A3(new_n694), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G141gat), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n840), .A2(new_n841), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n841), .B1(new_n840), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n835), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n853), .A2(G141gat), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT120), .B1(new_n834), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n840), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n840), .A2(new_n854), .A3(new_n841), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n857), .A2(new_n864), .ZN(G1344gat));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n796), .A2(new_n439), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(new_n844), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n646), .B1(new_n846), .B2(new_n792), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n842), .B(new_n439), .C1(new_n871), .C2(new_n757), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n869), .A2(new_n605), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n867), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n867), .A2(G148gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n843), .A2(new_n852), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n605), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n837), .A2(new_n839), .ZN(new_n880));
  NOR4_X1   g679(.A1(new_n880), .A2(G148gat), .A3(new_n606), .A4(new_n711), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n866), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n711), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n303), .A3(new_n605), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(KEYINPUT121), .C1(new_n874), .C2(new_n878), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n885), .ZN(G1345gat));
  NAND3_X1  g685(.A1(new_n883), .A2(new_n296), .A3(new_n646), .ZN(new_n887));
  OAI21_X1  g686(.A(G155gat), .B1(new_n876), .B2(new_n548), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n876), .B2(new_n642), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n823), .A2(new_n297), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n880), .B2(new_n891), .ZN(G1347gat));
  AND3_X1   g691(.A1(new_n796), .A2(new_n612), .A3(new_n711), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(new_n822), .ZN(new_n894));
  INV_X1    g693(.A(G169gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n694), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT122), .Z(new_n897));
  NAND2_X1  g696(.A1(new_n612), .A2(new_n651), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n798), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n796), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n279), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n897), .A2(new_n901), .ZN(G1348gat));
  AND2_X1   g701(.A1(new_n899), .A2(new_n796), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(G176gat), .A3(new_n605), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT123), .ZN(new_n905));
  AOI21_X1  g704(.A(G176gat), .B1(new_n894), .B2(new_n605), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(G1349gat));
  NAND3_X1  g706(.A1(new_n894), .A2(new_n379), .A3(new_n646), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n900), .B2(new_n548), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G183gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n900), .A2(new_n909), .A3(new_n548), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n900), .B2(new_n642), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT61), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n894), .A2(new_n380), .A3(new_n576), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n893), .A2(new_n829), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n279), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n898), .A2(new_n624), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n869), .A2(new_n872), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n694), .A2(G197gat), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n920), .A2(G197gat), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g724(.A(new_n919), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  AOI21_X1  g726(.A(G204gat), .B1(new_n927), .B2(KEYINPUT62), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n605), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n869), .A2(new_n605), .A3(new_n872), .ZN(new_n932));
  INV_X1    g731(.A(new_n921), .ZN(new_n933));
  OAI21_X1  g732(.A(G204gat), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(G1353gat));
  OAI21_X1  g734(.A(G211gat), .B1(new_n922), .B2(new_n548), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g737(.A(KEYINPUT63), .B(G211gat), .C1(new_n922), .C2(new_n548), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(KEYINPUT127), .A3(new_n939), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n919), .A2(G211gat), .A3(new_n548), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n940), .B(new_n941), .C1(KEYINPUT127), .C2(new_n938), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n926), .B2(new_n576), .ZN(new_n943));
  INV_X1    g742(.A(new_n922), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n576), .A2(new_n387), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(G1355gat));
endmodule


