//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT91), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n206), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n213));
  NOR2_X1   g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(KEYINPUT14), .Z(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n213), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(KEYINPUT90), .ZN(new_n222));
  XOR2_X1   g021(.A(G43gat), .B(G50gat), .Z(new_n223));
  NOR2_X1   g022(.A1(KEYINPUT89), .A2(KEYINPUT15), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT89), .A2(KEYINPUT15), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT88), .A3(KEYINPUT15), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n229), .B(new_n230), .C1(new_n215), .C2(KEYINPUT90), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n221), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT17), .B(new_n221), .C1(new_n227), .C2(new_n231), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n211), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n210), .A2(new_n232), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n232), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n211), .A2(KEYINPUT92), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n210), .B2(new_n232), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n238), .A3(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n237), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n238), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n241), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G197gat), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT11), .B(G169gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT12), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n241), .A2(new_n248), .A3(new_n255), .A4(new_n249), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT82), .ZN(new_n261));
  XNOR2_X1  g060(.A(G1gat), .B(G29gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT0), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G148gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT76), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT76), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G148gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n270), .A3(G141gat), .ZN(new_n271));
  INV_X1    g070(.A(G141gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G148gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT77), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NOR2_X1   g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n275), .A2(new_n277), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n267), .A2(G141gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n273), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(KEYINPUT2), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n278), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n281), .B(KEYINPUT75), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(G127gat), .A2(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G134gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n292), .B1(new_n297), .B2(G127gat), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G113gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n302), .A3(KEYINPUT68), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT68), .B1(new_n300), .B2(new_n302), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n298), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT69), .B(G120gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n300), .B1(new_n308), .B2(new_n299), .ZN(new_n309));
  INV_X1    g108(.A(new_n292), .ZN(new_n310));
  NAND2_X1  g109(.A1(G127gat), .A2(G134gat), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT1), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n291), .A2(new_n314), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n307), .A2(KEYINPUT78), .A3(new_n313), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT78), .B1(new_n307), .B2(new_n313), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n315), .B1(new_n318), .B2(new_n291), .ZN(new_n319));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT5), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n271), .A2(new_n276), .A3(new_n273), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n276), .B1(new_n271), .B2(new_n273), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n322), .A2(new_n323), .A3(new_n282), .ZN(new_n324));
  INV_X1    g123(.A(new_n290), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT3), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n284), .A2(new_n327), .A3(new_n290), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n300), .A2(new_n302), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(new_n304), .A3(new_n303), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n334), .A2(new_n298), .B1(new_n309), .B2(new_n312), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n326), .A2(new_n328), .A3(new_n330), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n291), .B2(new_n314), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n282), .B1(new_n274), .B2(KEYINPUT77), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n340), .A2(new_n277), .B1(new_n289), .B2(new_n288), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT4), .A3(new_n335), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n337), .A2(new_n320), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n339), .A2(new_n342), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n346), .A2(KEYINPUT79), .A3(new_n320), .A4(new_n337), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n321), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n337), .A2(new_n349), .A3(new_n320), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT80), .B1(new_n339), .B2(new_n342), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n339), .A2(KEYINPUT80), .A3(new_n342), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n266), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n347), .ZN(new_n358));
  INV_X1    g157(.A(new_n321), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n354), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT6), .B1(new_n360), .B2(new_n265), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT81), .B(new_n266), .C1(new_n348), .C2(new_n354), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT6), .B(new_n266), .C1(new_n348), .C2(new_n354), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G8gat), .B(G36gat), .Z(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT73), .ZN(new_n367));
  XOR2_X1   g166(.A(G64gat), .B(G92gat), .Z(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT72), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT72), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n375), .B(new_n370), .C1(new_n371), .C2(new_n372), .ZN(new_n376));
  XNOR2_X1  g175(.A(G197gat), .B(G204gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G211gat), .B(G218gat), .Z(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n381), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G183gat), .ZN(new_n385));
  INV_X1    g184(.A(G190gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G169gat), .ZN(new_n388));
  INV_X1    g187(.A(G176gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n390), .A2(KEYINPUT26), .A3(new_n391), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n387), .B(new_n392), .C1(KEYINPUT26), .C2(new_n391), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT27), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n385), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT66), .B(G183gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n394), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT28), .B1(new_n397), .B2(new_n386), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT27), .B(G183gat), .Z(new_n399));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n399), .A2(new_n400), .A3(G190gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n393), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT24), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(G183gat), .A3(G190gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n387), .B2(new_n403), .ZN(new_n405));
  INV_X1    g204(.A(new_n396), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(G190gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT23), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n408), .A2(KEYINPUT65), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n408), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n391), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n391), .A2(KEYINPUT23), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n407), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n385), .A2(new_n386), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n411), .B1(new_n405), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n413), .A2(KEYINPUT64), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n413), .A2(KEYINPUT64), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT25), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n414), .A2(KEYINPUT25), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n402), .A2(new_n420), .B1(new_n424), .B2(new_n421), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n384), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n402), .A2(new_n420), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n421), .A2(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n383), .A3(new_n422), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n369), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n430), .A3(new_n369), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n433), .B2(KEYINPUT30), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n432), .A2(KEYINPUT74), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT74), .B1(new_n432), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n434), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n261), .B1(new_n365), .B2(new_n439), .ZN(new_n440));
  AOI211_X1 g239(.A(KEYINPUT82), .B(new_n438), .C1(new_n363), .C2(new_n364), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n383), .A2(new_n424), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n341), .B1(new_n442), .B2(new_n327), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n383), .B1(new_n328), .B2(new_n424), .ZN(new_n444));
  INV_X1    g243(.A(G228gat), .ZN(new_n445));
  INV_X1    g244(.A(G233gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G22gat), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n341), .B2(new_n327), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n383), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n328), .B2(new_n424), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n443), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n447), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n449), .B(new_n450), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n443), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n328), .A2(new_n452), .A3(new_n424), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n384), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n463), .B2(new_n454), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n448), .B1(new_n464), .B2(new_n447), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(new_n450), .ZN(new_n466));
  XNOR2_X1  g265(.A(G78gat), .B(G106gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n460), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT83), .B1(new_n465), .B2(new_n450), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n449), .B1(new_n456), .B2(new_n457), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G22gat), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n467), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n468), .B1(new_n460), .B2(new_n466), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n472), .A3(new_n467), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n427), .A2(new_n335), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n402), .A2(new_n420), .A3(new_n314), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(G227gat), .A3(G233gat), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT32), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G15gat), .B(G43gat), .Z(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n488), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n482), .B(KEYINPUT32), .C1(new_n484), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n480), .A2(new_n481), .ZN(new_n495));
  INV_X1    g294(.A(G227gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(new_n446), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n492), .B2(new_n493), .ZN(new_n502));
  OAI22_X1  g301(.A1(new_n476), .A2(new_n479), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n440), .A2(new_n441), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  INV_X1    g304(.A(new_n320), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n327), .B1(new_n284), .B2(new_n290), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n507), .A2(new_n316), .A3(new_n317), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n508), .B2(new_n328), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT79), .B1(new_n509), .B2(new_n346), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n337), .A2(new_n320), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n339), .A2(new_n342), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n511), .A2(new_n344), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n359), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n354), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n265), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n516), .A2(new_n355), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n514), .A2(new_n515), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n266), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n364), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n517), .B1(new_n361), .B2(new_n355), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n475), .B1(new_n469), .B2(new_n473), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n477), .A2(new_n478), .A3(new_n474), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n489), .A2(new_n531), .A3(new_n491), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n500), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n499), .A2(new_n492), .A3(KEYINPUT71), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n529), .A2(new_n505), .A3(new_n439), .A4(new_n535), .ZN(new_n536));
  OAI22_X1  g335(.A1(new_n504), .A2(new_n505), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n529), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n440), .B2(new_n441), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT36), .B1(new_n501), .B2(new_n502), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT36), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n533), .A2(new_n541), .A3(new_n534), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT38), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n369), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n426), .A2(new_n430), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT86), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n384), .A2(KEYINPUT86), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT37), .B1(new_n426), .B2(new_n549), .ZN(new_n550));
  OAI221_X1 g349(.A(new_n544), .B1(new_n431), .B2(new_n546), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n431), .A2(new_n546), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n545), .B1(new_n426), .B2(new_n430), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT38), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n432), .A3(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n524), .A2(new_n525), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n353), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n337), .B1(new_n557), .B2(new_n351), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n506), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT39), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n319), .B2(new_n320), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n560), .A3(new_n506), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n265), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT40), .A4(new_n265), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n566), .A2(new_n438), .A3(new_n355), .A4(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(new_n476), .B2(new_n479), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n539), .B(new_n543), .C1(new_n556), .C2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n260), .B1(new_n537), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT94), .ZN(new_n573));
  INV_X1    g372(.A(G71gat), .ZN(new_n574));
  INV_X1    g373(.A(G78gat), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT93), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G57gat), .B(G64gat), .Z(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n573), .A2(new_n576), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n576), .B2(new_n573), .ZN(new_n581));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT95), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT9), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n572), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT96), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G99gat), .B(G106gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n596), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n592), .A2(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n593), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n598), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n607), .A3(new_n586), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n581), .A2(new_n586), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n603), .B2(new_n604), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n597), .A2(KEYINPUT103), .A3(new_n598), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n610), .A2(new_n605), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n588), .A2(new_n608), .ZN(new_n617));
  INV_X1    g416(.A(new_n606), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n609), .B2(new_n614), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n621), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n616), .B2(new_n619), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n623), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(KEYINPUT104), .A3(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n627), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n632), .B2(new_n623), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT105), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT104), .B1(new_n633), .B2(new_n627), .ZN(new_n639));
  NOR4_X1   g438(.A1(new_n632), .A2(new_n629), .A3(new_n623), .A4(new_n636), .ZN(new_n640));
  OAI211_X1 g439(.A(KEYINPUT105), .B(new_n637), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n210), .B1(new_n617), .B2(KEYINPUT21), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n645));
  NAND3_X1  g444(.A1(new_n588), .A2(new_n608), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(G231gat), .A3(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(G127gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n588), .A2(new_n608), .A3(new_n649), .A4(new_n645), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n648), .B1(new_n647), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n644), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  INV_X1    g454(.A(new_n644), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n656), .A3(new_n651), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G155gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G183gat), .B(G211gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n654), .A2(new_n657), .A3(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G232gat), .A2(G233gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(KEYINPUT41), .ZN(new_n669));
  XNOR2_X1  g468(.A(G134gat), .B(G162gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n618), .A2(new_n232), .B1(KEYINPUT41), .B2(new_n668), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n232), .A2(new_n233), .B1(new_n605), .B2(new_n599), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(KEYINPUT102), .A3(new_n235), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT102), .B1(new_n676), .B2(new_n235), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G190gat), .B(G218gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT100), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n675), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n676), .A2(new_n235), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n687), .B2(new_n677), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n681), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n674), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n688), .B2(new_n681), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n680), .A2(new_n682), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n673), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n643), .A2(KEYINPUT106), .A3(new_n666), .A4(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n641), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n666), .A2(new_n695), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n696), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n571), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n365), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g508(.A(new_n202), .B1(new_n706), .B2(new_n438), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT16), .B(G8gat), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n705), .A2(new_n439), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT42), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n712), .B2(KEYINPUT42), .ZN(G1325gat));
  AOI21_X1  g513(.A(G15gat), .B1(new_n706), .B2(new_n535), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n540), .A2(new_n542), .A3(G15gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT107), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(new_n706), .B2(new_n717), .ZN(G1326gat));
  AND2_X1   g517(.A1(new_n571), .A2(new_n538), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n704), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT43), .B(G22gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1327gat));
  AOI21_X1  g521(.A(new_n695), .B1(new_n537), .B2(new_n570), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n701), .A2(new_n666), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n260), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(G29gat), .A3(new_n365), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT45), .Z(new_n729));
  AND2_X1   g528(.A1(new_n690), .A2(new_n694), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n536), .A2(new_n526), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n365), .A2(new_n439), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT82), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n365), .A2(new_n261), .A3(new_n439), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n501), .A2(new_n502), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n528), .B2(new_n527), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n731), .B1(new_n737), .B2(KEYINPUT35), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n543), .B1(new_n556), .B2(new_n569), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n733), .A2(new_n734), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n538), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n730), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  OR2_X1    g541(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n730), .B(new_n745), .C1(new_n738), .C2(new_n741), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n726), .ZN(new_n748));
  OAI21_X1  g547(.A(G29gat), .B1(new_n748), .B2(new_n365), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n749), .ZN(G1328gat));
  NOR3_X1   g549(.A1(new_n727), .A2(G36gat), .A3(new_n439), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT46), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT109), .B1(new_n748), .B2(new_n439), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G36gat), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n748), .A2(KEYINPUT109), .A3(new_n439), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(G1329gat));
  NAND3_X1  g555(.A1(new_n540), .A2(new_n542), .A3(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(new_n535), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n727), .A2(new_n758), .ZN(new_n759));
  OAI22_X1  g558(.A1(new_n748), .A2(new_n757), .B1(new_n759), .B2(G43gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g560(.A(G50gat), .ZN(new_n762));
  INV_X1    g561(.A(new_n726), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n744), .B2(new_n746), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(new_n538), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n725), .A2(G50gat), .A3(new_n695), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n719), .A2(new_n767), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n765), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1331gat));
  NAND2_X1  g570(.A1(new_n537), .A2(new_n570), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n666), .A2(new_n260), .A3(new_n695), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n643), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n707), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g577(.A(new_n439), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n780), .B(new_n781), .Z(G1333gat));
  OAI21_X1  g581(.A(G71gat), .B1(new_n775), .B2(new_n543), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n535), .A2(new_n574), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1334gat));
  NOR2_X1   g586(.A1(new_n775), .A2(new_n529), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(new_n575), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n666), .A2(new_n259), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n643), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n744), .B2(new_n746), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795), .B2(new_n365), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n730), .B(new_n790), .C1(new_n738), .C2(new_n741), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n802), .A2(new_n590), .A3(new_n707), .A4(new_n701), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n803), .ZN(G1336gat));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n439), .B(new_n793), .C1(new_n744), .C2(new_n746), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n591), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n439), .A2(G92gat), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n723), .B2(new_n790), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n701), .B(new_n808), .C1(new_n809), .C2(new_n799), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n806), .B2(new_n591), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n811), .A3(KEYINPUT52), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI221_X1 g612(.A(new_n810), .B1(new_n805), .B2(new_n813), .C1(new_n806), .C2(new_n591), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n795), .B2(new_n543), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n758), .A2(G99gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n701), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1338gat));
  INV_X1    g618(.A(G106gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n794), .B2(new_n538), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n643), .A2(G106gat), .A3(new_n529), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT112), .Z(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n800), .B2(new_n801), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT53), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n802), .A2(new_n822), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n825), .B1(new_n828), .B2(new_n821), .ZN(G1339gat));
  INV_X1    g628(.A(new_n666), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n246), .A2(new_n247), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n254), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n258), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n638), .B2(new_n642), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n627), .B1(new_n632), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n622), .A2(KEYINPUT54), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n620), .A2(new_n621), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT55), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n635), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n259), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n730), .B1(new_n836), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n690), .A3(new_n694), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(new_n842), .A3(new_n834), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n830), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n773), .A2(new_n701), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n365), .A2(new_n438), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n538), .A2(new_n758), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n260), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n854), .A2(new_n707), .A3(new_n439), .A4(new_n736), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n259), .A2(new_n299), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT113), .Z(G1340gat));
  OAI21_X1  g661(.A(G120gat), .B1(new_n857), .B2(new_n643), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n643), .A2(new_n308), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n859), .B2(new_n864), .ZN(G1341gat));
  OAI21_X1  g664(.A(G127gat), .B1(new_n857), .B2(new_n830), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n666), .A2(new_n648), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n859), .B2(new_n867), .ZN(G1342gat));
  OR2_X1    g667(.A1(new_n695), .A2(new_n297), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n859), .A2(KEYINPUT114), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT114), .B1(new_n859), .B2(new_n869), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n857), .B2(new_n695), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n543), .A2(new_n538), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n438), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n854), .A2(new_n707), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n259), .A2(new_n272), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT58), .B1(new_n881), .B2(KEYINPUT115), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n855), .A2(new_n543), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n854), .B2(new_n538), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n834), .B1(new_n700), .B2(new_n641), .ZN(new_n887));
  AND4_X1   g686(.A1(new_n259), .A2(new_n846), .A3(new_n635), .A4(new_n841), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n695), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n850), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n666), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT57), .B(new_n538), .C1(new_n891), .C2(new_n852), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n259), .B(new_n885), .C1(new_n886), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(new_n881), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n883), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI211_X1 g696(.A(KEYINPUT116), .B(new_n881), .C1(new_n894), .C2(G141gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n882), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n891), .A2(new_n852), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n529), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n884), .B1(new_n902), .B2(new_n892), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n272), .B1(new_n903), .B2(new_n259), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT116), .B1(new_n904), .B2(new_n881), .ZN(new_n905));
  INV_X1    g704(.A(new_n882), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n895), .A2(new_n883), .A3(new_n896), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n899), .A2(new_n908), .ZN(G1344gat));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n843), .A2(new_n730), .A3(new_n910), .A4(new_n846), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT117), .B1(new_n849), .B2(new_n842), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n835), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n666), .B1(new_n913), .B2(new_n889), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n259), .B1(new_n696), .B2(new_n703), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n538), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n900), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(KEYINPUT118), .A3(new_n900), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n892), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n701), .A3(new_n885), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n268), .A2(new_n270), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n701), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n903), .B2(new_n701), .ZN(new_n926));
  OAI221_X1 g725(.A(new_n923), .B1(new_n879), .B2(new_n925), .C1(KEYINPUT59), .C2(new_n926), .ZN(G1345gat));
  NOR3_X1   g726(.A1(new_n879), .A2(G155gat), .A3(new_n830), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n903), .A2(new_n666), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(G155gat), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT119), .ZN(G1346gat));
  NOR3_X1   g730(.A1(new_n879), .A2(G162gat), .A3(new_n695), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  INV_X1    g732(.A(G162gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n934), .B1(new_n903), .B2(new_n730), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n933), .A2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n707), .A2(new_n439), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n854), .A2(new_n856), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n260), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n901), .A2(new_n707), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n438), .A3(new_n736), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n259), .A2(new_n388), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT121), .Z(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n938), .B2(new_n643), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n701), .A2(new_n389), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n941), .B2(new_n946), .ZN(G1349gat));
  NOR3_X1   g746(.A1(new_n941), .A2(new_n399), .A3(new_n830), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(KEYINPUT123), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT122), .ZN(new_n950));
  OR3_X1    g749(.A1(new_n938), .A2(new_n950), .A3(new_n830), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n938), .B2(new_n830), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n406), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT60), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT60), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n949), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n938), .B2(new_n695), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n730), .A2(new_n386), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n941), .B2(new_n961), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n937), .A2(new_n543), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n921), .A2(new_n259), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT125), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n893), .B1(new_n917), .B2(new_n918), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n963), .B1(new_n967), .B2(new_n920), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n968), .A2(new_n969), .A3(new_n259), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n970), .A3(G197gat), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n877), .A2(new_n439), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n940), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n973), .A2(G197gat), .A3(new_n260), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT124), .Z(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(new_n975), .ZN(G1352gat));
  XNOR2_X1  g775(.A(KEYINPUT126), .B(G204gat), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n973), .A2(new_n643), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT62), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n968), .A2(KEYINPUT127), .A3(new_n701), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n977), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT127), .B1(new_n968), .B2(new_n701), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n921), .A2(new_n666), .A3(new_n964), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n666), .A2(new_n371), .ZN(new_n987));
  OAI22_X1  g786(.A1(new_n985), .A2(new_n986), .B1(new_n973), .B2(new_n987), .ZN(G1354gat));
  AND2_X1   g787(.A1(new_n968), .A2(new_n730), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n730), .A2(new_n372), .ZN(new_n990));
  OAI22_X1  g789(.A1(new_n989), .A2(new_n372), .B1(new_n973), .B2(new_n990), .ZN(G1355gat));
endmodule


