

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n640), .A2(G651), .ZN(n643) );
  AND2_X2 U553 ( .A1(n529), .A2(G2104), .ZN(n895) );
  XOR2_X1 U554 ( .A(n583), .B(n582), .Z(n519) );
  NOR2_X2 U555 ( .A1(G2104), .A2(n529), .ZN(n889) );
  INV_X2 U556 ( .A(G2105), .ZN(n529) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U558 ( .A(n718), .B(n717), .ZN(n724) );
  XNOR2_X1 U559 ( .A(n686), .B(n685), .ZN(n796) );
  NAND2_X1 U560 ( .A1(G40), .A2(G160), .ZN(n686) );
  NOR2_X1 U561 ( .A1(n565), .A2(n523), .ZN(n566) );
  OR2_X1 U562 ( .A1(n810), .A2(n1019), .ZN(n520) );
  AND2_X1 U563 ( .A1(n643), .A2(G43), .ZN(n521) );
  AND2_X1 U564 ( .A1(n620), .A2(G137), .ZN(n522) );
  AND2_X1 U565 ( .A1(G126), .A2(n889), .ZN(n523) );
  AND2_X1 U566 ( .A1(n774), .A2(n773), .ZN(n524) );
  OR2_X1 U567 ( .A1(n761), .A2(n772), .ZN(n525) );
  XOR2_X1 U568 ( .A(KEYINPUT31), .B(n732), .Z(n526) );
  OR2_X1 U569 ( .A1(n688), .A2(n687), .ZN(n690) );
  AND2_X1 U570 ( .A1(n694), .A2(n693), .ZN(n696) );
  INV_X1 U571 ( .A(KEYINPUT99), .ZN(n740) );
  NAND2_X1 U572 ( .A1(n797), .A2(n796), .ZN(n699) );
  BUF_X1 U573 ( .A(n699), .Z(n734) );
  NAND2_X1 U574 ( .A1(n525), .A2(n968), .ZN(n762) );
  AND2_X1 U575 ( .A1(n811), .A2(n520), .ZN(n812) );
  INV_X1 U576 ( .A(KEYINPUT13), .ZN(n579) );
  NOR2_X1 U577 ( .A1(n581), .A2(n521), .ZN(n584) );
  NAND2_X1 U578 ( .A1(n584), .A2(n519), .ZN(n960) );
  AND2_X1 U579 ( .A1(n567), .A2(n566), .ZN(G164) );
  NAND2_X1 U580 ( .A1(G101), .A2(n895), .ZN(n527) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(n527), .Z(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT17), .B(n528), .Z(n620) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U584 ( .A1(G113), .A2(n888), .ZN(n531) );
  NAND2_X1 U585 ( .A1(G125), .A2(n889), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U587 ( .A1(n522), .A2(n532), .ZN(n533) );
  AND2_X2 U588 ( .A1(n534), .A2(n533), .ZN(G160) );
  NOR2_X2 U589 ( .A1(G543), .A2(G651), .ZN(n651) );
  NAND2_X1 U590 ( .A1(n651), .A2(G89), .ZN(n535) );
  XNOR2_X1 U591 ( .A(n535), .B(KEYINPUT4), .ZN(n537) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  INV_X1 U593 ( .A(G651), .ZN(n539) );
  NOR2_X2 U594 ( .A1(n640), .A2(n539), .ZN(n645) );
  NAND2_X1 U595 ( .A1(G76), .A2(n645), .ZN(n536) );
  NAND2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U597 ( .A(n538), .B(KEYINPUT5), .ZN(n546) );
  NOR2_X1 U598 ( .A1(n539), .A2(G543), .ZN(n540) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n540), .Z(n594) );
  INV_X1 U600 ( .A(n594), .ZN(n541) );
  INV_X1 U601 ( .A(n541), .ZN(n648) );
  NAND2_X1 U602 ( .A1(G63), .A2(n648), .ZN(n543) );
  NAND2_X1 U603 ( .A1(G51), .A2(n643), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U605 ( .A(KEYINPUT6), .B(n544), .Z(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U607 ( .A(n547), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G91), .A2(n651), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT66), .B(n548), .Z(n553) );
  NAND2_X1 U611 ( .A1(G65), .A2(n648), .ZN(n550) );
  NAND2_X1 U612 ( .A1(G53), .A2(n643), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT67), .B(n551), .Z(n552) );
  NOR2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n645), .A2(G78), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(G299) );
  NAND2_X1 U618 ( .A1(G85), .A2(n651), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G72), .A2(n645), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G60), .A2(n648), .ZN(n559) );
  NAND2_X1 U622 ( .A1(G47), .A2(n643), .ZN(n558) );
  NAND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n560) );
  OR2_X1 U624 ( .A1(n561), .A2(n560), .ZN(G290) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  INV_X1 U628 ( .A(G82), .ZN(G220) );
  NAND2_X1 U629 ( .A1(n620), .A2(G138), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT82), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G102), .A2(n895), .ZN(n564) );
  NAND2_X1 U632 ( .A1(G114), .A2(n888), .ZN(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U634 ( .A1(G88), .A2(n651), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G75), .A2(n645), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G62), .A2(n648), .ZN(n571) );
  NAND2_X1 U638 ( .A1(G50), .A2(n643), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(G166) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n832) );
  NAND2_X1 U644 ( .A1(n832), .A2(G567), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U646 ( .A1(n651), .A2(G81), .ZN(n576) );
  XNOR2_X1 U647 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U648 ( .A1(G68), .A2(n645), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n583) );
  NAND2_X1 U652 ( .A1(G56), .A2(n648), .ZN(n582) );
  INV_X1 U653 ( .A(G860), .ZN(n611) );
  OR2_X1 U654 ( .A1(n960), .A2(n611), .ZN(G153) );
  NAND2_X1 U655 ( .A1(G90), .A2(n651), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G77), .A2(n645), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT9), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G64), .A2(n648), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G52), .A2(n643), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT64), .B(n590), .Z(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n593), .B(KEYINPUT65), .ZN(G171) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U667 ( .A1(n594), .A2(G66), .ZN(n595) );
  XOR2_X1 U668 ( .A(KEYINPUT69), .B(n595), .Z(n597) );
  NAND2_X1 U669 ( .A1(n651), .A2(G92), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT70), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G79), .A2(n645), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G54), .A2(n643), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X2 U676 ( .A(KEYINPUT15), .B(n603), .Z(n951) );
  OR2_X1 U677 ( .A1(n951), .A2(G868), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(G284) );
  XNOR2_X1 U679 ( .A(KEYINPUT71), .B(G868), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G286), .A2(n606), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT72), .ZN(n609) );
  NOR2_X1 U682 ( .A1(G299), .A2(G868), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT73), .B(n610), .Z(G297) );
  NAND2_X1 U685 ( .A1(n611), .A2(G559), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n612), .A2(n951), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G868), .A2(n960), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G868), .A2(n951), .ZN(n614) );
  NOR2_X1 U690 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G123), .A2(n889), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT18), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n888), .A2(G111), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G99), .A2(n895), .ZN(n622) );
  BUF_X1 U697 ( .A(n620), .Z(n893) );
  NAND2_X1 U698 ( .A1(G135), .A2(n893), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n1015) );
  XNOR2_X1 U701 ( .A(n1015), .B(G2096), .ZN(n626) );
  INV_X1 U702 ( .A(G2100), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G93), .A2(n651), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n627), .B(KEYINPUT74), .ZN(n634) );
  NAND2_X1 U706 ( .A1(G67), .A2(n648), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G80), .A2(n645), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G55), .A2(n643), .ZN(n630) );
  XNOR2_X1 U710 ( .A(KEYINPUT75), .B(n630), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n666) );
  NAND2_X1 U713 ( .A1(n951), .A2(G559), .ZN(n663) );
  XNOR2_X1 U714 ( .A(n960), .B(n663), .ZN(n635) );
  NOR2_X1 U715 ( .A1(G860), .A2(n635), .ZN(n636) );
  XOR2_X1 U716 ( .A(n666), .B(n636), .Z(G145) );
  INV_X1 U717 ( .A(G166), .ZN(G303) );
  NAND2_X1 U718 ( .A1(G49), .A2(n643), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U721 ( .A1(n648), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n640), .A2(G87), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G48), .A2(n643), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n644), .B(KEYINPUT78), .ZN(n656) );
  NAND2_X1 U726 ( .A1(G73), .A2(n645), .ZN(n646) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  XNOR2_X1 U728 ( .A(n647), .B(KEYINPUT77), .ZN(n650) );
  NAND2_X1 U729 ( .A1(G61), .A2(n648), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n651), .A2(G86), .ZN(n652) );
  XOR2_X1 U732 ( .A(KEYINPUT76), .B(n652), .Z(n653) );
  NOR2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(G305) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(G303), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n657), .B(G288), .ZN(n660) );
  XOR2_X1 U737 ( .A(n960), .B(G305), .Z(n658) );
  XNOR2_X1 U738 ( .A(n666), .B(n658), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n660), .B(n659), .ZN(n662) );
  INV_X1 U740 ( .A(G299), .ZN(n948) );
  XNOR2_X1 U741 ( .A(G290), .B(n948), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n839) );
  XOR2_X1 U743 ( .A(n839), .B(n663), .Z(n664) );
  NAND2_X1 U744 ( .A1(G868), .A2(n664), .ZN(n668) );
  INV_X1 U745 ( .A(G868), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U747 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(KEYINPUT20), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n670), .B(KEYINPUT79), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U757 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U758 ( .A1(G96), .A2(n676), .ZN(n837) );
  AND2_X1 U759 ( .A1(G2106), .A2(n837), .ZN(n681) );
  NAND2_X1 U760 ( .A1(G120), .A2(G69), .ZN(n677) );
  NOR2_X1 U761 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G108), .A2(n678), .ZN(n836) );
  NAND2_X1 U763 ( .A1(G567), .A2(n836), .ZN(n679) );
  XOR2_X1 U764 ( .A(KEYINPUT80), .B(n679), .Z(n680) );
  NOR2_X1 U765 ( .A1(n681), .A2(n680), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n921) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U768 ( .A1(n921), .A2(n682), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT81), .B(n683), .Z(n835) );
  NAND2_X1 U770 ( .A1(n835), .A2(G36), .ZN(G176) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n797) );
  INV_X1 U772 ( .A(KEYINPUT84), .ZN(n685) );
  INV_X1 U773 ( .A(G1996), .ZN(n928) );
  NOR2_X1 U774 ( .A1(n699), .A2(n928), .ZN(n688) );
  XOR2_X1 U775 ( .A(KEYINPUT26), .B(KEYINPUT92), .Z(n687) );
  NAND2_X1 U776 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U777 ( .A1(n690), .A2(n689), .ZN(n694) );
  INV_X1 U778 ( .A(n960), .ZN(n692) );
  NAND2_X1 U779 ( .A1(n699), .A2(G1341), .ZN(n691) );
  AND2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U781 ( .A1(n696), .A2(n951), .ZN(n695) );
  XNOR2_X1 U782 ( .A(n695), .B(KEYINPUT95), .ZN(n706) );
  NAND2_X1 U783 ( .A1(n696), .A2(n951), .ZN(n703) );
  INV_X1 U784 ( .A(n699), .ZN(n720) );
  NAND2_X1 U785 ( .A1(n720), .A2(G2067), .ZN(n698) );
  INV_X1 U786 ( .A(KEYINPUT93), .ZN(n697) );
  XNOR2_X1 U787 ( .A(n698), .B(n697), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n734), .A2(G1348), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U791 ( .A(n704), .B(KEYINPUT94), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n711) );
  NAND2_X1 U793 ( .A1(n720), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U794 ( .A(n707), .B(KEYINPUT27), .ZN(n709) );
  INV_X1 U795 ( .A(G1956), .ZN(n975) );
  NOR2_X1 U796 ( .A1(n975), .A2(n720), .ZN(n708) );
  NOR2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U798 ( .A1(n948), .A2(n712), .ZN(n710) );
  NAND2_X1 U799 ( .A1(n711), .A2(n710), .ZN(n716) );
  NOR2_X1 U800 ( .A1(n948), .A2(n712), .ZN(n714) );
  XNOR2_X1 U801 ( .A(KEYINPUT28), .B(KEYINPUT91), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U803 ( .A1(n716), .A2(n715), .ZN(n718) );
  XNOR2_X1 U804 ( .A(KEYINPUT29), .B(KEYINPUT96), .ZN(n717) );
  NAND2_X1 U805 ( .A1(G1961), .A2(n734), .ZN(n722) );
  XOR2_X1 U806 ( .A(G2078), .B(KEYINPUT90), .Z(n719) );
  XNOR2_X1 U807 ( .A(KEYINPUT25), .B(n719), .ZN(n935) );
  NAND2_X1 U808 ( .A1(n720), .A2(n935), .ZN(n721) );
  NAND2_X1 U809 ( .A1(n722), .A2(n721), .ZN(n729) );
  NOR2_X1 U810 ( .A1(G301), .A2(n729), .ZN(n723) );
  NOR2_X2 U811 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U812 ( .A(n725), .B(KEYINPUT97), .ZN(n733) );
  NAND2_X1 U813 ( .A1(G8), .A2(n734), .ZN(n772) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n772), .ZN(n747) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n734), .ZN(n748) );
  NOR2_X1 U816 ( .A1(n747), .A2(n748), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U819 ( .A1(G168), .A2(n728), .ZN(n731) );
  AND2_X1 U820 ( .A1(G301), .A2(n729), .ZN(n730) );
  NOR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n733), .A2(n526), .ZN(n744) );
  NAND2_X1 U823 ( .A1(n744), .A2(G286), .ZN(n739) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n772), .ZN(n736) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n737), .A2(G303), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U829 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U831 ( .A(n743), .B(KEYINPUT32), .ZN(n753) );
  BUF_X1 U832 ( .A(n744), .Z(n745) );
  INV_X1 U833 ( .A(n745), .ZN(n746) );
  NOR2_X1 U834 ( .A1(n747), .A2(n746), .ZN(n750) );
  NAND2_X1 U835 ( .A1(G8), .A2(n748), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U837 ( .A(n751), .B(KEYINPUT98), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U839 ( .A(n754), .B(KEYINPUT100), .ZN(n767) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n957) );
  NOR2_X1 U842 ( .A1(n755), .A2(n957), .ZN(n756) );
  AND2_X1 U843 ( .A1(n767), .A2(n756), .ZN(n759) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n958) );
  INV_X1 U845 ( .A(n772), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n958), .A2(n757), .ZN(n758) );
  NOR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n760), .A2(KEYINPUT33), .ZN(n763) );
  NAND2_X1 U849 ( .A1(n957), .A2(KEYINPUT33), .ZN(n761) );
  XOR2_X1 U850 ( .A(G1981), .B(G305), .Z(n968) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  INV_X1 U852 ( .A(n764), .ZN(n775) );
  NAND2_X1 U853 ( .A1(G8), .A2(G166), .ZN(n765) );
  NOR2_X1 U854 ( .A1(G2090), .A2(n765), .ZN(n766) );
  XNOR2_X1 U855 ( .A(KEYINPUT101), .B(n766), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n769), .A2(n772), .ZN(n774) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XOR2_X1 U859 ( .A(n770), .B(KEYINPUT24), .Z(n771) );
  OR2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n775), .A2(n524), .ZN(n813) );
  XNOR2_X1 U862 ( .A(G1986), .B(KEYINPUT83), .ZN(n776) );
  XNOR2_X1 U863 ( .A(n776), .B(G290), .ZN(n949) );
  NAND2_X1 U864 ( .A1(G131), .A2(n893), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G119), .A2(n889), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G95), .A2(n895), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G107), .A2(n888), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  OR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n884) );
  NAND2_X1 U871 ( .A1(G1991), .A2(n884), .ZN(n783) );
  XOR2_X1 U872 ( .A(KEYINPUT86), .B(n783), .Z(n795) );
  NAND2_X1 U873 ( .A1(G117), .A2(n888), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G129), .A2(n889), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G105), .A2(n895), .ZN(n786) );
  XNOR2_X1 U877 ( .A(n786), .B(KEYINPUT87), .ZN(n787) );
  XNOR2_X1 U878 ( .A(n787), .B(KEYINPUT38), .ZN(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n790), .B(KEYINPUT88), .ZN(n792) );
  NAND2_X1 U881 ( .A1(G141), .A2(n893), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U883 ( .A(KEYINPUT89), .B(n793), .ZN(n869) );
  NOR2_X1 U884 ( .A1(n869), .A2(n928), .ZN(n794) );
  NOR2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n1020) );
  NAND2_X1 U886 ( .A1(n949), .A2(n1020), .ZN(n799) );
  INV_X1 U887 ( .A(n796), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n798), .A2(n797), .ZN(n828) );
  NAND2_X1 U889 ( .A1(n799), .A2(n828), .ZN(n811) );
  INV_X1 U890 ( .A(n828), .ZN(n810) );
  NAND2_X1 U891 ( .A1(n889), .A2(G128), .ZN(n800) );
  XOR2_X1 U892 ( .A(KEYINPUT85), .B(n800), .Z(n802) );
  NAND2_X1 U893 ( .A1(n888), .A2(G116), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U895 ( .A(n803), .B(KEYINPUT35), .ZN(n808) );
  NAND2_X1 U896 ( .A1(G104), .A2(n895), .ZN(n805) );
  NAND2_X1 U897 ( .A1(G140), .A2(n893), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U899 ( .A(KEYINPUT34), .B(n806), .Z(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U901 ( .A(n809), .B(KEYINPUT36), .ZN(n885) );
  XOR2_X1 U902 ( .A(G2067), .B(KEYINPUT37), .Z(n824) );
  NAND2_X1 U903 ( .A1(n885), .A2(n824), .ZN(n1019) );
  NAND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n814), .B(KEYINPUT102), .ZN(n830) );
  INV_X1 U906 ( .A(n869), .ZN(n815) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n815), .ZN(n1011) );
  INV_X1 U908 ( .A(n1020), .ZN(n819) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n884), .ZN(n1016) );
  NOR2_X1 U911 ( .A1(n816), .A2(n1016), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT103), .B(n817), .Z(n818) );
  NOR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n820), .B(KEYINPUT104), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n1011), .A2(n821), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n822), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n520), .ZN(n826) );
  NOR2_X1 U918 ( .A1(n885), .A2(n824), .ZN(n825) );
  XNOR2_X1 U919 ( .A(KEYINPUT105), .B(n825), .ZN(n1008) );
  NAND2_X1 U920 ( .A1(n826), .A2(n1008), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U926 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U929 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(G171), .B(n951), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n838), .B(G286), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  NOR2_X1 U938 ( .A1(G37), .A2(n841), .ZN(G397) );
  XOR2_X1 U939 ( .A(G2100), .B(G2096), .Z(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT42), .B(G2678), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2090), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1981), .B(G1966), .Z(n851) );
  XNOR2_X1 U949 ( .A(G1991), .B(G1986), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U951 ( .A(G1976), .B(G1971), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1961), .B(G1956), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U954 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U957 ( .A(G2474), .B(n858), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n859), .B(n928), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n889), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT44), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT110), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G136), .A2(n893), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G100), .A2(n895), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G112), .A2(n888), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(KEYINPUT111), .B(n868), .Z(G162) );
  XOR2_X1 U969 ( .A(n1015), .B(G162), .Z(n871) );
  XNOR2_X1 U970 ( .A(G160), .B(n869), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n904) );
  XNOR2_X1 U972 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n882) );
  NAND2_X1 U973 ( .A1(G103), .A2(n895), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G139), .A2(n893), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n874), .B(KEYINPUT115), .ZN(n880) );
  XNOR2_X1 U977 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G115), .A2(n888), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G127), .A2(n889), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(n878), .B(n877), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n1003) );
  XNOR2_X1 U983 ( .A(n1003), .B(KEYINPUT48), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n887) );
  XNOR2_X1 U986 ( .A(G164), .B(n885), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n902) );
  NAND2_X1 U988 ( .A1(G118), .A2(n888), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U991 ( .A(KEYINPUT112), .B(n892), .ZN(n900) );
  NAND2_X1 U992 ( .A1(n893), .A2(G142), .ZN(n894) );
  XOR2_X1 U993 ( .A(KEYINPUT113), .B(n894), .Z(n897) );
  NAND2_X1 U994 ( .A1(n895), .A2(G106), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n902), .B(n901), .Z(n903) );
  XOR2_X1 U999 ( .A(n904), .B(n903), .Z(n905) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n905), .ZN(n906) );
  XOR2_X1 U1001 ( .A(KEYINPUT117), .B(n906), .Z(G395) );
  XNOR2_X1 U1002 ( .A(G2454), .B(G2451), .ZN(n915) );
  XNOR2_X1 U1003 ( .A(G2430), .B(G2446), .ZN(n913) );
  XOR2_X1 U1004 ( .A(G2435), .B(G2427), .Z(n908) );
  XNOR2_X1 U1005 ( .A(KEYINPUT106), .B(G2438), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n909), .B(G2443), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n916), .A2(G14), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(KEYINPUT107), .B(n917), .ZN(G401) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n918) );
  XOR2_X1 U1015 ( .A(KEYINPUT119), .B(n918), .Z(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(KEYINPUT49), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G397), .A2(n920), .ZN(n925) );
  NOR2_X1 U1018 ( .A1(n921), .A2(G401), .ZN(n922) );
  XOR2_X1 U1019 ( .A(KEYINPUT118), .B(n922), .Z(n923) );
  NOR2_X1 U1020 ( .A1(G395), .A2(n923), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1024 ( .A(G2067), .B(G26), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(G33), .B(G2072), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(G32), .B(n928), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n929), .A2(G28), .ZN(n932) );
  XOR2_X1 U1029 ( .A(G25), .B(G1991), .Z(n930) );
  XNOR2_X1 U1030 ( .A(KEYINPUT123), .B(n930), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(G27), .B(n935), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1035 ( .A(KEYINPUT53), .B(n938), .Z(n941) );
  XOR2_X1 U1036 ( .A(G34), .B(KEYINPUT54), .Z(n939) );
  XNOR2_X1 U1037 ( .A(G2084), .B(n939), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(G35), .B(G2090), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT55), .B(n944), .ZN(n946) );
  INV_X1 U1042 ( .A(G29), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n947), .A2(G11), .ZN(n1002) );
  XNOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .ZN(n974) );
  XNOR2_X1 U1046 ( .A(n948), .B(G1956), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n966) );
  XOR2_X1 U1048 ( .A(n951), .B(G1348), .Z(n953) );
  XOR2_X1 U1049 ( .A(G171), .B(G1961), .Z(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT124), .B(n954), .ZN(n964) );
  XNOR2_X1 U1052 ( .A(G166), .B(G1971), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n955), .B(KEYINPUT125), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(G1341), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT126), .B(n967), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(KEYINPUT57), .B(n970), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n1000) );
  INV_X1 U1066 ( .A(G16), .ZN(n998) );
  XNOR2_X1 U1067 ( .A(G20), .B(n975), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G1981), .B(G6), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .Z(n980) );
  XNOR2_X1 U1073 ( .A(G4), .B(n980), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(KEYINPUT60), .B(n983), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G21), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G1961), .B(G5), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(G23), .B(G1976), .ZN(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n991) );
  XOR2_X1 U1083 ( .A(G1986), .B(G24), .Z(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(KEYINPUT58), .B(n992), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1087 ( .A(n995), .B(KEYINPUT127), .Z(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT61), .B(n996), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1031) );
  XOR2_X1 U1092 ( .A(G164), .B(G2078), .Z(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT120), .B(n1003), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G2072), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1007), .B(KEYINPUT50), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1014) );
  XOR2_X1 U1098 ( .A(G2090), .B(G162), .Z(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1012), .B(KEYINPUT51), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1024) );
  XNOR2_X1 U1102 ( .A(G160), .B(G2084), .ZN(n1018) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1022) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT121), .B(n1025), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(KEYINPUT52), .B(n1026), .Z(n1027) );
  NOR2_X1 U1110 ( .A1(KEYINPUT55), .A2(n1027), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(KEYINPUT122), .B(n1028), .Z(n1029) );
  NAND2_X1 U1112 ( .A1(G29), .A2(n1029), .ZN(n1030) );
  NAND2_X1 U1113 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

