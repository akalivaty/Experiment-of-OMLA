//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G137), .A4(new_n463), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n464), .A2(new_n465), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NOR2_X1   g060(.A1(new_n480), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n480), .A2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(KEYINPUT69), .A2(KEYINPUT4), .A3(G138), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n470), .B2(new_n471), .ZN(new_n495));
  NAND2_X1  g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n463), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n470), .B2(new_n471), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n498), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n498), .A2(new_n503), .A3(new_n506), .A4(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n513), .A2(new_n514), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT6), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n525), .B(new_n527), .C1(new_n513), .C2(new_n514), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n523), .A2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n524), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n529), .A2(new_n545), .B1(new_n531), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n524), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n529), .A2(new_n551), .B1(new_n531), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(new_n531), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n531), .A2(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n531), .B(new_n562), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n568), .A2(KEYINPUT73), .A3(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n529), .B2(new_n571), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n519), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n572), .A2(new_n573), .B1(G651), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n570), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  OR2_X1    g155(.A1(new_n523), .A2(new_n533), .ZN(G303));
  NAND2_X1  g156(.A1(new_n568), .A2(G87), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n515), .A2(G74), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n528), .A2(G543), .ZN(new_n584));
  AOI22_X1  g159(.A1(G651), .A2(new_n583), .B1(new_n584), .B2(G49), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n519), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n584), .A2(G48), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n563), .A2(G86), .A3(new_n564), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n524), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT74), .B(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n529), .A2(new_n596), .B1(new_n531), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n568), .A2(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n519), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n584), .A2(G54), .B1(G651), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT76), .Z(G148));
  NAND2_X1  g195(.A1(new_n611), .A2(new_n618), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n472), .A2(new_n476), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n486), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n488), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(G156));
  INV_X1    g213(.A(G14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT77), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT78), .Z(new_n654));
  AOI211_X1 g229(.A(new_n639), .B(new_n654), .C1(new_n652), .C2(new_n650), .ZN(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT17), .Z(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  INV_X1    g236(.A(new_n658), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(new_n656), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n661), .C1(new_n659), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n656), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n636), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(G227));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT79), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT80), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  OR2_X1    g253(.A1(new_n671), .A2(new_n673), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n676), .A3(new_n674), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n678), .B(new_n680), .C1(new_n676), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  INV_X1    g260(.A(G1981), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G32), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n488), .A2(G129), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT87), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n486), .A2(G141), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT86), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n696));
  NAND3_X1  g271(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G105), .B2(new_n476), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n693), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n691), .B1(new_n701), .B2(new_n690), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT27), .B(G1996), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n690), .A2(G27), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G164), .B2(new_n690), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n704), .B1(G2078), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G5), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G171), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G1961), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n690), .A2(G33), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(new_n463), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n714), .B(new_n716), .C1(G139), .C2(new_n486), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(new_n690), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n711), .B1(G2072), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n710), .A2(G1961), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT31), .B(G11), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT89), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(G28), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n724), .B2(G28), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n727), .B1(new_n690), .B2(new_n635), .C1(new_n718), .C2(G2072), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n690), .B1(KEYINPUT24), .B2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(KEYINPUT24), .B2(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n484), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n708), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n708), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1966), .ZN(new_n736));
  NOR4_X1   g311(.A1(new_n721), .A2(new_n728), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n707), .B(new_n737), .C1(G2078), .C2(new_n706), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT90), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT90), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT82), .B(G16), .Z(new_n741));
  INV_X1    g316(.A(G20), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n615), .B2(new_n708), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT91), .B(G1956), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n690), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n486), .A2(G140), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n488), .A2(G128), .ZN(new_n751));
  NOR2_X1   g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  AND3_X1   g329(.A1(new_n754), .A2(KEYINPUT85), .A3(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(KEYINPUT85), .B1(new_n754), .B2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n749), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n741), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n554), .B2(new_n741), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1341), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n690), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n690), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT29), .B(G2090), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n758), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G4), .A2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT84), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n610), .B2(new_n708), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1348), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n747), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n739), .A2(new_n740), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n708), .A2(G23), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n586), .B2(new_n708), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT33), .Z(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G1976), .ZN(new_n776));
  INV_X1    g351(.A(G22), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n741), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G303), .B2(new_n741), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G6), .B(G305), .S(G16), .Z(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT32), .B(G1981), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n775), .A2(G1976), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n776), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT83), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n776), .A2(KEYINPUT83), .A3(new_n785), .A4(new_n786), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n789), .A2(new_n790), .A3(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n486), .A2(G131), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n488), .A2(G119), .ZN(new_n793));
  NOR2_X1   g368(.A1(G95), .A2(G2105), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G25), .B(new_n796), .S(G29), .Z(new_n797));
  XOR2_X1   g372(.A(KEYINPUT35), .B(G1991), .Z(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT81), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n797), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n741), .A2(G24), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n599), .B2(new_n741), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1986), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT34), .B1(new_n789), .B2(new_n790), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT36), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n808), .A2(new_n809), .A3(new_n791), .A4(new_n804), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n772), .B1(new_n807), .B2(new_n810), .ZN(G311));
  XNOR2_X1  g386(.A(G311), .B(KEYINPUT92), .ZN(G150));
  AOI22_X1  g387(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n524), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT93), .B(G55), .Z(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n529), .A2(new_n815), .B1(new_n531), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n554), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n611), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  AOI21_X1  g398(.A(G860), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT94), .ZN(new_n826));
  OAI21_X1  g401(.A(G860), .B1(new_n814), .B2(new_n817), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT95), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT96), .ZN(G145));
  XNOR2_X1  g406(.A(new_n754), .B(new_n507), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n717), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n486), .A2(G142), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n488), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(G106), .A2(G2105), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(new_n626), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n833), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n700), .B(new_n796), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n635), .B(new_n492), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G160), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(G37), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n846), .B2(new_n842), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g424(.A(new_n610), .B(G299), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT41), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(KEYINPUT41), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(KEYINPUT99), .A3(KEYINPUT41), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n621), .B(new_n819), .Z(new_n857));
  MUX2_X1   g432(.A(new_n850), .B(new_n856), .S(new_n857), .Z(new_n858));
  XNOR2_X1  g433(.A(G166), .B(new_n586), .ZN(new_n859));
  XOR2_X1   g434(.A(G305), .B(new_n599), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT42), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G868), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(G868), .B2(new_n818), .ZN(G295));
  OAI21_X1  g440(.A(new_n864), .B1(G868), .B2(new_n818), .ZN(G331));
  XNOR2_X1  g441(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G171), .B(G168), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n819), .A2(new_n869), .A3(KEYINPUT101), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n819), .B(new_n869), .Z(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n854), .A2(new_n855), .A3(new_n870), .A4(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n850), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n861), .B(KEYINPUT102), .Z(new_n878));
  AND2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n861), .A3(new_n876), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n868), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n851), .A2(new_n885), .A3(new_n853), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n851), .A2(new_n885), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n886), .A2(new_n871), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n850), .B1(new_n873), .B2(new_n870), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n883), .B1(new_n891), .B2(new_n868), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT44), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(KEYINPUT104), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n884), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(KEYINPUT43), .A3(new_n896), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n879), .A2(new_n882), .A3(new_n868), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n893), .B1(new_n899), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT105), .B(G1384), .Z(new_n902));
  AND2_X1   g477(.A1(new_n507), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n903), .B2(KEYINPUT106), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n475), .A2(new_n483), .A3(G40), .A4(new_n477), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n507), .A2(KEYINPUT106), .A3(new_n902), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G1996), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(new_n700), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n907), .B(KEYINPUT107), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n754), .B(G2067), .Z(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n701), .B2(new_n908), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n798), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n796), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n796), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1986), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n599), .B(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n907), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n924));
  INV_X1    g499(.A(G1384), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n507), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n905), .B1(new_n926), .B2(new_n901), .ZN(new_n927));
  AND3_X1   g502(.A1(KEYINPUT69), .A2(KEYINPUT4), .A3(G138), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n464), .B2(new_n465), .ZN(new_n929));
  AOI21_X1  g504(.A(G2105), .B1(new_n929), .B2(new_n496), .ZN(new_n930));
  OAI21_X1  g505(.A(G126), .B1(new_n464), .B2(new_n465), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n463), .B1(new_n931), .B2(new_n501), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT70), .B1(new_n933), .B2(new_n506), .ZN(new_n934));
  INV_X1    g509(.A(new_n510), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n925), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n927), .B1(new_n936), .B2(new_n901), .ZN(new_n937));
  INV_X1    g512(.A(G1966), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(KEYINPUT50), .ZN(new_n940));
  AOI21_X1  g515(.A(G1384), .B1(new_n933), .B2(new_n506), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n905), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n732), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(G8), .B(new_n924), .C1(new_n945), .C2(G286), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(G8), .A3(G286), .ZN(new_n947));
  INV_X1    g522(.A(G8), .ZN(new_n948));
  INV_X1    g523(.A(new_n945), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(G168), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT119), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT51), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n946), .B(new_n947), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT45), .B1(new_n511), .B2(new_n925), .ZN(new_n955));
  INV_X1    g530(.A(new_n905), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n507), .A2(new_n902), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n901), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT108), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n905), .B1(new_n903), .B2(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  AOI21_X1  g536(.A(G1384), .B1(new_n509), .B2(new_n510), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n960), .B(new_n961), .C1(KEYINPUT45), .C2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G2078), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1961), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n940), .B2(new_n943), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n942), .B1(new_n511), .B2(new_n925), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n956), .B1(KEYINPUT50), .B2(new_n926), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n972), .A2(KEYINPUT113), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n969), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G2078), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT53), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n937), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT120), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT113), .B1(new_n972), .B2(new_n973), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n943), .B(new_n970), .C1(new_n962), .C2(new_n942), .ZN(new_n982));
  AOI21_X1  g557(.A(G1961), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n983), .A2(new_n984), .A3(new_n978), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n968), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G171), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n954), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n959), .A2(new_n780), .A3(new_n963), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n962), .A2(new_n942), .ZN(new_n990));
  INV_X1    g565(.A(G2090), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n905), .B1(new_n926), .B2(KEYINPUT50), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G8), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n996));
  NAND3_X1  g571(.A1(G303), .A2(new_n996), .A3(G8), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT55), .B1(G166), .B2(new_n948), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(G303), .B2(G8), .ZN(new_n1001));
  NOR3_X1   g576(.A1(G166), .A2(KEYINPUT55), .A3(new_n948), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT110), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n997), .A2(new_n1004), .A3(new_n998), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n989), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n943), .B(new_n991), .C1(new_n962), .C2(new_n942), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT109), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n940), .A2(new_n1010), .A3(new_n991), .A4(new_n943), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(G8), .B(new_n1006), .C1(new_n1007), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n591), .A2(new_n592), .A3(new_n686), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n561), .A2(G86), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n686), .B1(new_n591), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1018), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n926), .A2(new_n905), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(new_n948), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n586), .A2(G1976), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n586), .B2(G1976), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1030), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OR3_X1    g607(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1029), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1013), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n988), .A2(new_n1000), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1013), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1034), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G288), .A2(G1976), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1024), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1023), .B1(new_n1042), .B2(new_n1016), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n949), .A2(new_n948), .A3(G286), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1000), .A2(new_n1013), .A3(new_n1034), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n945), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n999), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1035), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1038), .B(new_n1045), .C1(new_n1049), .C2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1047), .A2(new_n1048), .B1(new_n1035), .B2(new_n1052), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT112), .B1(new_n1055), .B2(new_n1044), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1035), .A2(new_n953), .A3(new_n1000), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n904), .A2(new_n906), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n903), .A2(KEYINPUT45), .ZN(new_n1060));
  INV_X1    g635(.A(new_n482), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n463), .B1(new_n1061), .B2(KEYINPUT122), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(KEYINPUT122), .B2(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(G40), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n977), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1060), .A2(new_n478), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n981), .A2(new_n982), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n969), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n968), .A2(new_n1058), .A3(G301), .A4(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1069), .B(G301), .C1(new_n964), .C2(new_n966), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT54), .B1(new_n1071), .B2(KEYINPUT123), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n987), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n968), .A2(G171), .A3(new_n1069), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n975), .A2(KEYINPUT120), .A3(new_n979), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n984), .B1(new_n983), .B2(new_n978), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n967), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1074), .B(KEYINPUT54), .C1(new_n1077), .C2(G171), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1057), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1348), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n971), .B2(new_n974), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1022), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(G2067), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(KEYINPUT114), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1348), .B1(new_n981), .B2(new_n982), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n1083), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n990), .A2(new_n992), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G299), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n570), .A2(KEYINPUT57), .A3(new_n577), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n936), .A2(new_n901), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n960), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1091), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1085), .A2(new_n1088), .A3(new_n611), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1094), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n570), .B2(new_n577), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1096), .A2(new_n960), .A3(new_n1097), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1956), .B1(new_n990), .B2(new_n992), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT115), .B1(new_n1091), .B2(new_n1098), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1103), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1100), .A2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT117), .B(KEYINPUT61), .Z(new_n1111));
  OAI21_X1  g686(.A(new_n1103), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1099), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n960), .B(new_n908), .C1(KEYINPUT45), .C2(new_n962), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT116), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1096), .A2(new_n1116), .A3(new_n908), .A4(new_n960), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n1082), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n554), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT59), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1123), .A3(new_n554), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1113), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT114), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1087), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1127));
  OAI211_X1 g702(.A(KEYINPUT60), .B(new_n610), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1105), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1091), .A2(KEYINPUT115), .A3(new_n1098), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1095), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1099), .A2(KEYINPUT61), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1133), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1109), .A2(new_n1135), .A3(KEYINPUT118), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1125), .A2(new_n1128), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1085), .A2(new_n1138), .A3(new_n1088), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n610), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1110), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1054), .A2(new_n1056), .B1(new_n1079), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1037), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1079), .A2(new_n1142), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1146), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n923), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n701), .A2(new_n912), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT126), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n909), .B(KEYINPUT46), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1155));
  XNOR2_X1  g730(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n907), .A2(new_n921), .A3(new_n599), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT48), .Z(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n920), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n754), .A2(G2067), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n914), .B2(new_n917), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT125), .Z(new_n1162));
  AOI21_X1  g737(.A(new_n1159), .B1(new_n911), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1149), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g739(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n892), .A2(new_n1166), .A3(new_n688), .A4(new_n848), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


