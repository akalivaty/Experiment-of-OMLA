

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  INV_X1 U321 ( .A(KEYINPUT112), .ZN(n380) );
  XNOR2_X1 U322 ( .A(n392), .B(n391), .ZN(n461) );
  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n391) );
  XNOR2_X1 U324 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U325 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U326 ( .A(n389), .B(n388), .ZN(n560) );
  XNOR2_X1 U327 ( .A(n452), .B(KEYINPUT120), .ZN(n473) );
  XNOR2_X1 U328 ( .A(n433), .B(KEYINPUT55), .ZN(n451) );
  XNOR2_X1 U329 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U330 ( .A(KEYINPUT45), .B(n362), .Z(n289) );
  XOR2_X1 U331 ( .A(n349), .B(n348), .Z(n290) );
  XOR2_X1 U332 ( .A(n398), .B(n366), .Z(n291) );
  INV_X1 U333 ( .A(KEYINPUT70), .ZN(n308) );
  XNOR2_X1 U334 ( .A(n309), .B(n308), .ZN(n310) );
  NOR2_X1 U335 ( .A1(n570), .A2(n384), .ZN(n385) );
  XNOR2_X1 U336 ( .A(n405), .B(n310), .ZN(n314) );
  INV_X1 U337 ( .A(n370), .ZN(n371) );
  XNOR2_X1 U338 ( .A(n318), .B(n437), .ZN(n319) );
  INV_X1 U339 ( .A(KEYINPUT79), .ZN(n356) );
  XNOR2_X1 U340 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U341 ( .A(n336), .B(n369), .ZN(n337) );
  XNOR2_X1 U342 ( .A(n374), .B(n373), .ZN(n376) );
  XNOR2_X1 U343 ( .A(n338), .B(n337), .ZN(n341) );
  INV_X1 U344 ( .A(G218GAT), .ZN(n464) );
  INV_X1 U345 ( .A(G190GAT), .ZN(n474) );
  XNOR2_X1 U346 ( .A(n378), .B(n377), .ZN(n575) );
  XOR2_X1 U347 ( .A(n450), .B(n449), .Z(n539) );
  XNOR2_X1 U348 ( .A(n464), .B(KEYINPUT62), .ZN(n465) );
  XNOR2_X1 U349 ( .A(n474), .B(KEYINPUT58), .ZN(n475) );
  XNOR2_X1 U350 ( .A(n466), .B(n465), .ZN(G1355GAT) );
  XNOR2_X1 U351 ( .A(n476), .B(n475), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n292) );
  XNOR2_X1 U353 ( .A(n292), .B(G183GAT), .ZN(n293) );
  XOR2_X1 U354 ( .A(n293), .B(KEYINPUT19), .Z(n295) );
  XNOR2_X1 U355 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n294) );
  XNOR2_X1 U356 ( .A(n295), .B(n294), .ZN(n448) );
  XOR2_X1 U357 ( .A(G169GAT), .B(G8GAT), .Z(n370) );
  XOR2_X1 U358 ( .A(KEYINPUT95), .B(n370), .Z(n297) );
  NAND2_X1 U359 ( .A1(G226GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U360 ( .A(n297), .B(n296), .ZN(n300) );
  XOR2_X1 U361 ( .A(G64GAT), .B(G92GAT), .Z(n299) );
  XNOR2_X1 U362 ( .A(G176GAT), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n317) );
  XOR2_X1 U364 ( .A(n300), .B(n317), .Z(n305) );
  XOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT21), .Z(n302) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G218GAT), .ZN(n301) );
  XNOR2_X1 U367 ( .A(n302), .B(n301), .ZN(n407) );
  XNOR2_X1 U368 ( .A(G36GAT), .B(G190GAT), .ZN(n303) );
  XOR2_X1 U369 ( .A(n303), .B(KEYINPUT76), .Z(n339) );
  XOR2_X1 U370 ( .A(n407), .B(n339), .Z(n304) );
  XNOR2_X1 U371 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U372 ( .A(n448), .B(n306), .Z(n537) );
  XOR2_X1 U373 ( .A(n537), .B(KEYINPUT118), .Z(n390) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(G78GAT), .ZN(n307) );
  XNOR2_X1 U375 ( .A(n307), .B(G148GAT), .ZN(n405) );
  NAND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n309) );
  XOR2_X1 U377 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n312) );
  XNOR2_X1 U378 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n311) );
  XNOR2_X1 U379 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U380 ( .A(n314), .B(n313), .Z(n320) );
  XOR2_X1 U381 ( .A(G57GAT), .B(KEYINPUT13), .Z(n316) );
  XNOR2_X1 U382 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n315) );
  XNOR2_X1 U383 ( .A(n316), .B(n315), .ZN(n355) );
  XNOR2_X1 U384 ( .A(n355), .B(n317), .ZN(n318) );
  XOR2_X1 U385 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XOR2_X1 U386 ( .A(G99GAT), .B(G85GAT), .Z(n323) );
  XOR2_X1 U387 ( .A(n321), .B(n323), .Z(n578) );
  XNOR2_X1 U388 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n322) );
  XNOR2_X1 U389 ( .A(n322), .B(G162GAT), .ZN(n406) );
  XNOR2_X1 U390 ( .A(n406), .B(G134GAT), .ZN(n326) );
  INV_X1 U391 ( .A(n323), .ZN(n324) );
  XNOR2_X1 U392 ( .A(n324), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U393 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U394 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n328) );
  NAND2_X1 U395 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U396 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U397 ( .A(n330), .B(n329), .Z(n338) );
  XOR2_X1 U398 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n332) );
  XNOR2_X1 U399 ( .A(G106GAT), .B(G92GAT), .ZN(n331) );
  XNOR2_X1 U400 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U401 ( .A(n333), .B(KEYINPUT9), .ZN(n336) );
  XOR2_X1 U402 ( .A(G29GAT), .B(G43GAT), .Z(n335) );
  XNOR2_X1 U403 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n334) );
  XNOR2_X1 U404 ( .A(n335), .B(n334), .ZN(n369) );
  INV_X1 U405 ( .A(n339), .ZN(n340) );
  XOR2_X1 U406 ( .A(n341), .B(n340), .Z(n472) );
  XNOR2_X1 U407 ( .A(KEYINPUT36), .B(n472), .ZN(n458) );
  XOR2_X1 U408 ( .A(KEYINPUT80), .B(KEYINPUT14), .Z(n343) );
  XNOR2_X1 U409 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n342) );
  XNOR2_X1 U410 ( .A(n343), .B(n342), .ZN(n361) );
  XOR2_X1 U411 ( .A(G155GAT), .B(G211GAT), .Z(n345) );
  XNOR2_X1 U412 ( .A(G22GAT), .B(G71GAT), .ZN(n344) );
  XNOR2_X1 U413 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U414 ( .A(KEYINPUT77), .B(G64GAT), .Z(n347) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U417 ( .A(G15GAT), .B(G1GAT), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n350), .B(KEYINPUT66), .ZN(n366) );
  XOR2_X1 U419 ( .A(G127GAT), .B(G183GAT), .Z(n352) );
  NAND2_X1 U420 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n366), .B(n353), .ZN(n354) );
  XNOR2_X1 U423 ( .A(n290), .B(n354), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n355), .B(KEYINPUT12), .ZN(n357) );
  XOR2_X1 U425 ( .A(n361), .B(n360), .Z(n582) );
  INV_X1 U426 ( .A(n582), .ZN(n490) );
  NOR2_X1 U427 ( .A1(n458), .A2(n490), .ZN(n362) );
  NOR2_X1 U428 ( .A1(n578), .A2(n289), .ZN(n363) );
  XNOR2_X1 U429 ( .A(n363), .B(KEYINPUT111), .ZN(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n365) );
  XNOR2_X1 U431 ( .A(G113GAT), .B(G197GAT), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n365), .B(n364), .ZN(n378) );
  XOR2_X1 U433 ( .A(G141GAT), .B(G22GAT), .Z(n398) );
  NAND2_X1 U434 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n291), .B(n367), .ZN(n368) );
  XOR2_X1 U436 ( .A(n368), .B(KEYINPUT67), .Z(n374) );
  XNOR2_X1 U437 ( .A(n369), .B(KEYINPUT30), .ZN(n372) );
  XNOR2_X1 U438 ( .A(G36GAT), .B(G50GAT), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n377) );
  NOR2_X1 U440 ( .A1(n379), .A2(n575), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n387) );
  INV_X1 U442 ( .A(n472), .ZN(n570) );
  XOR2_X1 U443 ( .A(KEYINPUT41), .B(n578), .Z(n467) );
  NAND2_X1 U444 ( .A1(n575), .A2(n467), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n382), .B(KEYINPUT46), .ZN(n383) );
  NAND2_X1 U446 ( .A1(n383), .A2(n490), .ZN(n384) );
  XNOR2_X1 U447 ( .A(KEYINPUT47), .B(n385), .ZN(n386) );
  NAND2_X1 U448 ( .A1(n387), .A2(n386), .ZN(n389) );
  XNOR2_X1 U449 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n388) );
  NAND2_X1 U450 ( .A1(n390), .A2(n560), .ZN(n392) );
  XOR2_X1 U451 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n394) );
  XNOR2_X1 U452 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n402) );
  XOR2_X1 U454 ( .A(KEYINPUT23), .B(G204GAT), .Z(n396) );
  XNOR2_X1 U455 ( .A(KEYINPUT91), .B(KEYINPUT88), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U457 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U458 ( .A1(G228GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n411) );
  XOR2_X1 U461 ( .A(G155GAT), .B(KEYINPUT90), .Z(n404) );
  XNOR2_X1 U462 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n420) );
  XOR2_X1 U464 ( .A(n405), .B(n420), .Z(n409) );
  XNOR2_X1 U465 ( .A(n406), .B(n407), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n484) );
  XOR2_X1 U468 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n413) );
  XNOR2_X1 U469 ( .A(G1GAT), .B(G57GAT), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n430) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G148GAT), .Z(n415) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(G120GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U474 ( .A(G29GAT), .B(G162GAT), .Z(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n426) );
  XOR2_X1 U476 ( .A(G127GAT), .B(KEYINPUT0), .Z(n419) );
  XNOR2_X1 U477 ( .A(G113GAT), .B(G134GAT), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n440) );
  XNOR2_X1 U479 ( .A(n440), .B(n420), .ZN(n424) );
  XOR2_X1 U480 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n422) );
  XNOR2_X1 U481 ( .A(KEYINPUT94), .B(KEYINPUT1), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n428) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n563) );
  INV_X1 U488 ( .A(n563), .ZN(n431) );
  NOR2_X1 U489 ( .A1(n484), .A2(n431), .ZN(n432) );
  NAND2_X1 U490 ( .A1(n461), .A2(n432), .ZN(n433) );
  XOR2_X1 U491 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n435) );
  XNOR2_X1 U492 ( .A(G15GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U494 ( .A(n436), .B(G190GAT), .Z(n439) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n444) );
  XOR2_X1 U497 ( .A(G169GAT), .B(n440), .Z(n442) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U500 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U501 ( .A(G176GAT), .B(KEYINPUT83), .Z(n446) );
  XNOR2_X1 U502 ( .A(KEYINPUT82), .B(KEYINPUT87), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U505 ( .A(n539), .ZN(n545) );
  NAND2_X1 U506 ( .A1(n451), .A2(n545), .ZN(n452) );
  INV_X1 U507 ( .A(n575), .ZN(n519) );
  NOR2_X1 U508 ( .A1(n473), .A2(n519), .ZN(n454) );
  XNOR2_X1 U509 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(G1348GAT) );
  NOR2_X1 U511 ( .A1(n473), .A2(n490), .ZN(n457) );
  XNOR2_X1 U512 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(G183GAT), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(G1350GAT) );
  XOR2_X1 U515 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n460) );
  NAND2_X1 U516 ( .A1(n484), .A2(n539), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(n477) );
  NAND2_X1 U518 ( .A1(n461), .A2(n563), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n477), .A2(n462), .ZN(n583) );
  INV_X1 U520 ( .A(n583), .ZN(n463) );
  NOR2_X1 U521 ( .A1(n458), .A2(n463), .ZN(n466) );
  INV_X1 U522 ( .A(n467), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n468), .A2(n473), .ZN(n471) );
  XNOR2_X1 U524 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(G176GAT), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n471), .B(n470), .ZN(G1349GAT) );
  NOR2_X1 U527 ( .A1(n473), .A2(n472), .ZN(n476) );
  XNOR2_X1 U528 ( .A(KEYINPUT27), .B(n537), .ZN(n485) );
  NOR2_X1 U529 ( .A1(n477), .A2(n485), .ZN(n561) );
  NOR2_X1 U530 ( .A1(n537), .A2(n539), .ZN(n478) );
  NOR2_X1 U531 ( .A1(n484), .A2(n478), .ZN(n479) );
  XOR2_X1 U532 ( .A(n479), .B(KEYINPUT98), .Z(n480) );
  XNOR2_X1 U533 ( .A(KEYINPUT25), .B(n480), .ZN(n481) );
  NOR2_X1 U534 ( .A1(n561), .A2(n481), .ZN(n482) );
  XNOR2_X1 U535 ( .A(KEYINPUT99), .B(n482), .ZN(n483) );
  NAND2_X1 U536 ( .A1(n483), .A2(n563), .ZN(n489) );
  XOR2_X1 U537 ( .A(n484), .B(KEYINPUT28), .Z(n542) );
  NOR2_X1 U538 ( .A1(n563), .A2(n485), .ZN(n486) );
  NAND2_X1 U539 ( .A1(n542), .A2(n486), .ZN(n547) );
  XOR2_X1 U540 ( .A(KEYINPUT96), .B(n547), .Z(n487) );
  NAND2_X1 U541 ( .A1(n487), .A2(n539), .ZN(n488) );
  NAND2_X1 U542 ( .A1(n489), .A2(n488), .ZN(n506) );
  NOR2_X1 U543 ( .A1(n490), .A2(n570), .ZN(n491) );
  XNOR2_X1 U544 ( .A(n491), .B(KEYINPUT81), .ZN(n492) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(n492), .Z(n493) );
  AND2_X1 U546 ( .A1(n506), .A2(n493), .ZN(n521) );
  NOR2_X1 U547 ( .A1(n578), .A2(n519), .ZN(n494) );
  XNOR2_X1 U548 ( .A(n494), .B(KEYINPUT72), .ZN(n508) );
  NAND2_X1 U549 ( .A1(n521), .A2(n508), .ZN(n495) );
  XNOR2_X1 U550 ( .A(KEYINPUT100), .B(n495), .ZN(n503) );
  NOR2_X1 U551 ( .A1(n503), .A2(n563), .ZN(n496) );
  XOR2_X1 U552 ( .A(G1GAT), .B(n496), .Z(n497) );
  XNOR2_X1 U553 ( .A(KEYINPUT34), .B(n497), .ZN(G1324GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n499) );
  NOR2_X1 U555 ( .A1(n537), .A2(n503), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U557 ( .A(G8GAT), .B(n500), .ZN(G1325GAT) );
  NOR2_X1 U558 ( .A1(n503), .A2(n539), .ZN(n502) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NOR2_X1 U561 ( .A1(n542), .A2(n503), .ZN(n504) );
  XOR2_X1 U562 ( .A(G22GAT), .B(n504), .Z(G1327GAT) );
  NOR2_X1 U563 ( .A1(n582), .A2(n458), .ZN(n505) );
  NAND2_X1 U564 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U565 ( .A(KEYINPUT37), .B(n507), .ZN(n533) );
  NAND2_X1 U566 ( .A1(n533), .A2(n508), .ZN(n510) );
  XOR2_X1 U567 ( .A(KEYINPUT38), .B(KEYINPUT103), .Z(n509) );
  XNOR2_X1 U568 ( .A(n510), .B(n509), .ZN(n516) );
  NOR2_X1 U569 ( .A1(n516), .A2(n563), .ZN(n512) );
  XNOR2_X1 U570 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  NOR2_X1 U572 ( .A1(n537), .A2(n516), .ZN(n513) );
  XOR2_X1 U573 ( .A(G36GAT), .B(n513), .Z(G1329GAT) );
  NOR2_X1 U574 ( .A1(n516), .A2(n539), .ZN(n514) );
  XOR2_X1 U575 ( .A(KEYINPUT40), .B(n514), .Z(n515) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n515), .ZN(G1330GAT) );
  NOR2_X1 U577 ( .A1(n542), .A2(n516), .ZN(n517) );
  XOR2_X1 U578 ( .A(KEYINPUT104), .B(n517), .Z(n518) );
  XNOR2_X1 U579 ( .A(G50GAT), .B(n518), .ZN(G1331GAT) );
  NAND2_X1 U580 ( .A1(n467), .A2(n519), .ZN(n520) );
  XNOR2_X1 U581 ( .A(n520), .B(KEYINPUT105), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n532), .A2(n521), .ZN(n522) );
  XNOR2_X1 U583 ( .A(n522), .B(KEYINPUT106), .ZN(n528) );
  NOR2_X1 U584 ( .A1(n528), .A2(n563), .ZN(n523) );
  XOR2_X1 U585 ( .A(KEYINPUT42), .B(n523), .Z(n524) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n524), .ZN(G1332GAT) );
  NOR2_X1 U587 ( .A1(n537), .A2(n528), .ZN(n525) );
  XOR2_X1 U588 ( .A(G64GAT), .B(n525), .Z(G1333GAT) );
  NOR2_X1 U589 ( .A1(n528), .A2(n539), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(G1334GAT) );
  XNOR2_X1 U592 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n530) );
  NOR2_X1 U593 ( .A1(n542), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G78GAT), .B(n531), .ZN(G1335GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n541) );
  NOR2_X1 U597 ( .A1(n563), .A2(n541), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(n536), .ZN(G1336GAT) );
  NOR2_X1 U601 ( .A1(n537), .A2(n541), .ZN(n538) );
  XOR2_X1 U602 ( .A(G92GAT), .B(n538), .Z(G1337GAT) );
  NOR2_X1 U603 ( .A1(n539), .A2(n541), .ZN(n540) );
  XOR2_X1 U604 ( .A(G99GAT), .B(n540), .Z(G1338GAT) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT44), .B(n543), .Z(n544) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n544), .ZN(G1339GAT) );
  XOR2_X1 U608 ( .A(G113GAT), .B(KEYINPUT113), .Z(n549) );
  NAND2_X1 U609 ( .A1(n545), .A2(n560), .ZN(n546) );
  NOR2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n557), .A2(n575), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n551) );
  XNOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT114), .B(n552), .Z(n554) );
  NAND2_X1 U617 ( .A1(n557), .A2(n467), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1341GAT) );
  NAND2_X1 U619 ( .A1(n557), .A2(n582), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT50), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G127GAT), .B(n556), .ZN(G1342GAT) );
  XOR2_X1 U622 ( .A(G134GAT), .B(KEYINPUT51), .Z(n559) );
  NAND2_X1 U623 ( .A1(n557), .A2(n570), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1343GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT117), .B(n564), .Z(n571) );
  NAND2_X1 U628 ( .A1(n575), .A2(n571), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n567) );
  NAND2_X1 U631 ( .A1(n571), .A2(n467), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G148GAT), .B(n568), .ZN(G1345GAT) );
  NAND2_X1 U634 ( .A1(n571), .A2(n582), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT59), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(n574), .Z(n577) );
  NAND2_X1 U641 ( .A1(n583), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n583), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
endmodule

