//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND3_X1  g0015(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n206), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n215), .B1(new_n217), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n210), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(new_n256), .B1(G150), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n203), .A2(G20), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n210), .A3(G1), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n209), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n262), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(G50), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n250), .B1(G33), .B2(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n269), .A2(new_n273), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G226), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT65), .B(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(G222), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(G1698), .ZN(new_n283));
  OAI221_X1 g0083(.A(new_n281), .B1(new_n226), .B2(new_n279), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n278), .B1(new_n284), .B2(new_n269), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n268), .B1(new_n285), .B2(G169), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n268), .B(KEYINPUT9), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(G190), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n295), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT3), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT3), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n280), .A2(G226), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G232), .A2(G1698), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n299), .A2(new_n205), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n269), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(G238), .A2(new_n275), .B1(new_n271), .B2(new_n273), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  INV_X1    g0116(.A(new_n314), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G179), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT14), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n319), .A3(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n262), .A2(new_n220), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT12), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n226), .B2(new_n255), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n263), .A2(G68), .A3(new_n264), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT11), .B1(new_n325), .B2(new_n251), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n317), .A2(G190), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n314), .A2(G200), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n274), .B1(new_n276), .B2(new_n227), .ZN(new_n336));
  INV_X1    g0136(.A(G41), .ZN(new_n337));
  OAI211_X1 g0137(.A(G1), .B(G13), .C1(new_n299), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n279), .A2(new_n280), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n339), .A2(new_n234), .B1(new_n206), .B2(new_n279), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n283), .A2(new_n221), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT66), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n338), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OR3_X1    g0144(.A1(new_n340), .A2(new_n343), .A3(new_n341), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n336), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n287), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n254), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n256), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n252), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n263), .A2(G77), .A3(new_n264), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(G77), .B2(new_n266), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n346), .B2(G169), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n348), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n344), .A2(new_n345), .ZN(new_n360));
  INV_X1    g0160(.A(new_n336), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n357), .B1(new_n346), .B2(G190), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n298), .A2(new_n332), .A3(new_n335), .A4(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n253), .B1(new_n209), .B2(G20), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n263), .B1(new_n262), .B2(new_n253), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n279), .A2(new_n280), .A3(G223), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G226), .A2(G1698), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n303), .A2(new_n370), .B1(new_n299), .B2(new_n222), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n269), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT69), .ZN(new_n373));
  INV_X1    g0173(.A(new_n370), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n279), .A2(new_n374), .B1(G33), .B2(G87), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n279), .A2(new_n280), .A3(G223), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n338), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n338), .A2(G232), .A3(new_n272), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n274), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n373), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n274), .A2(new_n381), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n292), .B1(new_n384), .B2(new_n377), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n279), .B2(G20), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n301), .A2(G33), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n299), .A2(KEYINPUT3), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT7), .B(new_n210), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n220), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G58), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n220), .ZN(new_n395));
  OAI21_X1  g0195(.A(G20), .B1(new_n395), .B2(new_n201), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n257), .A2(G159), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n387), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT68), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT68), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n387), .C1(new_n393), .C2(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n279), .A2(new_n388), .A3(G20), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n303), .B2(new_n210), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT67), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT67), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n393), .A2(new_n410), .A3(new_n407), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n251), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n368), .B(new_n386), .C1(new_n403), .C2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT71), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT67), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n410), .B1(new_n393), .B2(new_n407), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n252), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n400), .A3(new_n402), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n419), .A2(KEYINPUT71), .A3(new_n368), .A4(new_n386), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT17), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n368), .B1(new_n403), .B2(new_n412), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n274), .A2(new_n287), .A3(new_n381), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n373), .A2(new_n379), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT70), .ZN(new_n426));
  INV_X1    g0226(.A(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n384), .B2(new_n377), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n428), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT70), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT18), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n426), .B1(new_n425), .B2(new_n428), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n423), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n413), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n422), .A2(new_n433), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n441), .A2(KEYINPUT72), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(KEYINPUT72), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n366), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n210), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT82), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT82), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n449), .A3(new_n210), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n222), .A2(new_n205), .A3(new_n206), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n279), .A2(new_n210), .A3(G68), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT19), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n255), .B2(new_n205), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n251), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n350), .A2(new_n262), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n263), .B1(G1), .B2(new_n299), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n222), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n209), .A2(new_n270), .A3(G45), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n223), .B1(new_n463), .B2(G1), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n338), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT80), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n338), .A2(new_n467), .A3(new_n462), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n279), .A2(G244), .A3(G1698), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G116), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n339), .C2(new_n221), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n269), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G200), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT84), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n469), .B1(new_n269), .B2(new_n473), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n292), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n480), .B2(new_n460), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n475), .A2(new_n380), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n477), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n475), .A2(new_n427), .ZN(new_n485));
  XOR2_X1   g0285(.A(new_n350), .B(KEYINPUT83), .Z(new_n486));
  OAI211_X1 g0286(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n287), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n479), .A2(KEYINPUT81), .A3(new_n287), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  XOR2_X1   g0296(.A(KEYINPUT65), .B(G1698), .Z(new_n497));
  NAND3_X1  g0297(.A1(new_n300), .A2(new_n302), .A3(G244), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT4), .A4(G244), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n269), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT5), .ZN(new_n505));
  OR3_X1    g0305(.A1(new_n505), .A2(KEYINPUT77), .A3(G41), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT77), .B1(new_n505), .B2(G41), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n271), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n209), .B(G45), .C1(new_n337), .C2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT76), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n510), .B(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n337), .A2(KEYINPUT5), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n269), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n509), .A2(new_n512), .B1(G257), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(G169), .B1(new_n504), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n257), .A2(G77), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n207), .A2(new_n520), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n520), .A2(new_n522), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n205), .A2(G107), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n518), .B1(new_n527), .B2(new_n210), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT74), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n518), .C1(new_n527), .C2(new_n210), .ZN(new_n531));
  OAI21_X1  g0331(.A(G107), .B1(new_n404), .B2(new_n405), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n251), .ZN(new_n534));
  MUX2_X1   g0334(.A(new_n266), .B(new_n459), .S(G97), .Z(new_n535));
  AOI21_X1  g0335(.A(new_n517), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n503), .A2(KEYINPUT75), .A3(new_n269), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT75), .B1(new_n503), .B2(new_n269), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n512), .A2(new_n271), .A3(new_n508), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n515), .A2(G257), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n540), .A2(new_n287), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT78), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n504), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n503), .A2(KEYINPUT75), .A3(new_n269), .ZN(new_n546));
  AND4_X1   g0346(.A1(KEYINPUT78), .A2(new_n545), .A3(new_n546), .A4(new_n542), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n536), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT79), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT79), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n536), .B(new_n550), .C1(new_n543), .C2(new_n547), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n534), .A2(new_n535), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n504), .A2(new_n516), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n545), .A2(new_n546), .A3(new_n516), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n552), .B(new_n554), .C1(new_n292), .C2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n495), .A2(new_n549), .A3(new_n551), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n279), .A2(G257), .A3(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G294), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n339), .C2(new_n223), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n269), .B1(new_n515), .B2(G264), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n540), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G169), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n287), .B2(new_n562), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n279), .A2(new_n210), .A3(G87), .ZN(new_n567));
  NOR2_X1   g0367(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n472), .A2(G20), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n210), .B2(G107), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g0374(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n569), .B(new_n574), .C1(new_n567), .C2(new_n575), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n576), .B(KEYINPUT24), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n251), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT25), .B1(new_n262), .B2(new_n206), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n459), .A2(new_n206), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n563), .B(KEYINPUT86), .C1(new_n287), .C2(new_n562), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n566), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n561), .A2(G190), .A3(new_n540), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n562), .A2(G200), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n578), .A2(new_n583), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n279), .A2(new_n280), .A3(G257), .ZN(new_n591));
  INV_X1    g0391(.A(G303), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n279), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n283), .A2(new_n228), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n269), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n515), .A2(G270), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n540), .A3(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n263), .B(G116), .C1(G1), .C2(new_n299), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n262), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n501), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n251), .C1(new_n210), .C2(G116), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n598), .B(new_n600), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n597), .A2(KEYINPUT21), .A3(G169), .A4(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n540), .A2(new_n596), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n608), .A2(new_n606), .A3(G179), .A4(new_n595), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n597), .A2(G169), .A3(new_n606), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n606), .B1(new_n597), .B2(G200), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n380), .B2(new_n597), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n610), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NOR4_X1   g0417(.A1(new_n445), .A2(new_n557), .A3(new_n590), .A4(new_n617), .ZN(G372));
  NOR2_X1   g0418(.A1(new_n432), .A2(KEYINPUT18), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n437), .B1(new_n436), .B2(new_n423), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n333), .A2(new_n330), .A3(new_n334), .ZN(new_n622));
  INV_X1    g0422(.A(new_n359), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n332), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT91), .ZN(new_n625));
  INV_X1    g0425(.A(new_n440), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n421), .B2(KEYINPUT17), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n624), .A2(KEYINPUT91), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n621), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n296), .A2(new_n297), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n289), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n489), .A2(new_n487), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n473), .A2(new_n634), .A3(new_n269), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n473), .B2(new_n269), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n470), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n427), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  INV_X1    g0440(.A(new_n613), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n607), .A2(new_n609), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n610), .A2(KEYINPUT89), .A3(new_n613), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n584), .A2(new_n564), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n460), .B(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n482), .B1(G200), .B2(new_n637), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n649), .A2(new_n650), .B1(new_n633), .B2(new_n638), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n589), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n549), .A2(new_n551), .A3(new_n556), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n639), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n548), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT26), .B1(new_n657), .B2(new_n651), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n494), .B1(new_n549), .B2(new_n551), .ZN(new_n659));
  XNOR2_X1  g0459(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n632), .B1(new_n445), .B2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n606), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n643), .A2(new_n644), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n617), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n670), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n578), .B2(new_n583), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n590), .A2(new_n677), .B1(new_n586), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n676), .B1(new_n641), .B2(new_n642), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n590), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n646), .A2(new_n670), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  INV_X1    g0485(.A(new_n213), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(G41), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n213), .A2(KEYINPUT92), .A3(new_n337), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n451), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n218), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT93), .B1(new_n659), .B2(new_n661), .ZN(new_n694));
  INV_X1    g0494(.A(new_n551), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n539), .A2(KEYINPUT78), .A3(new_n542), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n545), .A2(new_n546), .A3(new_n542), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT78), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n550), .B1(new_n700), .B2(new_n536), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n495), .B1(new_n695), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(new_n703), .A3(new_n660), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n657), .A2(KEYINPUT26), .A3(new_n651), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n694), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n639), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n641), .A2(new_n642), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n652), .B1(new_n586), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n655), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n670), .B1(new_n706), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n663), .B2(new_n670), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n479), .A2(new_n561), .ZN(new_n716));
  AND4_X1   g0516(.A1(G179), .A2(new_n595), .A3(new_n540), .A4(new_n596), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n553), .A4(KEYINPUT30), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n479), .A2(new_n504), .A3(new_n516), .A4(new_n561), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n608), .A2(G179), .A3(new_n595), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n637), .A2(new_n287), .A3(new_n562), .A4(new_n597), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n718), .B(new_n722), .C1(new_n555), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n670), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n616), .A2(new_n586), .A3(new_n589), .A4(new_n676), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n727), .B(new_n728), .C1(new_n557), .C2(new_n729), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n713), .A2(new_n715), .B1(G330), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n693), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(new_n689), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n261), .A2(G20), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G45), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(G1), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n675), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G330), .B2(new_n673), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n250), .B1(G20), .B2(new_n427), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n247), .A2(G45), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT95), .Z(new_n749));
  NOR2_X1   g0549(.A1(new_n686), .A2(new_n279), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n749), .B(new_n750), .C1(G45), .C2(new_n218), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n686), .A2(new_n303), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(G355), .B1(new_n599), .B2(new_n686), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n747), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n739), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n210), .A2(new_n287), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n210), .A2(G179), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(new_n380), .A3(G200), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n759), .A2(new_n220), .B1(new_n761), .B2(new_n206), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n222), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n756), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n756), .A2(G190), .A3(new_n292), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n279), .B1(new_n766), .B2(new_n226), .C1(new_n394), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n757), .A2(new_n380), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n764), .B(new_n768), .C1(G50), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n760), .A2(new_n765), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n380), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n210), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n762), .B(new_n775), .C1(G97), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n767), .ZN(new_n780));
  INV_X1    g0580(.A(new_n771), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n780), .A2(G322), .B1(new_n781), .B2(G329), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n782), .B(new_n303), .C1(new_n783), .C2(new_n766), .ZN(new_n784));
  INV_X1    g0584(.A(new_n763), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n778), .A2(G294), .B1(new_n785), .B2(G303), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n787), .B2(new_n761), .C1(new_n759), .C2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n769), .B(KEYINPUT96), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n784), .B(new_n789), .C1(G326), .C2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n754), .B(new_n755), .C1(new_n793), .C2(new_n745), .ZN(new_n794));
  INV_X1    g0594(.A(new_n744), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n673), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n741), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  INV_X1    g0598(.A(new_n662), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n652), .B1(new_n646), .B2(new_n645), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n707), .B1(new_n800), .B2(new_n710), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n670), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n358), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n803), .A2(new_n347), .A3(new_n676), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n363), .A2(new_n364), .B1(new_n357), .B2(new_n670), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(new_n359), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n802), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n730), .A2(G330), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n739), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n806), .A2(new_n742), .ZN(new_n812));
  INV_X1    g0612(.A(new_n761), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G68), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n279), .C1(new_n815), .C2(new_n771), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n777), .A2(new_n394), .B1(new_n763), .B2(new_n202), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT99), .B(G143), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n767), .A2(new_n819), .B1(new_n766), .B2(new_n772), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(new_n769), .ZN(new_n822));
  INV_X1    g0622(.A(G150), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n821), .A2(new_n822), .B1(new_n759), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n818), .B1(new_n827), .B2(KEYINPUT34), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(KEYINPUT34), .B2(new_n827), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G97), .A2(new_n778), .B1(new_n769), .B2(G303), .ZN(new_n830));
  INV_X1    g0630(.A(new_n766), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n279), .B1(new_n831), .B2(G116), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n780), .A2(G294), .B1(new_n781), .B2(G311), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n761), .A2(new_n222), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n759), .A2(new_n787), .B1(new_n763), .B2(new_n206), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT97), .Z(new_n838));
  OAI21_X1  g0638(.A(new_n745), .B1(new_n829), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n745), .A2(new_n742), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n226), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n812), .A2(new_n739), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n811), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n734), .A2(new_n209), .ZN(new_n844));
  INV_X1    g0644(.A(G330), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n331), .A2(new_n670), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n332), .A2(new_n335), .A3(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n331), .B(new_n670), .C1(new_n622), .C2(new_n321), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n806), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n728), .B1(new_n557), .B2(new_n729), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n725), .A2(KEYINPUT103), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT103), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n724), .A2(new_n852), .A3(new_n670), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n851), .A2(new_n726), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n849), .B(KEYINPUT104), .C1(new_n850), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n851), .A2(new_n726), .A3(new_n853), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n857), .B(new_n728), .C1(new_n557), .C2(new_n729), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT104), .B1(new_n858), .B2(new_n849), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(new_n668), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n423), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n432), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n421), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n418), .A2(new_n399), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n368), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n436), .B2(new_n863), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n415), .A3(new_n420), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n866), .B1(KEYINPUT37), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n433), .A2(new_n438), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n439), .B1(new_n415), .B2(new_n420), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n872), .A2(new_n873), .A3(new_n626), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n868), .A2(new_n863), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT100), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT100), .ZN(new_n877));
  INV_X1    g0677(.A(new_n875), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n441), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n861), .B(new_n871), .C1(new_n876), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n879), .ZN(new_n881));
  INV_X1    g0681(.A(new_n871), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n860), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n887));
  INV_X1    g0687(.A(new_n864), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n441), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n432), .A2(new_n413), .A3(new_n864), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT101), .B1(new_n891), .B2(new_n866), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT37), .B1(new_n436), .B2(new_n423), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(new_n415), .A3(new_n420), .A4(new_n864), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT101), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n889), .A2(new_n892), .A3(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n898), .A2(KEYINPUT102), .A3(new_n861), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT102), .B1(new_n898), .B2(new_n861), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n887), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n858), .A2(new_n849), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(KEYINPUT40), .A3(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n444), .A2(new_n858), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n845), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n321), .A2(new_n331), .A3(new_n676), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n881), .A2(new_n882), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n861), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n909), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n804), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n802), .B2(new_n807), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n847), .A2(new_n848), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n913), .A2(new_n887), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n872), .B2(new_n668), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n713), .A2(new_n715), .A3(new_n444), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n632), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n844), .B1(new_n907), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n926), .B2(new_n907), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n217), .A2(new_n599), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT35), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n527), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n930), .B2(new_n527), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT36), .Z(new_n933));
  NOR3_X1   g0733(.A1(new_n395), .A2(new_n218), .A3(new_n226), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n220), .A2(G50), .ZN(new_n935));
  OAI211_X1 g0735(.A(G1), .B(new_n261), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n928), .A2(new_n933), .A3(new_n936), .ZN(G367));
  INV_X1    g0737(.A(new_n750), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n746), .B1(new_n213), .B2(new_n350), .C1(new_n938), .C2(new_n240), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT108), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n739), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n279), .B1(new_n771), .B2(new_n821), .C1(new_n202), .C2(new_n766), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n759), .A2(new_n772), .B1(new_n763), .B2(new_n394), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n944), .B(new_n945), .C1(G77), .C2(new_n813), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n777), .A2(new_n220), .B1(new_n767), .B2(new_n823), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT111), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n946), .B(new_n948), .C1(new_n790), .C2(new_n819), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n791), .A2(G311), .B1(G303), .B2(new_n780), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n778), .A2(G107), .B1(new_n813), .B2(G97), .ZN(new_n952));
  INV_X1    g0752(.A(G294), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n759), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT46), .B1(new_n785), .B2(G116), .ZN(new_n955));
  INV_X1    g0755(.A(G317), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n303), .B1(new_n771), .B2(new_n956), .C1(new_n787), .C2(new_n766), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n785), .A2(KEYINPUT46), .A3(G116), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT110), .Z(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n950), .A2(KEYINPUT109), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n949), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n941), .B(new_n943), .C1(new_n964), .C2(new_n745), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n649), .A2(new_n676), .ZN(new_n966));
  MUX2_X1   g0766(.A(new_n651), .B(new_n707), .S(new_n966), .Z(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n967), .B2(new_n795), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n710), .B1(new_n552), .B2(new_n676), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n657), .A2(new_n670), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n681), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT42), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n971), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n586), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n549), .A2(new_n551), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n676), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n975), .A2(new_n679), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n980), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n982), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n985), .B1(new_n984), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n689), .B(KEYINPUT41), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT105), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n971), .A2(new_n993), .A3(new_n683), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n971), .B2(new_n683), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT45), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n971), .A2(new_n683), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT44), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n996), .B1(new_n994), .B2(new_n995), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(new_n675), .A3(new_n678), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n681), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n680), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n678), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1003), .B(new_n1006), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n731), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n997), .A2(new_n999), .A3(new_n679), .A4(new_n1000), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1002), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n992), .B1(new_n1011), .B2(new_n731), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n738), .B(KEYINPUT107), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n968), .B1(new_n991), .B2(new_n1014), .ZN(G387));
  NOR2_X1   g0815(.A1(new_n1009), .A2(new_n689), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n731), .B2(new_n1007), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n690), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n752), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(G107), .B2(new_n213), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n237), .A2(new_n463), .ZN(new_n1021));
  AOI211_X1 g0821(.A(G45), .B(new_n1018), .C1(G68), .C2(G77), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n253), .A2(G50), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n938), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1020), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n739), .B1(new_n1026), .B2(new_n747), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n767), .A2(new_n202), .B1(new_n771), .B2(new_n823), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n303), .B(new_n1028), .C1(G68), .C2(new_n831), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n763), .A2(new_n226), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G97), .B2(new_n813), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n486), .A2(new_n777), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G159), .A2(new_n769), .B1(new_n758), .B2(new_n254), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n780), .A2(G317), .B1(new_n831), .B2(G303), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n783), .B2(new_n759), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n791), .B2(G322), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT112), .Z(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(KEYINPUT48), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(KEYINPUT48), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n777), .A2(new_n787), .B1(new_n763), .B2(new_n953), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(KEYINPUT49), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n279), .B1(new_n781), .B2(G326), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n599), .C2(new_n761), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1043), .A2(KEYINPUT49), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1034), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1027), .B1(new_n1048), .B2(new_n745), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n678), .A2(new_n795), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1049), .A2(new_n1050), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1017), .A2(new_n1051), .ZN(G393));
  NAND3_X1  g0852(.A1(new_n1002), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n746), .B1(new_n205), .B2(new_n213), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n750), .B2(new_n244), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n822), .A2(new_n956), .B1(new_n783), .B2(new_n767), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n766), .A2(new_n953), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n279), .B(new_n1058), .C1(G322), .C2(new_n781), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n758), .A2(G303), .B1(new_n813), .B2(G107), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n778), .A2(G116), .B1(new_n785), .B2(G283), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n822), .A2(new_n823), .B1(new_n772), .B2(new_n767), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT51), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n771), .A2(new_n819), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n303), .B(new_n1065), .C1(new_n254), .C2(new_n831), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n759), .A2(new_n202), .B1(new_n763), .B2(new_n220), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n777), .A2(new_n226), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1067), .A2(new_n835), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n755), .B(new_n1055), .C1(new_n1071), .C2(new_n745), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n971), .B2(new_n795), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1053), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1011), .A2(new_n733), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n1008), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  NAND3_X1  g0879(.A1(new_n858), .A2(G330), .A3(new_n849), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n676), .B1(new_n656), .B2(new_n662), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n805), .A2(new_n359), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n804), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n911), .B1(new_n1084), .B2(new_n918), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n909), .B2(new_n914), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n901), .A2(new_n910), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1083), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n916), .B1(new_n712), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n919), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1081), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n910), .B1(new_n917), .B2(new_n919), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT102), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n897), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n864), .B1(new_n627), .B2(new_n621), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n896), .B1(new_n894), .B2(new_n895), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1094), .B1(new_n1098), .B2(KEYINPUT38), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n898), .A2(KEYINPUT102), .A3(new_n861), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT39), .B1(new_n1101), .B2(new_n887), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n883), .A2(new_n880), .A3(new_n908), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1093), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n901), .B(new_n910), .C1(new_n919), .C2(new_n1089), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n730), .A2(G330), .A3(new_n807), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1106), .A2(new_n919), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1104), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n858), .A2(G330), .A3(new_n807), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n919), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n919), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1080), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1111), .A2(new_n1089), .B1(new_n1084), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n444), .A2(G330), .A3(new_n858), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n924), .A2(new_n632), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1092), .A2(new_n1109), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT113), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT113), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1092), .A2(new_n1109), .A3(new_n1120), .A4(new_n1117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1092), .A2(new_n1109), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1117), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n689), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1013), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n742), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n840), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n739), .B1(new_n254), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1068), .B1(G283), .B2(new_n769), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n206), .B2(new_n759), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n767), .A2(new_n599), .B1(new_n771), .B2(new_n953), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n279), .B(new_n1134), .C1(G97), .C2(new_n831), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n764), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n814), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n758), .A2(G137), .B1(new_n831), .B2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT114), .Z(new_n1141));
  NOR2_X1   g0941(.A1(new_n763), .A2(new_n823), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT53), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n279), .B1(new_n767), .B2(new_n815), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G125), .B2(new_n781), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n813), .A2(G50), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G159), .A2(new_n778), .B1(new_n769), .B2(G128), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1133), .A2(new_n1137), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1131), .B1(new_n1149), .B2(new_n745), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1128), .B1(new_n1129), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1126), .A2(new_n1151), .ZN(G378));
  NOR2_X1   g0952(.A1(new_n279), .A2(G41), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n787), .B2(new_n771), .C1(new_n206), .C2(new_n767), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1030), .B(new_n1154), .C1(G68), .C2(new_n778), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n822), .A2(new_n599), .B1(new_n761), .B2(new_n394), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G97), .B2(new_n758), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(new_n486), .C2(new_n766), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT58), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G150), .A2(new_n778), .B1(new_n769), .B2(G125), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT115), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n780), .A2(G128), .B1(new_n831), .B2(G137), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n763), .B2(new_n1138), .C1(new_n815), .C2(new_n759), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT116), .Z(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  OR2_X1    g0967(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(KEYINPUT117), .A2(G124), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n781), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1170), .A2(new_n299), .A3(new_n337), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1167), .B(new_n1171), .C1(new_n772), .C2(new_n761), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1159), .B1(new_n1153), .B2(new_n1160), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT118), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n745), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1174), .A2(KEYINPUT118), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n739), .B1(G50), .B2(new_n1130), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n268), .A2(new_n863), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n298), .B(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT119), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(KEYINPUT119), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1178), .B1(new_n1187), .B2(new_n742), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT120), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n880), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n1191));
  OAI21_X1  g0991(.A(G330), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT40), .B1(new_n921), .B2(new_n860), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT121), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT121), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n886), .A2(new_n903), .A3(new_n1195), .A4(G330), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1187), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n923), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1186), .B(KEYINPUT121), .C1(new_n1193), .C2(new_n1192), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1198), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1189), .B1(new_n1202), .B2(new_n1013), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n924), .A2(new_n632), .A3(new_n1115), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1122), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT57), .B1(new_n1205), .B2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n923), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(KEYINPUT57), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1116), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n733), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1203), .B1(new_n1206), .B2(new_n1212), .ZN(G375));
  INV_X1    g1013(.A(new_n992), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1124), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n739), .B1(G68), .B2(new_n1130), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n777), .A2(new_n202), .B1(new_n763), .B2(new_n772), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G132), .B2(new_n769), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n303), .B1(new_n781), .B2(G128), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n780), .A2(G137), .B1(new_n831), .B2(G150), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n758), .A2(new_n1139), .B1(new_n813), .B2(G58), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1032), .B1(new_n787), .B2(new_n767), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT122), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n759), .A2(new_n599), .B1(new_n761), .B2(new_n226), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n822), .A2(new_n953), .B1(new_n763), .B2(new_n205), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n303), .B1(new_n771), .B2(new_n592), .C1(new_n206), .C2(new_n766), .ZN(new_n1228));
  OR3_X1    g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1223), .B1(new_n1225), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1217), .B1(new_n1230), .B2(new_n745), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n918), .B2(new_n743), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1114), .B2(new_n1127), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1216), .A2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT123), .ZN(G381));
  INV_X1    g1036(.A(new_n1189), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(new_n1127), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT57), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1200), .A2(new_n1201), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n689), .B1(new_n1205), .B2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1211), .B2(new_n1238), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1239), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT124), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n990), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1078), .A3(new_n968), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G381), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .A4(new_n1250), .ZN(G407));
  NAND2_X1  g1051(.A1(new_n669), .A2(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1244), .A2(new_n1245), .A3(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(G407), .A2(G213), .A3(new_n1254), .ZN(G409));
  XNOR2_X1  g1055(.A(G393), .B(new_n797), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1248), .A2(new_n1078), .A3(new_n968), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1078), .B1(new_n1248), .B2(new_n968), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G387), .A2(G390), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1256), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1249), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT126), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1215), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1111), .A2(new_n1089), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1084), .A2(new_n1113), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n689), .B1(new_n1204), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1114), .A2(new_n1116), .A3(KEYINPUT60), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1266), .A2(new_n1270), .A3(KEYINPUT125), .A4(new_n1271), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G384), .B1(new_n1276), .B2(new_n1234), .ZN(new_n1277));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1278), .B(new_n1233), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1264), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n733), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT60), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT125), .B1(new_n1283), .B2(new_n1271), .ZN(new_n1284));
  AND4_X1   g1084(.A1(KEYINPUT125), .A2(new_n1266), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1234), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1278), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1276), .A2(G384), .A3(new_n1234), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(KEYINPUT126), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1253), .A2(G2897), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1280), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G2897), .A3(new_n1253), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1205), .A2(new_n1214), .A3(new_n1202), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G378), .B1(new_n1295), .B2(new_n1203), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1244), .B2(G378), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1297), .B2(new_n1253), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G378), .B(new_n1203), .C1(new_n1206), .C2(new_n1212), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1211), .A2(new_n1238), .A3(new_n992), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1245), .B1(new_n1301), .B2(new_n1239), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  AND2_X1   g1104(.A1(new_n1280), .A2(new_n1289), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1252), .A4(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1298), .A2(new_n1299), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1253), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1304), .B1(new_n1308), .B2(new_n1305), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1263), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1259), .A2(new_n1262), .A3(new_n1299), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1311), .B(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1308), .A2(new_n1305), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1308), .A2(KEYINPUT63), .A3(new_n1305), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1313), .A2(new_n1316), .A3(new_n1298), .A4(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1310), .A2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1245), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1300), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1305), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1292), .A3(new_n1300), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1263), .ZN(G402));
endmodule


