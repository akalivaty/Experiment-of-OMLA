

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U551 ( .A(n667), .B(n666), .ZN(G160) );
  AND2_X2 U552 ( .A1(n652), .A2(G2105), .ZN(n724) );
  NOR2_X1 U553 ( .A1(n825), .A2(G171), .ZN(n827) );
  INV_X1 U554 ( .A(KEYINPUT103), .ZN(n826) );
  NOR2_X1 U555 ( .A1(G2084), .A2(n840), .ZN(n852) );
  INV_X1 U556 ( .A(KEYINPUT17), .ZN(n650) );
  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n651) );
  XOR2_X1 U558 ( .A(n662), .B(n661), .Z(n518) );
  XOR2_X1 U559 ( .A(KEYINPUT74), .B(n541), .Z(n519) );
  XOR2_X1 U560 ( .A(n964), .B(n616), .Z(n520) );
  INV_X1 U561 ( .A(n817), .ZN(n805) );
  XNOR2_X1 U562 ( .A(n819), .B(KEYINPUT99), .ZN(n817) );
  INV_X1 U563 ( .A(G168), .ZN(n831) );
  NOR2_X1 U564 ( .A1(G651), .A2(n533), .ZN(n607) );
  NOR2_X1 U565 ( .A1(G397), .A2(n747), .ZN(n748) );
  XNOR2_X1 U566 ( .A(KEYINPUT69), .B(G651), .ZN(n527) );
  XNOR2_X1 U567 ( .A(KEYINPUT70), .B(n529), .ZN(n604) );
  XNOR2_X1 U568 ( .A(KEYINPUT75), .B(n545), .ZN(n797) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n533) );
  NAND2_X1 U570 ( .A1(G48), .A2(n607), .ZN(n523) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n521) );
  XOR2_X1 U572 ( .A(KEYINPUT65), .B(n521), .Z(n603) );
  NAND2_X1 U573 ( .A1(G86), .A2(n603), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n523), .A2(n522), .ZN(n526) );
  NOR2_X1 U575 ( .A1(n533), .A2(n527), .ZN(n608) );
  NAND2_X1 U576 ( .A1(n608), .A2(G73), .ZN(n524) );
  XOR2_X1 U577 ( .A(KEYINPUT2), .B(n524), .Z(n525) );
  NOR2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n531) );
  NOR2_X1 U579 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n528), .Z(n529) );
  NAND2_X1 U581 ( .A1(G61), .A2(n604), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(G305) );
  NAND2_X1 U583 ( .A1(G74), .A2(G651), .ZN(n532) );
  XNOR2_X1 U584 ( .A(n532), .B(KEYINPUT88), .ZN(n538) );
  NAND2_X1 U585 ( .A1(G49), .A2(n607), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G87), .A2(n533), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U588 ( .A1(n604), .A2(n536), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(G288) );
  NAND2_X1 U590 ( .A1(n608), .A2(G78), .ZN(n544) );
  NAND2_X1 U591 ( .A1(G53), .A2(n607), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G91), .A2(n603), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n604), .A2(G65), .ZN(n541) );
  NOR2_X1 U595 ( .A1(n542), .A2(n519), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n545) );
  INV_X1 U597 ( .A(n797), .ZN(G299) );
  NAND2_X1 U598 ( .A1(G50), .A2(n607), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G88), .A2(n603), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G62), .A2(n604), .ZN(n548) );
  XNOR2_X1 U602 ( .A(KEYINPUT89), .B(n548), .ZN(n549) );
  NOR2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n608), .A2(G75), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(G303) );
  INV_X1 U606 ( .A(G303), .ZN(G166) );
  NAND2_X1 U607 ( .A1(n607), .A2(G47), .ZN(n553) );
  XOR2_X1 U608 ( .A(KEYINPUT71), .B(n553), .Z(n555) );
  NAND2_X1 U609 ( .A1(G60), .A2(n604), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U611 ( .A(KEYINPUT72), .B(n556), .Z(n560) );
  NAND2_X1 U612 ( .A1(G85), .A2(n603), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G72), .A2(n608), .ZN(n557) );
  AND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(G290) );
  NAND2_X1 U616 ( .A1(G51), .A2(n607), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G63), .A2(n604), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U619 ( .A(KEYINPUT6), .B(n563), .ZN(n570) );
  NAND2_X1 U620 ( .A1(n603), .A2(G89), .ZN(n564) );
  XNOR2_X1 U621 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U622 ( .A1(G76), .A2(n608), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U624 ( .A(KEYINPUT5), .B(n567), .Z(n568) );
  XNOR2_X1 U625 ( .A(KEYINPUT80), .B(n568), .ZN(n569) );
  NOR2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U627 ( .A(KEYINPUT7), .B(n571), .Z(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U629 ( .A1(G52), .A2(n607), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G64), .A2(n604), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U632 ( .A(KEYINPUT73), .B(n574), .Z(n579) );
  NAND2_X1 U633 ( .A1(G90), .A2(n603), .ZN(n576) );
  NAND2_X1 U634 ( .A1(G77), .A2(n608), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U637 ( .A1(n579), .A2(n578), .ZN(G171) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G56), .A2(n604), .ZN(n580) );
  XNOR2_X1 U640 ( .A(KEYINPUT14), .B(n580), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n603), .A2(G81), .ZN(n581) );
  XNOR2_X1 U642 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G68), .A2(n608), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U645 ( .A(KEYINPUT13), .B(n584), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U647 ( .A(n587), .B(KEYINPUT77), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n607), .A2(G43), .ZN(n588) );
  NAND2_X1 U649 ( .A1(n589), .A2(n588), .ZN(n964) );
  NAND2_X1 U650 ( .A1(G80), .A2(n608), .ZN(n590) );
  XNOR2_X1 U651 ( .A(n590), .B(KEYINPUT86), .ZN(n597) );
  NAND2_X1 U652 ( .A1(G55), .A2(n607), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G93), .A2(n603), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G67), .A2(n604), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT87), .B(n593), .ZN(n594) );
  NOR2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U658 ( .A1(n597), .A2(n596), .ZN(n779) );
  XNOR2_X1 U659 ( .A(KEYINPUT19), .B(G305), .ZN(n598) );
  XNOR2_X1 U660 ( .A(n598), .B(G288), .ZN(n599) );
  XNOR2_X1 U661 ( .A(n779), .B(n599), .ZN(n601) );
  XOR2_X1 U662 ( .A(G299), .B(G166), .Z(n600) );
  XNOR2_X1 U663 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U664 ( .A(n602), .B(G290), .ZN(n776) );
  XOR2_X1 U665 ( .A(n776), .B(G286), .Z(n615) );
  NAND2_X1 U666 ( .A1(n603), .A2(G92), .ZN(n606) );
  NAND2_X1 U667 ( .A1(G66), .A2(n604), .ZN(n605) );
  NAND2_X1 U668 ( .A1(n606), .A2(n605), .ZN(n612) );
  NAND2_X1 U669 ( .A1(G54), .A2(n607), .ZN(n610) );
  NAND2_X1 U670 ( .A1(G79), .A2(n608), .ZN(n609) );
  NAND2_X1 U671 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U672 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U673 ( .A(KEYINPUT15), .B(n613), .ZN(n756) );
  INV_X1 U674 ( .A(n756), .ZN(n969) );
  XOR2_X1 U675 ( .A(G301), .B(n969), .Z(n614) );
  XNOR2_X1 U676 ( .A(n615), .B(n614), .ZN(n616) );
  NOR2_X1 U677 ( .A1(G37), .A2(n520), .ZN(n617) );
  XOR2_X1 U678 ( .A(KEYINPUT119), .B(n617), .Z(G397) );
  XOR2_X1 U679 ( .A(G2446), .B(G2451), .Z(n619) );
  XNOR2_X1 U680 ( .A(G2454), .B(KEYINPUT111), .ZN(n618) );
  XNOR2_X1 U681 ( .A(n619), .B(n618), .ZN(n626) );
  XOR2_X1 U682 ( .A(G2438), .B(G2430), .Z(n621) );
  XNOR2_X1 U683 ( .A(G2435), .B(G2443), .ZN(n620) );
  XNOR2_X1 U684 ( .A(n621), .B(n620), .ZN(n622) );
  XOR2_X1 U685 ( .A(n622), .B(G2427), .Z(n624) );
  XNOR2_X1 U686 ( .A(G1341), .B(G1348), .ZN(n623) );
  XNOR2_X1 U687 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U688 ( .A(n626), .B(n625), .ZN(n627) );
  AND2_X1 U689 ( .A1(n627), .A2(G14), .ZN(G401) );
  XNOR2_X1 U690 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U691 ( .A(G82), .ZN(G220) );
  INV_X1 U692 ( .A(G132), .ZN(G219) );
  INV_X1 U693 ( .A(G57), .ZN(G237) );
  XOR2_X1 U694 ( .A(KEYINPUT113), .B(G2678), .Z(n629) );
  XNOR2_X1 U695 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n629), .B(n628), .ZN(n633) );
  XOR2_X1 U697 ( .A(KEYINPUT114), .B(G2090), .Z(n631) );
  XNOR2_X1 U698 ( .A(G2067), .B(G2072), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n631), .B(n630), .ZN(n632) );
  XOR2_X1 U700 ( .A(n633), .B(n632), .Z(n635) );
  INV_X1 U701 ( .A(G2100), .ZN(n770) );
  XOR2_X1 U702 ( .A(G2096), .B(n770), .Z(n634) );
  XNOR2_X1 U703 ( .A(n635), .B(n634), .ZN(n637) );
  XOR2_X1 U704 ( .A(G2078), .B(G2084), .Z(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(G227) );
  XOR2_X1 U706 ( .A(G1976), .B(G1971), .Z(n639) );
  INV_X1 U707 ( .A(G1956), .ZN(n959) );
  XOR2_X1 U708 ( .A(G1986), .B(n959), .Z(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U710 ( .A(n640), .B(G2474), .Z(n642) );
  XNOR2_X1 U711 ( .A(G1966), .B(G1981), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(n646) );
  XOR2_X1 U713 ( .A(KEYINPUT41), .B(G1961), .Z(n644) );
  XNOR2_X1 U714 ( .A(G1996), .B(G1991), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(G229) );
  INV_X1 U717 ( .A(G2104), .ZN(n652) );
  NAND2_X1 U718 ( .A1(G126), .A2(n724), .ZN(n648) );
  AND2_X1 U719 ( .A1(G2104), .A2(G2105), .ZN(n725) );
  NAND2_X1 U720 ( .A1(G114), .A2(n725), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U722 ( .A(KEYINPUT94), .B(n649), .ZN(n656) );
  XNOR2_X2 U723 ( .A(n651), .B(n650), .ZN(n733) );
  NAND2_X1 U724 ( .A1(G138), .A2(n733), .ZN(n654) );
  NOR2_X1 U725 ( .A1(G2105), .A2(n652), .ZN(n660) );
  BUF_X1 U726 ( .A(n660), .Z(n728) );
  NAND2_X1 U727 ( .A1(G102), .A2(n728), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n656), .A2(n655), .ZN(G164) );
  NAND2_X1 U730 ( .A1(G113), .A2(n725), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n733), .A2(G137), .ZN(n657) );
  AND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n665) );
  NAND2_X1 U733 ( .A1(G125), .A2(n724), .ZN(n659) );
  XNOR2_X1 U734 ( .A(KEYINPUT67), .B(n659), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT23), .B(KEYINPUT68), .Z(n662) );
  NAND2_X1 U736 ( .A1(G101), .A2(n660), .ZN(n661) );
  NOR2_X1 U737 ( .A1(n663), .A2(n518), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n667) );
  INV_X1 U739 ( .A(KEYINPUT66), .ZN(n666) );
  NAND2_X1 U740 ( .A1(G112), .A2(n725), .ZN(n669) );
  NAND2_X1 U741 ( .A1(G100), .A2(n728), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n675) );
  NAND2_X1 U743 ( .A1(n724), .A2(G124), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n670), .B(KEYINPUT44), .ZN(n672) );
  NAND2_X1 U745 ( .A1(G136), .A2(n733), .ZN(n671) );
  NAND2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U747 ( .A(KEYINPUT115), .B(n673), .Z(n674) );
  NOR2_X1 U748 ( .A1(n675), .A2(n674), .ZN(G162) );
  NAND2_X1 U749 ( .A1(G119), .A2(n724), .ZN(n677) );
  NAND2_X1 U750 ( .A1(G131), .A2(n733), .ZN(n676) );
  NAND2_X1 U751 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U752 ( .A1(G107), .A2(n725), .ZN(n679) );
  NAND2_X1 U753 ( .A1(G95), .A2(n728), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n679), .A2(n678), .ZN(n680) );
  OR2_X1 U755 ( .A1(n681), .A2(n680), .ZN(n903) );
  XOR2_X1 U756 ( .A(KEYINPUT116), .B(KEYINPUT48), .Z(n683) );
  XNOR2_X1 U757 ( .A(KEYINPUT46), .B(KEYINPUT118), .ZN(n682) );
  XNOR2_X1 U758 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U759 ( .A(n903), .B(n684), .ZN(n695) );
  NAND2_X1 U760 ( .A1(G128), .A2(n724), .ZN(n686) );
  NAND2_X1 U761 ( .A1(G116), .A2(n725), .ZN(n685) );
  NAND2_X1 U762 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U763 ( .A(n687), .B(KEYINPUT35), .ZN(n692) );
  NAND2_X1 U764 ( .A1(G140), .A2(n733), .ZN(n689) );
  NAND2_X1 U765 ( .A1(G104), .A2(n728), .ZN(n688) );
  NAND2_X1 U766 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U767 ( .A(KEYINPUT34), .B(n690), .Z(n691) );
  NAND2_X1 U768 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U769 ( .A(n693), .B(KEYINPUT36), .Z(n913) );
  XOR2_X1 U770 ( .A(G164), .B(n913), .Z(n694) );
  XNOR2_X1 U771 ( .A(n695), .B(n694), .ZN(n723) );
  NAND2_X1 U772 ( .A1(n724), .A2(G123), .ZN(n696) );
  XNOR2_X1 U773 ( .A(n696), .B(KEYINPUT18), .ZN(n698) );
  NAND2_X1 U774 ( .A1(G135), .A2(n733), .ZN(n697) );
  NAND2_X1 U775 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U776 ( .A(KEYINPUT84), .B(n699), .ZN(n703) );
  NAND2_X1 U777 ( .A1(G111), .A2(n725), .ZN(n701) );
  NAND2_X1 U778 ( .A1(G99), .A2(n728), .ZN(n700) );
  NAND2_X1 U779 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U780 ( .A1(n703), .A2(n702), .ZN(n937) );
  NAND2_X1 U781 ( .A1(G130), .A2(n724), .ZN(n705) );
  NAND2_X1 U782 ( .A1(G118), .A2(n725), .ZN(n704) );
  NAND2_X1 U783 ( .A1(n705), .A2(n704), .ZN(n710) );
  NAND2_X1 U784 ( .A1(G142), .A2(n733), .ZN(n707) );
  NAND2_X1 U785 ( .A1(G106), .A2(n728), .ZN(n706) );
  NAND2_X1 U786 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U787 ( .A(KEYINPUT45), .B(n708), .Z(n709) );
  NOR2_X1 U788 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U789 ( .A(n937), .B(n711), .ZN(n721) );
  NAND2_X1 U790 ( .A1(G139), .A2(n733), .ZN(n713) );
  NAND2_X1 U791 ( .A1(G103), .A2(n728), .ZN(n712) );
  NAND2_X1 U792 ( .A1(n713), .A2(n712), .ZN(n718) );
  NAND2_X1 U793 ( .A1(G127), .A2(n724), .ZN(n715) );
  NAND2_X1 U794 ( .A1(G115), .A2(n725), .ZN(n714) );
  NAND2_X1 U795 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U796 ( .A(KEYINPUT47), .B(n716), .Z(n717) );
  NOR2_X1 U797 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U798 ( .A(KEYINPUT117), .B(n719), .Z(n931) );
  XNOR2_X1 U799 ( .A(G160), .B(n931), .ZN(n720) );
  XNOR2_X1 U800 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U801 ( .A(n723), .B(n722), .ZN(n737) );
  NAND2_X1 U802 ( .A1(G129), .A2(n724), .ZN(n727) );
  NAND2_X1 U803 ( .A1(G117), .A2(n725), .ZN(n726) );
  NAND2_X1 U804 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n728), .A2(G105), .ZN(n729) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(n729), .Z(n730) );
  NOR2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U808 ( .A(n732), .B(KEYINPUT96), .ZN(n735) );
  NAND2_X1 U809 ( .A1(G141), .A2(n733), .ZN(n734) );
  NAND2_X1 U810 ( .A1(n735), .A2(n734), .ZN(n902) );
  XNOR2_X1 U811 ( .A(n902), .B(G162), .ZN(n736) );
  XNOR2_X1 U812 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U813 ( .A1(G37), .A2(n738), .ZN(G395) );
  NOR2_X1 U814 ( .A1(G220), .A2(G219), .ZN(n739) );
  XOR2_X1 U815 ( .A(KEYINPUT22), .B(n739), .Z(n740) );
  NOR2_X1 U816 ( .A1(G218), .A2(n740), .ZN(n741) );
  NAND2_X1 U817 ( .A1(G96), .A2(n741), .ZN(n925) );
  NAND2_X1 U818 ( .A1(n925), .A2(G2106), .ZN(n745) );
  NAND2_X1 U819 ( .A1(G69), .A2(G120), .ZN(n742) );
  NOR2_X1 U820 ( .A1(G237), .A2(n742), .ZN(n743) );
  NAND2_X1 U821 ( .A1(G108), .A2(n743), .ZN(n924) );
  NAND2_X1 U822 ( .A1(n924), .A2(G567), .ZN(n744) );
  NAND2_X1 U823 ( .A1(n745), .A2(n744), .ZN(n927) );
  NOR2_X1 U824 ( .A1(G401), .A2(n927), .ZN(n749) );
  NOR2_X1 U825 ( .A1(G227), .A2(G229), .ZN(n746) );
  XNOR2_X1 U826 ( .A(KEYINPUT49), .B(n746), .ZN(n747) );
  NAND2_X1 U827 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U828 ( .A1(n750), .A2(G395), .ZN(n751) );
  XNOR2_X1 U829 ( .A(n751), .B(KEYINPUT120), .ZN(G308) );
  INV_X1 U830 ( .A(G308), .ZN(G225) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U832 ( .A1(G7), .A2(G661), .ZN(n752) );
  XNOR2_X1 U833 ( .A(n752), .B(KEYINPUT10), .ZN(n753) );
  XOR2_X1 U834 ( .A(KEYINPUT76), .B(n753), .Z(n920) );
  NAND2_X1 U835 ( .A1(n920), .A2(G567), .ZN(n754) );
  XOR2_X1 U836 ( .A(KEYINPUT11), .B(n754), .Z(G234) );
  XOR2_X1 U837 ( .A(G860), .B(KEYINPUT78), .Z(n764) );
  NOR2_X1 U838 ( .A1(n964), .A2(n764), .ZN(n755) );
  XNOR2_X1 U839 ( .A(n755), .B(KEYINPUT79), .ZN(G153) );
  NAND2_X1 U840 ( .A1(G868), .A2(G301), .ZN(n758) );
  INV_X1 U841 ( .A(G868), .ZN(n780) );
  NAND2_X1 U842 ( .A1(n756), .A2(n780), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n758), .A2(n757), .ZN(G284) );
  NOR2_X1 U844 ( .A1(G868), .A2(G299), .ZN(n759) );
  XOR2_X1 U845 ( .A(KEYINPUT82), .B(n759), .Z(n762) );
  NOR2_X1 U846 ( .A1(G286), .A2(n780), .ZN(n760) );
  XNOR2_X1 U847 ( .A(KEYINPUT81), .B(n760), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U849 ( .A(KEYINPUT83), .B(n763), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n764), .A2(G559), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n765), .A2(n969), .ZN(n766) );
  XNOR2_X1 U852 ( .A(n766), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U853 ( .A1(G868), .A2(n964), .ZN(n769) );
  NAND2_X1 U854 ( .A1(G868), .A2(n969), .ZN(n767) );
  NOR2_X1 U855 ( .A1(G559), .A2(n767), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n769), .A2(n768), .ZN(G282) );
  XNOR2_X1 U857 ( .A(n937), .B(G2096), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(G156) );
  XNOR2_X1 U859 ( .A(n964), .B(KEYINPUT85), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G559), .A2(n969), .ZN(n772) );
  XOR2_X1 U861 ( .A(n773), .B(n772), .Z(n775) );
  NOR2_X1 U862 ( .A1(G860), .A2(n775), .ZN(n774) );
  XOR2_X1 U863 ( .A(n779), .B(n774), .Z(G145) );
  XOR2_X1 U864 ( .A(n776), .B(n775), .Z(n777) );
  NAND2_X1 U865 ( .A1(n777), .A2(G868), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT90), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(G295) );
  NAND2_X1 U869 ( .A1(G2078), .A2(G2084), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT20), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(KEYINPUT91), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n785), .A2(G2090), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT21), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(KEYINPUT92), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n788), .A2(G2072), .ZN(G158) );
  NAND2_X1 U876 ( .A1(G661), .A2(G483), .ZN(n789) );
  XOR2_X1 U877 ( .A(KEYINPUT93), .B(n789), .Z(n790) );
  NOR2_X1 U878 ( .A1(n927), .A2(n790), .ZN(n923) );
  NAND2_X1 U879 ( .A1(n923), .A2(G36), .ZN(G176) );
  NOR2_X1 U880 ( .A1(G164), .A2(G1384), .ZN(n863) );
  INV_X1 U881 ( .A(n863), .ZN(n791) );
  NAND2_X1 U882 ( .A1(G40), .A2(G160), .ZN(n862) );
  NOR2_X2 U883 ( .A1(n791), .A2(n862), .ZN(n819) );
  NAND2_X1 U884 ( .A1(n805), .A2(G2072), .ZN(n792) );
  XNOR2_X1 U885 ( .A(n792), .B(KEYINPUT27), .ZN(n794) );
  NOR2_X1 U886 ( .A1(n959), .A2(n805), .ZN(n793) );
  NOR2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n796) );
  NOR2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n795) );
  XOR2_X1 U889 ( .A(n795), .B(KEYINPUT28), .Z(n815) );
  NAND2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n813) );
  INV_X1 U891 ( .A(n819), .ZN(n840) );
  NAND2_X1 U892 ( .A1(G1341), .A2(n840), .ZN(n798) );
  XNOR2_X1 U893 ( .A(n798), .B(KEYINPUT102), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n819), .A2(G1996), .ZN(n799) );
  XNOR2_X1 U895 ( .A(n799), .B(KEYINPUT26), .ZN(n800) );
  XNOR2_X1 U896 ( .A(KEYINPUT64), .B(n800), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U898 ( .A1(n964), .A2(n803), .ZN(n804) );
  OR2_X1 U899 ( .A1(n969), .A2(n804), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n969), .A2(n804), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G2067), .A2(n805), .ZN(n807) );
  NAND2_X1 U902 ( .A1(G1348), .A2(n840), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U908 ( .A(n816), .B(KEYINPUT29), .ZN(n824) );
  XOR2_X1 U909 ( .A(KEYINPUT25), .B(G2078), .Z(n1012) );
  NOR2_X1 U910 ( .A1(n817), .A2(n1012), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(KEYINPUT100), .ZN(n821) );
  NOR2_X1 U912 ( .A1(n819), .A2(G1961), .ZN(n820) );
  NOR2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U914 ( .A(n822), .B(KEYINPUT101), .ZN(n825) );
  AND2_X1 U915 ( .A1(G171), .A2(n825), .ZN(n823) );
  NOR2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n837) );
  XNOR2_X1 U917 ( .A(n827), .B(n826), .ZN(n834) );
  NAND2_X1 U918 ( .A1(G8), .A2(n840), .ZN(n879) );
  NOR2_X1 U919 ( .A1(G1966), .A2(n879), .ZN(n851) );
  XOR2_X1 U920 ( .A(KEYINPUT98), .B(n852), .Z(n828) );
  NAND2_X1 U921 ( .A1(G8), .A2(n828), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n851), .A2(n829), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n830), .B(KEYINPUT30), .ZN(n832) );
  AND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U925 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U926 ( .A(n835), .B(KEYINPUT31), .ZN(n836) );
  NOR2_X1 U927 ( .A1(n837), .A2(n836), .ZN(n839) );
  INV_X1 U928 ( .A(KEYINPUT104), .ZN(n838) );
  XNOR2_X1 U929 ( .A(n839), .B(n838), .ZN(n849) );
  NAND2_X1 U930 ( .A1(n849), .A2(G286), .ZN(n845) );
  NOR2_X1 U931 ( .A1(G1971), .A2(n879), .ZN(n842) );
  NOR2_X1 U932 ( .A1(G2090), .A2(n840), .ZN(n841) );
  NOR2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U934 ( .A1(n843), .A2(G303), .ZN(n844) );
  NAND2_X1 U935 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U936 ( .A(n846), .B(KEYINPUT106), .ZN(n847) );
  NAND2_X1 U937 ( .A1(n847), .A2(G8), .ZN(n848) );
  XNOR2_X1 U938 ( .A(n848), .B(KEYINPUT32), .ZN(n885) );
  XNOR2_X1 U939 ( .A(n849), .B(KEYINPUT105), .ZN(n850) );
  NOR2_X1 U940 ( .A1(n851), .A2(n850), .ZN(n855) );
  XNOR2_X1 U941 ( .A(n852), .B(KEYINPUT98), .ZN(n853) );
  NAND2_X1 U942 ( .A1(G8), .A2(n853), .ZN(n854) );
  NAND2_X1 U943 ( .A1(n855), .A2(n854), .ZN(n883) );
  INV_X1 U944 ( .A(n879), .ZN(n856) );
  NAND2_X1 U945 ( .A1(G1976), .A2(G288), .ZN(n962) );
  AND2_X1 U946 ( .A1(n856), .A2(n962), .ZN(n857) );
  NOR2_X1 U947 ( .A1(KEYINPUT33), .A2(n857), .ZN(n860) );
  NOR2_X1 U948 ( .A1(G1976), .A2(G288), .ZN(n871) );
  NAND2_X1 U949 ( .A1(n871), .A2(KEYINPUT33), .ZN(n858) );
  NOR2_X1 U950 ( .A1(n879), .A2(n858), .ZN(n859) );
  NOR2_X1 U951 ( .A1(n860), .A2(n859), .ZN(n867) );
  XNOR2_X1 U952 ( .A(G1981), .B(KEYINPUT107), .ZN(n861) );
  XNOR2_X1 U953 ( .A(n861), .B(G305), .ZN(n954) );
  NOR2_X1 U954 ( .A1(n863), .A2(n862), .ZN(n916) );
  XNOR2_X1 U955 ( .A(G2067), .B(KEYINPUT37), .ZN(n912) );
  OR2_X1 U956 ( .A1(n912), .A2(n913), .ZN(n864) );
  XNOR2_X1 U957 ( .A(n864), .B(KEYINPUT95), .ZN(n949) );
  NAND2_X1 U958 ( .A1(n916), .A2(n949), .ZN(n910) );
  XNOR2_X1 U959 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U960 ( .A1(n916), .A2(n971), .ZN(n865) );
  AND2_X1 U961 ( .A1(n910), .A2(n865), .ZN(n880) );
  AND2_X1 U962 ( .A1(n954), .A2(n880), .ZN(n866) );
  AND2_X1 U963 ( .A1(n867), .A2(n866), .ZN(n869) );
  AND2_X1 U964 ( .A1(n883), .A2(n869), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n885), .A2(n868), .ZN(n876) );
  INV_X1 U966 ( .A(n869), .ZN(n874) );
  NOR2_X1 U967 ( .A1(G1971), .A2(G303), .ZN(n870) );
  NOR2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n972) );
  INV_X1 U969 ( .A(KEYINPUT33), .ZN(n872) );
  AND2_X1 U970 ( .A1(n972), .A2(n872), .ZN(n873) );
  OR2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n875) );
  AND2_X1 U972 ( .A1(n876), .A2(n875), .ZN(n895) );
  NOR2_X1 U973 ( .A1(G1981), .A2(G305), .ZN(n877) );
  XOR2_X1 U974 ( .A(n877), .B(KEYINPUT24), .Z(n878) );
  NOR2_X1 U975 ( .A1(n879), .A2(n878), .ZN(n887) );
  OR2_X1 U976 ( .A1(n887), .A2(n879), .ZN(n881) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n891) );
  INV_X1 U978 ( .A(n891), .ZN(n882) );
  AND2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  NAND2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n893) );
  NOR2_X1 U981 ( .A1(G2090), .A2(G303), .ZN(n886) );
  NAND2_X1 U982 ( .A1(G8), .A2(n886), .ZN(n889) );
  INV_X1 U983 ( .A(n887), .ZN(n888) );
  AND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  OR2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n892) );
  AND2_X1 U986 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U987 ( .A1(n895), .A2(n894), .ZN(n900) );
  NAND2_X1 U988 ( .A1(G1991), .A2(n903), .ZN(n897) );
  NAND2_X1 U989 ( .A1(G1996), .A2(n902), .ZN(n896) );
  NAND2_X1 U990 ( .A1(n897), .A2(n896), .ZN(n941) );
  NAND2_X1 U991 ( .A1(n941), .A2(n916), .ZN(n898) );
  XOR2_X1 U992 ( .A(KEYINPUT97), .B(n898), .Z(n899) );
  NAND2_X1 U993 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n901), .B(KEYINPUT108), .ZN(n918) );
  NOR2_X1 U995 ( .A1(G1996), .A2(n902), .ZN(n929) );
  NOR2_X1 U996 ( .A1(G1991), .A2(n903), .ZN(n904) );
  XNOR2_X1 U997 ( .A(KEYINPUT110), .B(n904), .ZN(n936) );
  NOR2_X1 U998 ( .A1(G1986), .A2(G290), .ZN(n905) );
  XOR2_X1 U999 ( .A(n905), .B(KEYINPUT109), .Z(n906) );
  NOR2_X1 U1000 ( .A1(n936), .A2(n906), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(n907), .A2(n941), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(n929), .A2(n908), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(n909), .B(KEYINPUT39), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n914) );
  NAND2_X1 U1005 ( .A1(n913), .A2(n912), .ZN(n942) );
  NAND2_X1 U1006 ( .A1(n914), .A2(n942), .ZN(n915) );
  NAND2_X1 U1007 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1008 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1009 ( .A(n919), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U1010 ( .A1(G2106), .A2(n920), .ZN(G217) );
  INV_X1 U1011 ( .A(n920), .ZN(G223) );
  AND2_X1 U1012 ( .A1(G15), .A2(G2), .ZN(n921) );
  NAND2_X1 U1013 ( .A1(G661), .A2(n921), .ZN(G259) );
  NAND2_X1 U1014 ( .A1(G3), .A2(G1), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(G188) );
  INV_X1 U1017 ( .A(G120), .ZN(G236) );
  INV_X1 U1018 ( .A(G96), .ZN(G221) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1021 ( .A(n926), .B(KEYINPUT112), .Z(G261) );
  INV_X1 U1022 ( .A(G261), .ZN(G325) );
  INV_X1 U1023 ( .A(n927), .ZN(G319) );
  INV_X1 U1024 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n930), .Z(n947) );
  XNOR2_X1 U1028 ( .A(G164), .B(G2078), .ZN(n934) );
  XOR2_X1 U1029 ( .A(G2072), .B(n931), .Z(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT121), .B(n932), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT50), .ZN(n945) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G160), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n950), .ZN(n952) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n951) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1044 ( .A1(n953), .A2(G29), .ZN(n1032) );
  XOR2_X1 U1045 ( .A(KEYINPUT56), .B(G16), .Z(n977) );
  XNOR2_X1 U1046 ( .A(G1966), .B(G168), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n956), .B(KEYINPUT57), .ZN(n968) );
  XOR2_X1 U1049 ( .A(G301), .B(G1961), .Z(n958) );
  NAND2_X1 U1050 ( .A1(G1971), .A2(G303), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1052 ( .A(n959), .B(G299), .Z(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n963) );
  NAND2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G1341), .B(n964), .ZN(n965) );
  NOR2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n975) );
  XOR2_X1 U1058 ( .A(G1348), .B(n969), .Z(n970) );
  NOR2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1060 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1061 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1062 ( .A1(n977), .A2(n976), .ZN(n1030) );
  XOR2_X1 U1063 ( .A(G20), .B(G1956), .Z(n981) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n979) );
  XNOR2_X1 U1065 ( .A(G1981), .B(G6), .ZN(n978) );
  NOR2_X1 U1066 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1067 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1068 ( .A(KEYINPUT59), .B(G1348), .Z(n982) );
  XNOR2_X1 U1069 ( .A(G4), .B(n982), .ZN(n983) );
  NOR2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n986) );
  XOR2_X1 U1071 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n985) );
  XNOR2_X1 U1072 ( .A(n986), .B(n985), .ZN(n990) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G21), .ZN(n988) );
  XNOR2_X1 U1074 ( .A(G5), .B(G1961), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n997) );
  XNOR2_X1 U1077 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(G23), .B(G1976), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n994) );
  XOR2_X1 U1080 ( .A(G1986), .B(G24), .Z(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n995), .ZN(n996) );
  NOR2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1084 ( .A(KEYINPUT61), .B(n998), .Z(n1000) );
  XNOR2_X1 U1085 ( .A(G16), .B(KEYINPUT126), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1023) );
  XOR2_X1 U1087 ( .A(G34), .B(KEYINPUT125), .Z(n1002) );
  XNOR2_X1 U1088 ( .A(G2084), .B(KEYINPUT54), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(n1002), .B(n1001), .ZN(n1020) );
  XNOR2_X1 U1090 ( .A(G2090), .B(G35), .ZN(n1017) );
  XNOR2_X1 U1091 ( .A(G2067), .B(G26), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G33), .B(G2072), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(G1991), .B(G25), .Z(n1005) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(G28), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(KEYINPUT122), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G1996), .B(G32), .Z(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT123), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G27), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT124), .B(n1018), .Z(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(KEYINPUT55), .A2(n1024), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(G11), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1028) );
  INV_X1 U1110 ( .A(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1033), .ZN(G150) );
  INV_X1 U1117 ( .A(G150), .ZN(G311) );
endmodule

