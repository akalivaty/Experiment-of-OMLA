//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n202));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(G204gat), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(new_n205), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT75), .B(G218gat), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT22), .B1(new_n213), .B2(G211gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n204), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n217));
  OAI21_X1  g016(.A(G211gat), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT22), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n220), .A2(new_n208), .A3(new_n211), .A4(new_n203), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT3), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G141gat), .B(G148gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n226), .B(new_n229), .C1(new_n230), .C2(KEYINPUT2), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G141gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n229), .A2(new_n226), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n226), .A2(KEYINPUT2), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n231), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n225), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G228gat), .A2(G233gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n231), .A2(new_n239), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n224), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n242), .B1(new_n245), .B2(new_n222), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT29), .B1(new_n215), .B2(new_n221), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n243), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n249));
  INV_X1    g048(.A(new_n222), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n244), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n242), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n202), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n251), .B(new_n242), .C1(new_n225), .C2(new_n240), .ZN(new_n254));
  INV_X1    g053(.A(new_n202), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n249), .A2(new_n251), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n242), .ZN(new_n257));
  XOR2_X1   g056(.A(G78gat), .B(G106gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G50gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G22gat), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n253), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n253), .B2(new_n257), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT79), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n261), .B2(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT67), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n271), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g080(.A1(G183gat), .A2(G190gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G183gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT27), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n290));
  NOR2_X1   g089(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n289), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n284), .A2(new_n288), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT24), .A3(new_n282), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(G183gat), .A3(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n277), .A2(KEYINPUT23), .ZN(new_n300));
  AND4_X1   g099(.A1(new_n297), .A2(new_n299), .A3(new_n270), .A4(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT65), .B1(new_n277), .B2(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(new_n304), .C1(G169gat), .C2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT25), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n300), .A2(new_n299), .A3(new_n270), .ZN(new_n308));
  AND4_X1   g107(.A1(KEYINPUT25), .A2(new_n308), .A3(new_n306), .A4(new_n297), .ZN(new_n309));
  OAI22_X1  g108(.A1(new_n294), .A2(new_n295), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n269), .B1(new_n310), .B2(new_n224), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n280), .A2(new_n282), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT68), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(new_n283), .A3(new_n293), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n306), .A3(new_n297), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n306), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n268), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n250), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n322), .B(new_n323), .Z(new_n324));
  NAND2_X1  g123(.A1(new_n310), .A2(new_n269), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n314), .B2(new_n319), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(new_n222), .C1(new_n326), .C2(new_n269), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT30), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n321), .A2(KEYINPUT77), .A3(new_n327), .A4(new_n324), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT69), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(KEYINPUT1), .ZN(new_n341));
  INV_X1    g140(.A(G134gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n340), .B2(KEYINPUT1), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n341), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(G113gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n352), .B(new_n339), .C1(new_n345), .C2(new_n343), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n240), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI211_X1 g157(.A(KEYINPUT4), .B(new_n243), .C1(new_n353), .C2(new_n347), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n347), .A2(new_n353), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(new_n240), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n334), .B(new_n358), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT5), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n240), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n347), .A2(new_n243), .A3(new_n353), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n334), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n243), .B1(new_n347), .B2(new_n353), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n360), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(new_n364), .A3(new_n334), .A4(new_n358), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT0), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n376), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n370), .A2(new_n375), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n370), .B2(new_n375), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n381), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n324), .B1(new_n321), .B2(new_n327), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n321), .A2(new_n324), .A3(new_n327), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(KEYINPUT30), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n333), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n310), .A2(new_n361), .ZN(new_n392));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT64), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n314), .A2(new_n319), .A3(new_n354), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT32), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G71gat), .B(G99gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT72), .ZN(new_n401));
  XNOR2_X1  g200(.A(G15gat), .B(G43gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(KEYINPUT71), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n401), .B(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n397), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n396), .B(KEYINPUT32), .C1(new_n398), .C2(new_n404), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n395), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n354), .B1(new_n314), .B2(new_n319), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n393), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT34), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n394), .A2(KEYINPUT34), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n409), .B2(new_n410), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT73), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n416), .B(new_n413), .C1(new_n409), .C2(new_n410), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(KEYINPUT34), .A2(new_n411), .B1(new_n414), .B2(KEYINPUT73), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n406), .A3(new_n407), .A4(new_n417), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT36), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(KEYINPUT36), .A3(new_n421), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n267), .A2(new_n391), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n261), .A2(new_n262), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n324), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n321), .A2(new_n327), .ZN(new_n429));
  INV_X1    g228(.A(new_n324), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n321), .B2(new_n327), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT38), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT38), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n222), .B1(new_n311), .B2(new_n320), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n325), .B(new_n250), .C1(new_n326), .C2(new_n269), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(KEYINPUT37), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n436), .B(new_n439), .C1(new_n388), .C2(new_n428), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT82), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT82), .B1(new_n370), .B2(new_n375), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n380), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n385), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n443), .A2(new_n444), .B1(KEYINPUT6), .B2(new_n386), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n330), .A2(new_n332), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n435), .A2(new_n440), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n432), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n388), .B2(new_n428), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(KEYINPUT84), .A3(KEYINPUT38), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n426), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n334), .B1(new_n374), .B2(new_n358), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT80), .B(KEYINPUT39), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n380), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT39), .B1(new_n367), .B2(new_n368), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n358), .B1(new_n359), .B2(new_n362), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n368), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT81), .B(KEYINPUT39), .C1(new_n367), .C2(new_n368), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n455), .A2(KEYINPUT40), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT40), .B1(new_n455), .B2(new_n462), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n443), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n333), .A2(new_n390), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT83), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n376), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT82), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n382), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n472), .A2(new_n463), .A3(new_n464), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n333), .A2(new_n390), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n425), .B1(new_n452), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n426), .A2(new_n421), .A3(new_n419), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT35), .B1(new_n480), .B2(new_n391), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(KEYINPUT85), .B(KEYINPUT35), .C1(new_n480), .C2(new_n391), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n480), .A2(new_n475), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n478), .A2(new_n479), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n479), .B1(new_n478), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n492), .A2(G1gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT16), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n494), .B2(G1gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n492), .A2(G1gat), .ZN(new_n497));
  OAI21_X1  g296(.A(G8gat), .B1(new_n497), .B2(KEYINPUT90), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n496), .B(new_n498), .Z(new_n499));
  XOR2_X1   g298(.A(KEYINPUT87), .B(G29gat), .Z(new_n500));
  INV_X1    g299(.A(G36gat), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT15), .ZN(new_n505));
  NOR2_X1   g304(.A1(G29gat), .A2(G36gat), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n506), .A2(KEYINPUT14), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(KEYINPUT14), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT15), .B1(new_n503), .B2(new_n504), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n502), .A2(new_n505), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(new_n508), .C1(new_n500), .C2(new_n501), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT91), .B1(new_n499), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n496), .B(new_n498), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n512), .A2(new_n514), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(new_n515), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n520), .A2(new_n523), .A3(new_n524), .A4(new_n511), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n499), .A2(new_n518), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT13), .Z(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n518), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n523), .A2(KEYINPUT17), .A3(new_n511), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n520), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n528), .A4(new_n526), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n530), .A2(KEYINPUT92), .A3(new_n535), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n528), .A3(new_n526), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  INV_X1    g343(.A(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT11), .B(G169gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n540), .A2(new_n541), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT93), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n549), .A3(new_n535), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT93), .B1(new_n540), .B2(new_n541), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n491), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G64gat), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n562), .A2(G57gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(G57gat), .ZN(new_n564));
  AND2_X1   g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n563), .A2(new_n564), .B1(new_n565), .B2(KEYINPUT9), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n568));
  NOR2_X1   g367(.A1(G71gat), .A2(G78gat), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n567), .A2(new_n568), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n566), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G127gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n520), .B1(new_n572), .B2(new_n571), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT96), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n578), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT95), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G155gat), .ZN(new_n583));
  XOR2_X1   g382(.A(G183gat), .B(G211gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT97), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n579), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n579), .B2(new_n580), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  XNOR2_X1  g391(.A(G99gat), .B(G106gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g396(.A1(new_n592), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n593), .B1(new_n592), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n590), .B1(new_n518), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n532), .A2(new_n533), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(KEYINPUT98), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT99), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n606), .B(new_n601), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(KEYINPUT99), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G134gat), .B(G162gat), .Z(new_n612));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT100), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n609), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n609), .A2(new_n611), .B1(KEYINPUT100), .B2(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n571), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n600), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n571), .B1(new_n598), .B2(new_n599), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n620), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n623), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(new_n620), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT101), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n625), .A2(new_n626), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n619), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n628), .A2(new_n620), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n589), .A2(new_n618), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n561), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n387), .A2(KEYINPUT102), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n387), .A2(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(G1gat), .Z(G1324gat));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n561), .A2(new_n475), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n641), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G8gat), .B1(new_n650), .B2(new_n641), .ZN(new_n654));
  NOR2_X1   g453(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n655));
  MUX2_X1   g454(.A(KEYINPUT103), .B(new_n655), .S(new_n652), .Z(new_n656));
  AOI22_X1  g455(.A1(new_n653), .A2(new_n654), .B1(new_n651), .B2(new_n656), .ZN(G1325gat));
  INV_X1    g456(.A(new_n424), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n422), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(G15gat), .B1(new_n643), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n419), .ZN(new_n662));
  INV_X1    g461(.A(new_n421), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(G15gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n661), .B1(new_n643), .B2(new_n666), .ZN(G1326gat));
  NAND3_X1  g466(.A1(new_n561), .A2(new_n267), .A3(new_n642), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n618), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n589), .A2(new_n639), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n559), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n672), .B(new_n675), .C1(new_n489), .C2(new_n490), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n646), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(new_n500), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT45), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n618), .B1(new_n478), .B2(new_n488), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n266), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n264), .ZN(new_n685));
  INV_X1    g484(.A(new_n391), .ZN(new_n686));
  OAI22_X1  g485(.A1(new_n685), .A2(new_n686), .B1(new_n658), .B2(new_n422), .ZN(new_n687));
  INV_X1    g486(.A(new_n426), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n443), .A2(new_n444), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n689), .A2(new_n446), .A3(new_n440), .A4(new_n381), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT84), .B1(new_n449), .B2(KEYINPUT38), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n688), .B1(new_n692), .B2(new_n450), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n474), .B1(new_n473), .B2(new_n475), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n687), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT86), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n478), .A2(new_n479), .A3(new_n488), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n618), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n683), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n675), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n646), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n680), .B1(new_n705), .B2(new_n500), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n673), .A2(new_n501), .A3(new_n672), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n650), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n704), .B2(new_n467), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT46), .Z(new_n712));
  OAI211_X1 g511(.A(new_n710), .B(new_n711), .C1(new_n708), .C2(new_n712), .ZN(G1329gat));
  NOR3_X1   g512(.A1(new_n676), .A2(G43gat), .A3(new_n665), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n704), .A2(new_n660), .ZN(new_n716));
  INV_X1    g515(.A(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(KEYINPUT48), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n699), .A2(new_n700), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n702), .B1(new_n724), .B2(new_n672), .ZN(new_n725));
  INV_X1    g524(.A(new_n683), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n688), .B(new_n675), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G50gat), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n685), .A2(G50gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n677), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n723), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  INV_X1    g531(.A(new_n729), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n676), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n701), .A2(KEYINPUT107), .A3(new_n675), .A4(new_n729), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n723), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n703), .A2(new_n267), .A3(new_n675), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(G50gat), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT108), .B1(new_n731), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(G50gat), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n734), .A2(new_n723), .A3(new_n735), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n727), .A2(G50gat), .B1(new_n677), .B2(new_n729), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n742), .B(new_n743), .C1(new_n723), .C2(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n739), .A2(new_n745), .ZN(G1331gat));
  INV_X1    g545(.A(new_n589), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n747), .A2(new_n672), .A3(new_n559), .A4(new_n640), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n697), .B2(new_n698), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n646), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g550(.A(new_n749), .B(KEYINPUT109), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n467), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  NAND3_X1  g557(.A1(new_n752), .A2(G71gat), .A3(new_n659), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n749), .A2(new_n665), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(G71gat), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n752), .A2(new_n267), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n559), .A2(new_n589), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n703), .A2(new_n639), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n646), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n681), .A2(new_n765), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(KEYINPUT110), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n771));
  NAND3_X1  g570(.A1(new_n681), .A2(new_n765), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n595), .A3(new_n639), .A4(new_n678), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n767), .A2(new_n774), .ZN(G1336gat));
  AND4_X1   g574(.A1(new_n596), .A2(new_n773), .A3(new_n475), .A4(new_n639), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n703), .A2(new_n475), .A3(new_n639), .A4(new_n765), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(G92gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n778), .B(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n766), .B2(new_n660), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n665), .A2(G99gat), .A3(new_n640), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT112), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1338gat));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  INV_X1    g586(.A(G106gat), .ZN(new_n788));
  AND4_X1   g587(.A1(new_n788), .A2(new_n773), .A3(new_n688), .A4(new_n639), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n703), .A2(new_n267), .A3(new_n639), .A4(new_n765), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(G106gat), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n766), .A2(new_n426), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n788), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n787), .A2(new_n791), .B1(new_n792), .B2(new_n794), .ZN(G1339gat));
  NOR2_X1   g594(.A1(new_n641), .A2(new_n559), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n625), .A2(new_n626), .A3(new_n620), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n636), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n633), .B1(new_n627), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n638), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n798), .B2(new_n800), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n803), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n638), .A4(new_n801), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT93), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n542), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n811), .A2(new_n554), .A3(new_n556), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n534), .A2(new_n526), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n813), .A2(new_n528), .B1(new_n529), .B2(new_n527), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n548), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n809), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n558), .A2(KEYINPUT114), .A3(new_n815), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n808), .A2(new_n672), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n812), .A2(new_n816), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n808), .A2(new_n559), .B1(new_n639), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(new_n672), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n796), .B1(new_n822), .B2(new_n747), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n646), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n485), .ZN(new_n825));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n559), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT115), .B1(new_n823), .B2(new_n267), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n552), .B1(new_n536), .B2(new_n537), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n549), .B1(new_n828), .B2(new_n539), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n804), .B(new_n807), .C1(new_n829), .C2(new_n812), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n820), .A2(new_n639), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n672), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n818), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n804), .B(new_n807), .C1(new_n616), .C2(new_n617), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n747), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n796), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n839), .A3(new_n685), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n827), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n665), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n646), .A2(new_n475), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n559), .A2(G113gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n826), .B1(new_n846), .B2(new_n847), .ZN(G1340gat));
  AOI21_X1  g647(.A(G120gat), .B1(new_n825), .B2(new_n639), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n640), .A2(new_n349), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n846), .B2(new_n850), .ZN(G1341gat));
  OAI21_X1  g650(.A(G127gat), .B1(new_n845), .B2(new_n747), .ZN(new_n852));
  INV_X1    g651(.A(G127gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n825), .A2(new_n853), .A3(new_n589), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1342gat));
  OAI21_X1  g654(.A(G134gat), .B1(new_n845), .B2(new_n618), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n825), .A2(new_n342), .A3(new_n672), .ZN(new_n857));
  XOR2_X1   g656(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1343gat));
  NAND4_X1  g659(.A1(new_n824), .A2(new_n688), .A3(new_n467), .A4(new_n660), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n232), .A3(new_n559), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n823), .A2(KEYINPUT57), .A3(new_n426), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n802), .A2(new_n803), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n559), .A2(new_n865), .B1(new_n820), .B2(new_n639), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n819), .B1(new_n866), .B2(new_n672), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n796), .B1(new_n867), .B2(new_n747), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT57), .B1(new_n868), .B2(new_n685), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n659), .A2(new_n646), .A3(new_n475), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n864), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n559), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n863), .B1(new_n872), .B2(new_n232), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n234), .A3(new_n639), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n838), .A2(KEYINPUT57), .A3(new_n688), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT117), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n672), .A2(new_n865), .A3(new_n817), .A4(new_n818), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n866), .B2(new_n672), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n589), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n837), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n884), .B2(new_n267), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n639), .B(new_n870), .C1(new_n878), .C2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n876), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n234), .C1(new_n871), .C2(new_n639), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n875), .B1(new_n887), .B2(new_n888), .ZN(G1345gat));
  OR3_X1    g688(.A1(new_n861), .A2(KEYINPUT119), .A3(new_n747), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n861), .B2(new_n747), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n227), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n871), .A2(G155gat), .A3(new_n589), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT120), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n862), .B2(new_n672), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n618), .A2(new_n228), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n871), .B2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n678), .A2(new_n467), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n823), .A2(new_n480), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n559), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n839), .B1(new_n838), .B2(new_n685), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT115), .B(new_n267), .C1(new_n836), .C2(new_n837), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n664), .B(new_n899), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n559), .A2(G169gat), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(G1348gat));
  OAI21_X1  g707(.A(G176gat), .B1(new_n905), .B2(new_n640), .ZN(new_n909));
  INV_X1    g708(.A(G176gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n901), .A2(new_n910), .A3(new_n639), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(G1349gat));
  OAI21_X1  g711(.A(G183gat), .B1(new_n905), .B2(new_n747), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n589), .A2(new_n285), .A3(new_n287), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT121), .B1(new_n901), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n841), .A2(new_n664), .A3(new_n672), .A4(new_n899), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT122), .B1(new_n919), .B2(G190gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G190gat), .B1(new_n905), .B2(new_n618), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(KEYINPUT123), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n922), .A2(KEYINPUT61), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n918), .B(new_n929), .C1(new_n920), .C2(new_n921), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n901), .A2(new_n288), .A3(new_n672), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n900), .A2(new_n659), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n823), .A2(new_n934), .A3(new_n426), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n559), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n878), .B2(new_n885), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n560), .A2(new_n545), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  OAI21_X1  g739(.A(G204gat), .B1(new_n937), .B2(new_n640), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(new_n209), .A3(new_n639), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(KEYINPUT124), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g744(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n941), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT125), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n941), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1353gat));
  OAI21_X1  g751(.A(G211gat), .B1(new_n937), .B2(new_n747), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT63), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(KEYINPUT63), .ZN(new_n955));
  INV_X1    g754(.A(new_n935), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(G211gat), .A3(new_n747), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(G1354gat));
  AOI21_X1  g758(.A(G218gat), .B1(new_n935), .B2(new_n672), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n672), .A2(new_n213), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n961), .B(KEYINPUT127), .Z(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n938), .B2(new_n962), .ZN(G1355gat));
endmodule


