//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209));
  XOR2_X1   g008(.A(G141gat), .B(G148gat), .Z(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT2), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n210), .A2(new_n213), .B1(new_n214), .B2(KEYINPUT74), .ZN(new_n215));
  INV_X1    g014(.A(new_n214), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT74), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n216), .A2(new_n210), .A3(new_n217), .A4(new_n213), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n208), .B1(new_n209), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n203), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n206), .B(new_n207), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n219), .A2(new_n220), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT76), .A3(new_n224), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G225gat), .A2(G233gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(new_n227), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n221), .A2(new_n227), .A3(KEYINPUT4), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n228), .A2(new_n208), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n233), .ZN(new_n242));
  INV_X1    g041(.A(new_n232), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT0), .ZN(new_n248));
  XNOR2_X1  g047(.A(G57gat), .B(G85gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n237), .B1(new_n226), .B2(new_n230), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT5), .A3(new_n232), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT6), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n250), .B(KEYINPUT79), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AND4_X1   g057(.A1(KEYINPUT5), .A2(new_n231), .A3(new_n232), .A4(new_n238), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n244), .B1(new_n251), .B2(new_n232), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT81), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT81), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n262), .A3(new_n252), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n258), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n252), .ZN(new_n267));
  INV_X1    g066(.A(new_n250), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT6), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n256), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT67), .B1(new_n273), .B2(G183gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT27), .B(G183gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n272), .B(new_n274), .C1(new_n275), .C2(KEYINPUT67), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(KEYINPUT28), .A3(new_n272), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(new_n272), .ZN(new_n282));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT26), .ZN(new_n286));
  AOI211_X1 g085(.A(new_n282), .B(new_n286), .C1(KEYINPUT26), .C2(new_n285), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n285), .A2(KEYINPUT23), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n290), .A2(G169gat), .A3(G176gat), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n289), .A2(new_n291), .A3(new_n284), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n281), .B2(new_n272), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n294), .B(new_n295), .C1(G183gat), .C2(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n295), .B(new_n300), .ZN(new_n301));
  OR3_X1    g100(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n292), .B(KEYINPUT25), .C1(new_n301), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n208), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n306), .A3(new_n227), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G227gat), .ZN(new_n311));
  INV_X1    g110(.A(G233gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n271), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n310), .A2(new_n271), .A3(new_n313), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT32), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT33), .B1(new_n315), .B2(new_n316), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n308), .B(new_n309), .C1(new_n311), .C2(new_n312), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT34), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(G15gat), .B(G43gat), .Z(new_n323));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n319), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n320), .B(KEYINPUT34), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT33), .ZN(new_n329));
  INV_X1    g128(.A(new_n316), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(new_n314), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n331), .B2(new_n325), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n318), .B1(new_n327), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n322), .B1(new_n319), .B2(new_n326), .ZN(new_n334));
  INV_X1    g133(.A(new_n318), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n328), .A3(new_n325), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G228gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(new_n312), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n224), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G197gat), .B(G204gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(G211gat), .A2(G218gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT22), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(KEYINPUT70), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT70), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G211gat), .B(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n350), .A2(KEYINPUT71), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(new_n350), .B2(KEYINPUT71), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n343), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n352), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n351), .B1(new_n348), .B2(new_n349), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n342), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n221), .B1(new_n359), .B2(new_n223), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n341), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n353), .A2(new_n354), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(KEYINPUT72), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n343), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n340), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(KEYINPUT77), .A3(new_n342), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n342), .A3(new_n354), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT3), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n221), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n361), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G22gat), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n375), .B(new_n361), .C1(new_n367), .C2(new_n372), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n373), .B2(G22gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT31), .B(G50gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n377), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n374), .A2(new_n378), .A3(new_n376), .A4(new_n382), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n307), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT73), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n307), .A2(KEYINPUT73), .A3(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n307), .A2(new_n342), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n387), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n355), .B(new_n364), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n362), .A3(new_n389), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n363), .A2(new_n365), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n393), .B2(new_n395), .ZN(new_n406));
  INV_X1    g205(.A(new_n402), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(KEYINPUT30), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n406), .A2(new_n407), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n401), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT35), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n338), .A2(new_n386), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n202), .B1(new_n270), .B2(new_n414), .ZN(new_n415));
  AND4_X1   g214(.A1(new_n386), .A2(new_n413), .A3(new_n337), .A4(new_n333), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n261), .A2(new_n263), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n265), .B1(new_n417), .B2(new_n257), .ZN(new_n418));
  AOI211_X1 g217(.A(KEYINPUT82), .B(new_n258), .C1(new_n261), .C2(new_n263), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n269), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n255), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n421), .A3(KEYINPUT84), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n269), .A2(new_n253), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n423), .A2(new_n255), .B1(new_n409), .B2(new_n412), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n338), .A2(new_n386), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT35), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n415), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n401), .A2(KEYINPUT38), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n362), .B1(new_n395), .B2(new_n389), .ZN(new_n431));
  INV_X1    g230(.A(new_n396), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n405), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n429), .B(new_n430), .C1(new_n428), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n403), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n404), .B1(new_n410), .B2(new_n428), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT83), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(new_n404), .C1(new_n410), .C2(new_n428), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n439), .A3(new_n429), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(KEYINPUT38), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n255), .A3(new_n420), .ZN(new_n442));
  INV_X1    g241(.A(new_n386), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n251), .A2(new_n232), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT39), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n257), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n242), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n448), .B2(new_n232), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n251), .B2(new_n232), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n444), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n451), .A2(new_n452), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n409), .A2(new_n412), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n443), .B1(new_n456), .B2(new_n266), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT69), .B(KEYINPUT36), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n333), .A2(new_n337), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT69), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n333), .A2(new_n337), .B1(new_n462), .B2(KEYINPUT36), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n423), .A2(new_n255), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n455), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n443), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n458), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n427), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G169gat), .B(G197gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT12), .Z(new_n477));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(G29gat), .B2(G36gat), .ZN(new_n479));
  INV_X1    g278(.A(G29gat), .ZN(new_n480));
  INV_X1    g279(.A(G36gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT14), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT87), .B(G29gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n479), .B(new_n482), .C1(new_n483), .C2(new_n481), .ZN(new_n484));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n488));
  INV_X1    g287(.A(G50gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(KEYINPUT88), .A2(G43gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n491), .A2(new_n492), .B1(new_n485), .B2(KEYINPUT15), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n487), .B1(new_n493), .B2(new_n484), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n495), .A2(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(KEYINPUT17), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n493), .A2(new_n484), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(new_n495), .A3(KEYINPUT17), .A4(new_n487), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  XOR2_X1   g301(.A(G15gat), .B(G22gat), .Z(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G1gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505));
  INV_X1    g304(.A(G1gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT16), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT90), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT89), .B1(new_n504), .B2(new_n507), .ZN(new_n509));
  INV_X1    g308(.A(G8gat), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n502), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n507), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(KEYINPUT89), .A3(G8gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT92), .B1(new_n501), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n494), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n511), .A2(new_n515), .A3(KEYINPUT93), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT93), .B1(new_n511), .B2(new_n515), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n498), .A2(new_n500), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n511), .A4(new_n515), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n517), .A2(new_n521), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n522), .B(KEYINPUT13), .Z(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n519), .A2(new_n520), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n494), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n534), .B2(new_n521), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT86), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n477), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n530), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n540));
  INV_X1    g339(.A(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n477), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT86), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n211), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n520), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n511), .A2(new_n515), .A3(KEYINPUT93), .ZN(new_n551));
  NAND2_X1  g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(G71gat), .A2(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT9), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(KEYINPUT95), .A2(G57gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G64gat), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n559));
  AND2_X1   g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n552), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(new_n553), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n556), .A2(new_n558), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n550), .A2(new_n551), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT96), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n533), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n549), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n572));
  AND2_X1   g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G127gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n567), .A2(new_n569), .A3(new_n549), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n571), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n575), .B(new_n576), .ZN(new_n581));
  INV_X1    g380(.A(new_n579), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n570), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT97), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT7), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT8), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT8), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(G99gat), .B2(G106gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT97), .B(G85gat), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n604), .B1(new_n605), .B2(new_n590), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n600), .A3(new_n596), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n585), .B1(new_n494), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n523), .B2(new_n608), .ZN(new_n610));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT98), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n610), .A2(KEYINPUT99), .A3(new_n612), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT99), .B1(new_n610), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT100), .B1(new_n614), .B2(new_n615), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  OAI221_X1 g421(.A(new_n613), .B1(KEYINPUT100), .B2(new_n622), .C1(new_n614), .C2(new_n615), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n558), .A2(new_n556), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n561), .A2(new_n563), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n600), .B1(new_n606), .B2(new_n596), .ZN(new_n629));
  AND4_X1   g428(.A1(new_n600), .A2(new_n591), .A3(new_n596), .A4(new_n598), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n564), .A2(new_n602), .A3(new_n607), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(KEYINPUT101), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n602), .A2(new_n564), .A3(new_n607), .A4(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT10), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n625), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n633), .A2(G230gat), .A3(G233gat), .A4(new_n635), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  NOR2_X1   g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n584), .A2(new_n624), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n546), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n471), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n466), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n506), .ZN(G1324gat));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT16), .B(G8gat), .Z(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n468), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(G8gat), .B1(new_n650), .B2(new_n455), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n658), .A2(new_n660), .A3(KEYINPUT102), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT102), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(G1325gat));
  INV_X1    g462(.A(new_n338), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n650), .A2(G15gat), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n650), .B2(new_n465), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n386), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT103), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n624), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n471), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n647), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n545), .A2(new_n584), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n467), .A3(new_n483), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n461), .A2(new_n463), .B1(new_n386), .B2(new_n424), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n442), .B2(new_n457), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n416), .A2(new_n421), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n682), .A2(new_n202), .B1(KEYINPUT35), .B2(new_n425), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n683), .B2(new_n422), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n684), .A2(new_n685), .A3(new_n624), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n471), .B2(new_n672), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n687), .A3(new_n676), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n466), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n679), .B1(new_n483), .B2(new_n690), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n677), .A2(new_n481), .A3(new_n468), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT46), .Z(new_n693));
  OAI21_X1  g492(.A(G36gat), .B1(new_n689), .B2(new_n455), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1329gat));
  OAI21_X1  g494(.A(new_n685), .B1(new_n684), .B2(new_n624), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n471), .A2(KEYINPUT44), .A3(new_n672), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n696), .A2(new_n464), .A3(new_n697), .A4(new_n675), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n488), .A2(new_n490), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT47), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n677), .A2(new_n338), .A3(new_n488), .A4(new_n490), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n700), .B(new_n703), .C1(new_n701), .C2(KEYINPUT47), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1330gat));
  AOI21_X1  g506(.A(new_n489), .B1(new_n688), .B2(new_n443), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n386), .A2(G50gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n677), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(KEYINPUT48), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  INV_X1    g513(.A(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n708), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n584), .ZN(new_n718));
  NOR4_X1   g517(.A1(new_n546), .A2(new_n672), .A3(new_n718), .A4(new_n647), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n471), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n467), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g522(.A1(new_n720), .A2(new_n455), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  AND2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n724), .B2(new_n725), .ZN(G1333gat));
  INV_X1    g527(.A(G71gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n720), .B2(new_n664), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n465), .A2(new_n729), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n721), .A2(KEYINPUT106), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT106), .B1(new_n721), .B2(new_n731), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n721), .A2(new_n443), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g536(.A1(new_n684), .A2(new_n624), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n546), .A2(new_n584), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT51), .A4(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n471), .A2(KEYINPUT51), .A3(new_n672), .A4(new_n740), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT107), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  INV_X1    g543(.A(new_n740), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n673), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n741), .A2(new_n746), .A3(new_n743), .A4(KEYINPUT108), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n674), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n467), .A2(new_n605), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n686), .A2(new_n687), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n745), .A2(new_n647), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n466), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n751), .A2(new_n752), .B1(new_n605), .B2(new_n756), .ZN(G1336gat));
  NOR3_X1   g556(.A1(new_n455), .A2(G92gat), .A3(new_n647), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n747), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n696), .A2(new_n468), .A3(new_n697), .A4(new_n754), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(new_n760), .B2(G92gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n760), .A2(new_n763), .A3(G92gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n760), .B2(G92gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n758), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n746), .B2(new_n742), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n762), .B1(new_n768), .B2(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n755), .B2(new_n465), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n753), .A2(KEYINPUT110), .A3(new_n464), .A4(new_n754), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(G99gat), .A3(new_n773), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n664), .A2(G99gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n751), .B2(new_n775), .ZN(G1338gat));
  NOR3_X1   g575(.A1(new_n386), .A2(G106gat), .A3(new_n647), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n747), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n696), .A2(new_n443), .A3(new_n697), .A4(new_n754), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G106gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n746), .A2(new_n742), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n783), .A2(new_n777), .B1(new_n779), .B2(G106gat), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n778), .A2(new_n782), .B1(new_n784), .B2(new_n781), .ZN(G1339gat));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  INV_X1    g585(.A(new_n646), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n788), .B(new_n625), .C1(new_n636), .C2(new_n638), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  INV_X1    g589(.A(new_n644), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n636), .A2(new_n625), .A3(new_n638), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(KEYINPUT54), .A3(new_n639), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT55), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n787), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n789), .A2(new_n791), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT112), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n802), .B2(new_n796), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n786), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n639), .A2(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(new_n795), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n646), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n796), .B1(new_n792), .B2(new_n793), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n805), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n810), .A3(KEYINPUT113), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n804), .A2(new_n538), .A3(new_n544), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n521), .A2(new_n525), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n522), .B1(new_n814), .B2(new_n517), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n534), .A2(new_n521), .A3(new_n532), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n476), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n674), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n672), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n817), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n624), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n821), .A2(new_n804), .A3(new_n811), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n718), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n648), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT111), .B1(new_n824), .B2(new_n546), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n648), .A2(new_n545), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n823), .A2(KEYINPUT114), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n338), .A2(new_n386), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n466), .A2(new_n468), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n546), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n833), .B2(new_n443), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n823), .A2(KEYINPUT114), .A3(new_n828), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT114), .B1(new_n823), .B2(new_n828), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n386), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n836), .A2(new_n664), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n546), .A2(G113gat), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n838), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  AOI21_X1  g650(.A(G120gat), .B1(new_n837), .B2(new_n674), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n674), .A2(G120gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n849), .B2(new_n853), .ZN(G1341gat));
  AND2_X1   g653(.A1(new_n584), .A2(G127gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n845), .A2(new_n847), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n856), .A2(new_n857), .ZN(new_n859));
  AOI21_X1  g658(.A(G127gat), .B1(new_n837), .B2(new_n584), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n837), .A2(new_n862), .A3(new_n672), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n846), .A2(new_n624), .A3(new_n848), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n862), .ZN(G1343gat));
  INV_X1    g666(.A(G141gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n831), .A2(new_n443), .A3(new_n832), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n465), .A2(new_n835), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n868), .B1(new_n873), .B2(new_n545), .ZN(new_n874));
  INV_X1    g673(.A(new_n818), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n798), .A2(new_n803), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n546), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n672), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n718), .B1(new_n878), .B2(new_n822), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n828), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n386), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n870), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n872), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n545), .A2(new_n868), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n874), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n874), .B(KEYINPUT58), .C1(new_n887), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1344gat));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n674), .ZN(new_n895));
  OR3_X1    g694(.A1(new_n869), .A2(G148gat), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n831), .A2(new_n443), .A3(new_n832), .A4(new_n885), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n821), .A2(new_n876), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n877), .B2(new_n672), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n900), .A2(new_n718), .B1(new_n545), .B2(new_n648), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n881), .B1(new_n901), .B2(new_n386), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n895), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(G148gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n903), .B2(new_n904), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n897), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n897), .A2(G148gat), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n869), .A2(new_n884), .B1(new_n880), .B2(new_n882), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n871), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n911), .B2(new_n674), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n896), .B1(new_n908), .B2(new_n912), .ZN(G1345gat));
  NAND2_X1  g712(.A1(new_n584), .A2(G155gat), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT119), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n870), .A2(new_n584), .A3(new_n872), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n911), .A2(new_n915), .B1(new_n211), .B2(new_n916), .ZN(G1346gat));
  NOR3_X1   g716(.A1(new_n910), .A2(new_n624), .A3(new_n871), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G162gat), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n672), .A2(new_n212), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n873), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT120), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n923), .A2(KEYINPUT120), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n920), .A2(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n834), .A2(new_n455), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT122), .Z(new_n928));
  NAND3_X1  g727(.A1(new_n843), .A2(new_n466), .A3(new_n928), .ZN(new_n929));
  OR3_X1    g728(.A1(new_n929), .A2(G169gat), .A3(new_n545), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n467), .A2(new_n455), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n932), .A2(new_n664), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n845), .A2(new_n546), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT123), .B1(new_n934), .B2(G169gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  INV_X1    g736(.A(new_n929), .ZN(new_n938));
  INV_X1    g737(.A(G176gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n674), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n845), .A2(new_n674), .A3(new_n933), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n939), .ZN(G1349gat));
  XNOR2_X1  g741(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT115), .B1(new_n843), .B2(new_n386), .ZN(new_n944));
  NOR4_X1   g743(.A1(new_n841), .A2(new_n842), .A3(new_n839), .A4(new_n443), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n584), .B(new_n933), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G183gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n584), .A2(new_n275), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n929), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n943), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n943), .ZN(new_n952));
  AOI211_X1 g751(.A(new_n949), .B(new_n952), .C1(new_n946), .C2(G183gat), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n953), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n272), .A3(new_n672), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n845), .A2(new_n672), .A3(new_n933), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NOR2_X1   g759(.A1(new_n833), .A2(new_n467), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n464), .A2(new_n386), .A3(new_n455), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n545), .A2(G197gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT125), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n932), .A2(new_n464), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n967), .B1(new_n898), .B2(new_n902), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(G197gat), .B1(new_n969), .B2(new_n545), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n965), .A2(new_n970), .ZN(G1352gat));
  NAND3_X1  g770(.A1(new_n843), .A2(new_n466), .A3(new_n962), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n647), .A2(G204gat), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(KEYINPUT62), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n961), .A2(new_n976), .A3(new_n962), .A4(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(G204gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n979), .B1(new_n968), .B2(new_n674), .ZN(new_n980));
  OR3_X1    g779(.A1(new_n978), .A2(new_n980), .A3(KEYINPUT126), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT126), .B1(new_n978), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1353gat));
  OR3_X1    g782(.A1(new_n972), .A2(G211gat), .A3(new_n718), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n584), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1354gat));
  INV_X1    g787(.A(G218gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n989), .B1(new_n972), .B2(new_n624), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n968), .A2(G218gat), .A3(new_n672), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(G1355gat));
endmodule


