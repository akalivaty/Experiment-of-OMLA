//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  AOI21_X1  g007(.A(G128), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(KEYINPUT1), .A3(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n194), .A2(KEYINPUT85), .A3(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n198), .B2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT85), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(new_n193), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n201), .A2(KEYINPUT1), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(new_n200), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n206), .A2(G107), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n207), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n205), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT10), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT0), .B(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(new_n198), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n198), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n201), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n211), .A2(new_n214), .A3(new_n207), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(G101), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(G101), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n216), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n231), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT66), .B1(new_n239), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  OAI211_X1 g057(.A(KEYINPUT66), .B(new_n243), .C1(new_n239), .C2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G134), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n242), .A3(new_n244), .A4(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n246), .B1(new_n240), .B2(KEYINPUT11), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n242), .B1(new_n250), .B2(new_n244), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n238), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n244), .A3(new_n247), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n248), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n201), .A2(new_n202), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT67), .B1(new_n257), .B2(new_n195), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n194), .A2(new_n259), .A3(new_n196), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n204), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n221), .A2(new_n237), .A3(new_n256), .A4(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G140), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n265), .A2(G227), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n261), .A2(new_n218), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n203), .B1(KEYINPUT85), .B2(new_n199), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n217), .B1(new_n273), .B2(new_n197), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n271), .B1(new_n275), .B2(new_n256), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n271), .B1(new_n254), .B2(new_n248), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n272), .B2(new_n274), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT86), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(KEYINPUT86), .B(new_n277), .C1(new_n272), .C2(new_n274), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n270), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n262), .A2(new_n237), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n274), .A2(KEYINPUT10), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n255), .B(new_n252), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n263), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n267), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n189), .B1(new_n289), .B2(new_n187), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n269), .A2(KEYINPUT87), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT87), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n263), .A2(new_n292), .A3(new_n268), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n286), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n282), .A2(new_n263), .ZN(new_n295));
  OAI211_X1 g109(.A(G469), .B(new_n294), .C1(new_n295), .C2(new_n268), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(KEYINPUT84), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G113), .B(G122), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(new_n206), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n265), .A3(G214), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n307));
  AOI21_X1  g121(.A(G143), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n305), .A2(new_n265), .A3(KEYINPUT88), .A4(G214), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n306), .A2(new_n192), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n309), .B1(new_n308), .B2(new_n310), .ZN(new_n314));
  OAI21_X1  g128(.A(G131), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n314), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(new_n242), .A3(new_n312), .A4(new_n311), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT17), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT79), .A4(KEYINPUT16), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n321), .B2(KEYINPUT16), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n324), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G146), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n190), .B(new_n324), .C1(new_n325), .C2(new_n327), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n319), .B(new_n331), .C1(new_n318), .C2(new_n315), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT18), .B(G131), .C1(new_n313), .C2(new_n314), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT18), .A2(G131), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n316), .A2(new_n334), .A3(new_n312), .A4(new_n311), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n321), .A2(new_n323), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(G146), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(G146), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n335), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n304), .B1(new_n332), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n331), .B1(new_n315), .B2(new_n318), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n304), .B(new_n341), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n188), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G475), .ZN(new_n348));
  NOR2_X1   g162(.A1(G475), .A2(G902), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n304), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n333), .A2(new_n335), .A3(new_n340), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n337), .B(KEYINPUT19), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n329), .B1(G146), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n315), .B2(new_n317), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n351), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n350), .B1(new_n345), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n345), .A2(new_n356), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT91), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT91), .ZN(new_n362));
  AND4_X1   g176(.A1(new_n362), .A2(new_n358), .A3(new_n360), .A4(new_n349), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n348), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G952), .ZN(new_n366));
  AOI211_X1 g180(.A(G953), .B(new_n366), .C1(G234), .C2(G237), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT21), .B(G898), .Z(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT97), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI211_X1 g184(.A(new_n188), .B(new_n265), .C1(G234), .C2(G237), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n192), .A2(G128), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT13), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT92), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n202), .A2(G143), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n374), .A2(KEYINPUT92), .A3(new_n375), .ZN(new_n380));
  OAI21_X1  g194(.A(G134), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n377), .A3(new_n239), .ZN(new_n382));
  XNOR2_X1  g196(.A(G116), .B(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n213), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n383), .A2(new_n213), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n381), .B(new_n382), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n374), .A2(new_n377), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G134), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT93), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n382), .A2(new_n389), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(KEYINPUT93), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n395));
  INV_X1    g209(.A(G122), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n213), .B1(new_n397), .B2(KEYINPUT14), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(new_n394), .B2(new_n398), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n391), .B(new_n392), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G217), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n298), .A2(new_n402), .A3(G953), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n387), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n387), .B2(new_n401), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n188), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT95), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G478), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT15), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT95), .B(new_n188), .C1(new_n404), .C2(new_n405), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n413));
  OR3_X1    g227(.A1(new_n406), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n406), .B2(new_n410), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n365), .A2(new_n373), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G214), .B1(G237), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G210), .B1(G237), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G224), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n259), .B1(new_n194), .B2(new_n196), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT67), .B(new_n195), .C1(new_n198), .C2(G128), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n203), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n322), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n230), .A2(G125), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n425), .A3(new_n430), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(G116), .B(G119), .Z(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT2), .B(G113), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n236), .A3(new_n234), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n435), .A2(new_n436), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n440));
  INV_X1    g254(.A(G119), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(G116), .ZN(new_n442));
  OAI211_X1 g256(.A(G113), .B(new_n442), .C1(new_n435), .C2(new_n440), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n218), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n438), .A2(new_n446), .A3(new_n444), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n451), .A3(new_n447), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n434), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n432), .B2(new_n433), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n429), .A2(new_n430), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n455), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n443), .A2(new_n439), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n217), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n444), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n446), .B(KEYINPUT8), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n449), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n188), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n422), .B1(new_n454), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n464), .ZN(new_n467));
  INV_X1    g281(.A(new_n433), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n468), .A2(new_n431), .B1(KEYINPUT7), .B2(new_n424), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n421), .A3(new_n453), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n420), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n302), .A2(new_n418), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT74), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT28), .ZN(new_n476));
  INV_X1    g290(.A(new_n437), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n252), .A2(new_n255), .A3(new_n231), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n239), .A2(G137), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n479), .B2(new_n246), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n248), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n261), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n437), .B1(new_n261), .B2(new_n482), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n485), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n486), .B1(new_n485), .B2(new_n478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n484), .B1(new_n489), .B2(KEYINPUT73), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT73), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n487), .B2(new_n488), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n476), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT28), .B1(new_n485), .B2(new_n478), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n305), .A2(new_n265), .A3(G210), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT27), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT26), .B(G101), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n495), .A2(KEYINPUT29), .A3(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n475), .B(new_n188), .C1(new_n493), .C2(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n252), .A2(new_n231), .A3(new_n255), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n477), .B1(new_n428), .B2(new_n481), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT69), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n485), .A2(new_n478), .A3(new_n486), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(KEYINPUT73), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n484), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n492), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n500), .B1(new_n508), .B2(KEYINPUT28), .ZN(new_n509));
  OAI21_X1  g323(.A(KEYINPUT74), .B1(new_n509), .B2(G902), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n230), .B1(new_n254), .B2(new_n248), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n426), .A2(new_n427), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n481), .B1(new_n512), .B2(new_n204), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n437), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n489), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n499), .B(new_n495), .C1(new_n515), .C2(new_n476), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n478), .A2(KEYINPUT30), .A3(new_n483), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n511), .B2(new_n513), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n437), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n489), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n499), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT29), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n501), .A2(new_n510), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G472), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n520), .A2(new_n504), .A3(new_n505), .A4(new_n499), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT70), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n489), .A2(new_n529), .A3(new_n520), .A4(new_n499), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(KEYINPUT31), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n476), .B1(new_n489), .B2(new_n514), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n522), .B1(new_n532), .B2(new_n494), .ZN(new_n533));
  AND4_X1   g347(.A1(new_n520), .A2(new_n504), .A3(new_n505), .A4(new_n499), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT71), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT71), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n527), .A2(new_n537), .A3(KEYINPUT31), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n531), .B(new_n533), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n526), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G234), .ZN(new_n547));
  OAI21_X1  g361(.A(G217), .B1(new_n547), .B2(G902), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n202), .A2(G119), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n441), .A2(G128), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT76), .B1(new_n441), .B2(G128), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT24), .B(G110), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n329), .B2(new_n330), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT77), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT77), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(new_n562), .A3(KEYINPUT23), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n551), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n202), .A2(KEYINPUT78), .A3(G119), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n561), .A2(new_n563), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G110), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G110), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n572), .A3(new_n568), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n556), .A2(new_n557), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT80), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n337), .A2(G146), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n328), .B2(G146), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n571), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT22), .B(G137), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n188), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n575), .A2(new_n578), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT80), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n588), .A2(new_n589), .B1(new_n570), .B2(new_n559), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT81), .B1(new_n590), .B2(new_n584), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT81), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n592), .A3(new_n585), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n586), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n550), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g411(.A(new_n595), .B(new_n586), .C1(new_n591), .C2(new_n593), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n549), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT83), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(KEYINPUT83), .B(new_n549), .C1(new_n597), .C2(new_n598), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n591), .A2(new_n593), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n581), .B2(new_n585), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n548), .A2(new_n188), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n474), .A2(new_n546), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT98), .B(G101), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G3));
  INV_X1    g424(.A(new_n542), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n539), .A2(new_n188), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(G472), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n302), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n613), .A2(new_n607), .A3(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n404), .A2(new_n405), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT33), .B1(new_n616), .B2(KEYINPUT99), .ZN(new_n617));
  OAI211_X1 g431(.A(KEYINPUT99), .B(KEYINPUT33), .C1(new_n404), .C2(new_n405), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(G478), .B(new_n188), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n364), .A2(new_n472), .A3(new_n373), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT100), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n372), .B(new_n420), .C1(new_n466), .C2(new_n471), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n364), .A4(new_n622), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n615), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  XNOR2_X1  g445(.A(new_n357), .B(new_n360), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n632), .A2(new_n348), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n615), .A2(new_n416), .A3(new_n625), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NOR2_X1   g450(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n581), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n188), .A3(new_n548), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT101), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n601), .A2(new_n602), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT102), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n601), .A2(new_n643), .A3(new_n602), .A4(new_n640), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n474), .A2(new_n642), .A3(new_n613), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT37), .B(G110), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT103), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n645), .B(new_n648), .ZN(G12));
  AND2_X1   g463(.A1(new_n642), .A2(new_n644), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n611), .B2(KEYINPUT32), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n302), .B1(new_n652), .B2(new_n526), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n632), .A2(new_n348), .A3(new_n416), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n371), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n367), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n473), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n650), .A2(KEYINPUT105), .A3(new_n653), .A4(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n642), .A2(new_n546), .A3(new_n614), .A4(new_n644), .ZN(new_n663));
  INV_X1    g477(.A(new_n660), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  NAND2_X1  g481(.A1(new_n466), .A2(new_n471), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT38), .Z(new_n669));
  NOR2_X1   g483(.A1(new_n417), .A2(new_n420), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n364), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n658), .B(KEYINPUT39), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n302), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n669), .B(new_n671), .C1(new_n675), .C2(KEYINPUT40), .ZN(new_n676));
  INV_X1    g490(.A(new_n641), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n528), .A2(new_n530), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n522), .B2(new_n508), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n679), .B2(G902), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n652), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n677), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  NAND3_X1  g498(.A1(new_n364), .A2(new_n622), .A3(new_n658), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n473), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n653), .A2(new_n642), .A3(new_n644), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  AND2_X1   g502(.A1(new_n546), .A2(new_n607), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n289), .A2(new_n187), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n289), .A2(new_n187), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n301), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n624), .B2(new_n627), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  INV_X1    g510(.A(new_n625), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n692), .A2(new_n697), .A3(new_n654), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NAND4_X1  g514(.A1(new_n690), .A2(new_n472), .A3(new_n301), .A4(new_n691), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n418), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n642), .A2(new_n546), .A3(new_n702), .A4(new_n644), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  NAND3_X1  g518(.A1(new_n670), .A2(new_n364), .A3(new_n668), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n692), .A3(new_n372), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n494), .B1(new_n508), .B2(KEYINPUT28), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n531), .B1(new_n707), .B2(new_n499), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(KEYINPUT106), .B(new_n531), .C1(new_n707), .C2(new_n499), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n710), .B(new_n711), .C1(new_n536), .C2(new_n538), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n540), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n612), .A2(G472), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n706), .A2(new_n713), .A3(new_n607), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  AND2_X1   g530(.A1(new_n713), .A2(new_n714), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n701), .A2(new_n685), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n641), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  XOR2_X1   g534(.A(new_n189), .B(KEYINPUT107), .Z(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n289), .B2(new_n187), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n296), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n668), .A2(new_n420), .A3(new_n300), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n685), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n546), .A2(new_n727), .A3(new_n607), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n546), .A2(new_n607), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n611), .A2(KEYINPUT32), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n541), .A3(new_n526), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(KEYINPUT42), .A3(new_n607), .A4(new_n727), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NOR3_X1   g552(.A1(new_n726), .A2(new_n654), .A3(new_n659), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n546), .A3(new_n607), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NAND2_X1  g555(.A1(new_n365), .A2(new_n622), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT43), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n742), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n613), .A2(new_n677), .A3(KEYINPUT110), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT110), .B1(new_n613), .B2(new_n677), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n294), .B1(new_n295), .B2(new_n268), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n187), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n759), .B1(new_n765), .B2(new_n722), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n721), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n691), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n768), .A2(new_n301), .A3(new_n672), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n668), .A2(new_n420), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n756), .B2(new_n752), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n758), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  INV_X1    g588(.A(new_n770), .ZN(new_n775));
  OR3_X1    g589(.A1(new_n607), .A2(new_n685), .A3(new_n775), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n776), .A2(KEYINPUT113), .A3(new_n546), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT113), .B1(new_n776), .B2(new_n546), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n768), .A2(new_n301), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n768), .A2(new_n301), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  NAND2_X1  g601(.A1(new_n690), .A2(new_n691), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n301), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n607), .A2(new_n717), .A3(new_n367), .A4(new_n747), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(new_n770), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n791), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n692), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n669), .A2(new_n797), .A3(new_n420), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT50), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n652), .A2(new_n607), .A3(new_n680), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n692), .A2(new_n775), .A3(new_n657), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n364), .A2(new_n622), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n747), .A2(new_n804), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT119), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n717), .A2(new_n641), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n796), .A2(KEYINPUT51), .A3(new_n802), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n802), .A2(new_n811), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n790), .A2(new_n794), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n735), .A2(new_n607), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n809), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT48), .Z(new_n819));
  NAND3_X1  g633(.A1(new_n793), .A2(new_n472), .A3(new_n797), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n366), .A2(G953), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n364), .A2(new_n622), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n805), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n812), .A2(new_n816), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n546), .B(new_n607), .C1(new_n693), .C2(new_n698), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n703), .A3(new_n715), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n365), .A2(new_n416), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n697), .B1(new_n828), .B2(new_n822), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n613), .A2(new_n607), .A3(new_n829), .A4(new_n614), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n645), .A2(new_n608), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n713), .A2(new_n727), .A3(new_n714), .A4(new_n641), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n633), .A2(new_n770), .A3(new_n417), .A4(new_n658), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n740), .B(new_n833), .C1(new_n663), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n832), .A2(new_n737), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n661), .A2(new_n665), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n658), .B(KEYINPUT116), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n724), .A2(new_n301), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n677), .A2(KEYINPUT117), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n724), .A2(new_n301), .A3(new_n840), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n641), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n705), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n842), .A2(new_n681), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n719), .A2(new_n687), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n838), .A2(new_n839), .A3(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n719), .A2(new_n687), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(new_n850), .B2(new_n666), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n837), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n839), .B1(new_n838), .B2(new_n848), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n850), .A2(KEYINPUT52), .A3(new_n666), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n857), .B2(new_n837), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n827), .A2(KEYINPUT118), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n826), .A2(new_n861), .A3(new_n703), .A4(new_n715), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n835), .B1(new_n733), .B2(new_n736), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n831), .A2(new_n853), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n852), .A2(new_n853), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n825), .A2(new_n870), .B1(G952), .B2(G953), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT114), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n669), .A2(new_n874), .A3(new_n419), .A4(new_n301), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n742), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n803), .A3(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT115), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n878), .ZN(G75));
  NAND2_X1  g693(.A1(new_n450), .A2(new_n452), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n434), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT55), .Z(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(G210), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n188), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n855), .B2(new_n856), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n858), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(KEYINPUT121), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n890), .B(new_n885), .C1(new_n858), .C2(new_n887), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n265), .A2(G952), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n888), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT122), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n885), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT121), .B1(new_n867), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n891), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n882), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n895), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n897), .A2(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n283), .A2(new_n288), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n852), .A2(new_n853), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n857), .A2(new_n866), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n869), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n721), .B(KEYINPUT57), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n867), .A2(new_n188), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n765), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n893), .B1(new_n914), .B2(new_n916), .ZN(G54));
  NAND2_X1  g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT123), .Z(new_n919));
  AND3_X1   g733(.A1(new_n915), .A2(new_n358), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n358), .B1(new_n915), .B2(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n893), .ZN(G60));
  INV_X1    g736(.A(new_n893), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n859), .B2(new_n869), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n617), .A2(new_n619), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n927), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n925), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n911), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT124), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n911), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n928), .B1(new_n932), .B2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT60), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n909), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n604), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n909), .A2(new_n638), .A3(new_n937), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n923), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(KEYINPUT61), .A3(new_n923), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(G66));
  OAI21_X1  g759(.A(G953), .B1(new_n370), .B2(new_n423), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n832), .B2(G953), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n880), .B1(G898), .B2(new_n265), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G69));
  NAND2_X1  g763(.A1(new_n517), .A2(new_n519), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n353), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT125), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n828), .A2(new_n822), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n689), .A2(new_n674), .A3(new_n770), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n786), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n758), .B2(new_n772), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n666), .A2(new_n687), .A3(new_n719), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n683), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n952), .B1(new_n961), .B2(new_n265), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n770), .B(new_n769), .C1(new_n753), .C2(KEYINPUT44), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n757), .B2(new_n754), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n817), .A2(new_n846), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n965), .A2(new_n769), .B1(new_n689), .B2(new_n739), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n786), .A2(new_n957), .A3(new_n966), .A4(new_n737), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT126), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n786), .A2(new_n737), .A3(new_n966), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n773), .A2(new_n969), .A3(new_n970), .A4(new_n957), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n971), .A3(new_n265), .ZN(new_n972));
  INV_X1    g786(.A(new_n951), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(G900), .B2(G953), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n962), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n265), .B1(G227), .B2(G900), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n972), .A2(new_n974), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n976), .B1(new_n979), .B2(new_n962), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G72));
  NAND2_X1  g795(.A1(new_n521), .A2(new_n499), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n956), .A2(new_n959), .A3(new_n832), .A4(new_n960), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n988), .B(new_n982), .C1(new_n983), .C2(new_n985), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n521), .A2(new_n499), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n968), .A2(new_n832), .A3(new_n971), .ZN(new_n992));
  INV_X1    g806(.A(new_n985), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n854), .A2(new_n858), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n678), .B1(new_n521), .B2(new_n522), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n996), .A2(new_n993), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n893), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n990), .A2(new_n999), .ZN(G57));
endmodule


