//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n445, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G259));
  XOR2_X1   g021(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AND2_X1   g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n457), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n466), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OR2_X1    g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT69), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(G113), .A3(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(G2105), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT70), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2105), .C1(new_n476), .C2(new_n481), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n472), .B1(new_n483), .B2(new_n485), .ZN(G160));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(new_n466), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n493));
  INV_X1    g068(.A(G136), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n493), .C1(new_n494), .C2(new_n470), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n487), .B2(new_n488), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n501), .C1(new_n488), .C2(new_n487), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n505));
  OAI211_X1 g080(.A(G126), .B(G2105), .C1(new_n487), .C2(new_n488), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  AND3_X1   g083(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n503), .B2(new_n507), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(G164));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(G50), .A3(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT72), .A3(G543), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(new_n520), .B1(KEYINPUT5), .B2(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n514), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n515), .B1(new_n522), .B2(new_n523), .C1(new_n524), .C2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  AND2_X1   g102(.A1(new_n514), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n514), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n530), .B(KEYINPUT73), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n521), .A2(G89), .A3(new_n514), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n533), .A2(new_n534), .A3(new_n537), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n537), .A2(new_n541), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT73), .B1(new_n529), .B2(new_n530), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT74), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G168));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT75), .B(G52), .Z(new_n548));
  OAI22_X1  g123(.A1(new_n522), .A2(new_n547), .B1(new_n535), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT76), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n521), .A2(G64), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n525), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  AOI22_X1  g129(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n525), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n522), .A2(new_n557), .B1(new_n535), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  AOI22_X1  g140(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n525), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n521), .A2(new_n514), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G91), .ZN(new_n569));
  OAI211_X1 g144(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n570));
  NAND2_X1  g145(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n570), .B(new_n571), .Z(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n569), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  AND2_X1   g149(.A1(new_n542), .A2(new_n545), .ZN(G286));
  NAND2_X1  g150(.A1(new_n568), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n528), .A2(G49), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  AOI22_X1  g154(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n525), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n521), .A2(G86), .A3(new_n514), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  XNOR2_X1  g161(.A(KEYINPUT79), .B(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n568), .A2(G85), .B1(new_n528), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(KEYINPUT78), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(new_n521), .A2(G66), .ZN(new_n597));
  INV_X1    g172(.A(G79), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n517), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n521), .A2(G92), .A3(new_n514), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G321));
  XNOR2_X1  g183(.A(G299), .B(KEYINPUT81), .ZN(new_n609));
  MUX2_X1   g184(.A(G286), .B(new_n609), .S(new_n605), .Z(G297));
  MUX2_X1   g185(.A(G286), .B(new_n609), .S(new_n605), .Z(G280));
  INV_X1    g186(.A(new_n604), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g192(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n618));
  XNOR2_X1  g193(.A(G323), .B(new_n618), .ZN(G282));
  NAND2_X1  g194(.A1(new_n469), .A2(new_n467), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  INV_X1    g200(.A(new_n470), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n490), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n466), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n624), .A2(new_n625), .A3(new_n633), .ZN(G156));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G401));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n623), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n632), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  MUX2_X1   g249(.A(new_n674), .B(new_n673), .S(new_n666), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n585), .B2(G16), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT32), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1971), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n691), .A2(G23), .ZN(new_n697));
  INV_X1    g272(.A(G288), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n698), .B2(new_n691), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT33), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT86), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n694), .B2(new_n695), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n690), .A2(new_n696), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n691), .A2(G24), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT84), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n691), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT85), .B(G1986), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n626), .A2(G131), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n490), .A2(G119), .ZN(new_n716));
  OR2_X1    g291(.A1(G95), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(new_n713), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  NOR3_X1   g298(.A1(new_n711), .A2(new_n712), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n690), .A2(new_n725), .A3(new_n696), .A4(new_n703), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n705), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n691), .A2(G19), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT90), .Z(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n560), .B2(new_n691), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1341), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n713), .A2(G26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n626), .A2(G140), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n490), .A2(G128), .ZN(new_n738));
  OR2_X1    g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(new_n713), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n691), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n612), .B2(new_n691), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT89), .ZN(new_n747));
  INV_X1    g322(.A(G1348), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n734), .B(new_n744), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n730), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n691), .A2(G20), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT23), .ZN(new_n753));
  INV_X1    g328(.A(G299), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n691), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n713), .A2(G33), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT25), .ZN(new_n759));
  NAND2_X1  g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  INV_X1    g335(.A(G127), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n489), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(G2105), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n759), .B(new_n763), .C1(G139), .C2(new_n626), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(new_n713), .ZN(new_n765));
  NAND2_X1  g340(.A1(G162), .A2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G29), .B2(G35), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT29), .B(G2090), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n765), .A2(G2072), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G2072), .B2(new_n765), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n767), .A2(new_n769), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT31), .B(G11), .Z(new_n773));
  NOR2_X1   g348(.A1(new_n631), .A2(new_n713), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT30), .B(G28), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n773), .B(new_n774), .C1(new_n713), .C2(new_n775), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n713), .A2(G32), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n626), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n490), .A2(G129), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT26), .Z(new_n781));
  NAND3_X1  g356(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n777), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n772), .A2(new_n776), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n713), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n713), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2078), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n756), .A2(new_n771), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G34), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n713), .B1(new_n792), .B2(G34), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G160), .B2(G29), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(G2084), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT96), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(G2084), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT93), .Z(new_n802));
  NOR2_X1   g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n691), .A2(G5), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G171), .B2(new_n691), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT95), .B(G1961), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n791), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G21), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G168), .B2(G16), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT94), .B(G1966), .Z(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n751), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n728), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n705), .A2(new_n724), .A3(new_n815), .A4(new_n726), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n749), .A2(new_n730), .A3(new_n750), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n729), .A2(new_n814), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(G311));
  XNOR2_X1  g395(.A(new_n818), .B(KEYINPUT98), .ZN(G150));
  AOI22_X1  g396(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(new_n525), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n568), .A2(G93), .B1(new_n528), .B2(G55), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(new_n826), .C1(new_n556), .C2(new_n559), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT99), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n822), .A2(new_n525), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n522), .A2(new_n830), .B1(new_n535), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n826), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n560), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n827), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n612), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n840));
  AOI21_X1  g415(.A(G860), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT101), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n825), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XOR2_X1   g421(.A(KEYINPUT104), .B(G37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n505), .A2(new_n506), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n500), .B2(new_n502), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n741), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n782), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n764), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n719), .B(new_n621), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n626), .A2(G142), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT103), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n490), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n466), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n853), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n631), .B(KEYINPUT102), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G160), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n852), .A2(new_n860), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n852), .B(new_n868), .ZN(new_n869));
  OAI221_X1 g444(.A(new_n847), .B1(new_n865), .B2(new_n866), .C1(new_n869), .C2(new_n864), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g446(.A1(new_n698), .A2(KEYINPUT107), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  NAND2_X1  g448(.A1(G288), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n872), .A2(G305), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G305), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(G290), .A2(G166), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n594), .A2(G303), .A3(new_n595), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT108), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT42), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n835), .B(new_n615), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n604), .A2(G299), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n572), .A2(new_n569), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n887), .A2(new_n567), .A3(new_n600), .A4(new_n603), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT106), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(KEYINPUT41), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n895), .B2(new_n885), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT109), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n884), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n896), .B(KEYINPUT109), .Z(new_n899));
  NOR2_X1   g474(.A1(new_n884), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(G868), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n825), .A2(new_n605), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(G295));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(G331));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n892), .A2(KEYINPUT110), .ZN(new_n907));
  NAND2_X1  g482(.A1(G286), .A2(new_n835), .ZN(new_n908));
  NAND3_X1  g483(.A1(G168), .A2(new_n827), .A3(new_n834), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(G171), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G171), .B1(new_n908), .B2(new_n909), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n906), .B(new_n907), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n908), .A2(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G301), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n890), .A3(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n882), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n895), .B1(new_n911), .B2(new_n912), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n915), .A2(new_n886), .A3(new_n888), .A4(new_n910), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n878), .A2(new_n879), .ZN(new_n920));
  INV_X1    g495(.A(new_n877), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n919), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n925), .A3(new_n847), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT112), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n917), .A2(new_n925), .A3(new_n928), .A4(new_n847), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(KEYINPUT43), .A3(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n911), .A2(new_n912), .A3(new_n889), .ZN(new_n931));
  INV_X1    g506(.A(new_n895), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n915), .B2(new_n910), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n882), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n925), .A4(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n937), .A2(KEYINPUT44), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n930), .A2(new_n938), .A3(KEYINPUT113), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT113), .B1(new_n930), .B2(new_n938), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n934), .A2(new_n936), .A3(new_n925), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n917), .A2(new_n925), .A3(new_n935), .A4(new_n847), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI211_X1 g522(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  OAI22_X1  g523(.A1(new_n939), .A2(new_n940), .B1(new_n947), .B2(new_n948), .ZN(G397));
  INV_X1    g524(.A(KEYINPUT125), .ZN(new_n950));
  NAND2_X1  g525(.A1(G286), .A2(G8), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n952));
  INV_X1    g527(.A(new_n502), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n501), .B1(new_n469), .B2(new_n498), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT71), .B1(new_n955), .B2(new_n848), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n957));
  AOI211_X1 g532(.A(new_n952), .B(G1384), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n952), .B1(new_n849), .B2(G1384), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(G40), .A3(G160), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n811), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  OAI211_X1 g537(.A(KEYINPUT50), .B(new_n962), .C1(new_n509), .C2(new_n510), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n503), .B2(new_n507), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G2084), .ZN(new_n969));
  NAND3_X1  g544(.A1(G160), .A2(G40), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n961), .A2(new_n972), .A3(KEYINPUT119), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT119), .ZN(new_n974));
  INV_X1    g549(.A(new_n472), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n478), .B(new_n480), .C1(new_n489), .C2(new_n473), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n484), .B1(new_n976), .B2(G2105), .ZN(new_n977));
  INV_X1    g552(.A(new_n485), .ZN(new_n978));
  OAI211_X1 g553(.A(G40), .B(new_n975), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n506), .B(new_n505), .C1(new_n953), .C2(new_n954), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT45), .B1(new_n980), .B2(new_n962), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT45), .B(new_n962), .C1(new_n509), .C2(new_n510), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n812), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n970), .B1(new_n963), .B2(new_n967), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n974), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n951), .B1(new_n973), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n973), .A2(new_n986), .A3(G168), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT120), .ZN(new_n989));
  OAI21_X1  g564(.A(G8), .B1(new_n989), .B2(KEYINPUT51), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n989), .B2(KEYINPUT51), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n993));
  OAI21_X1  g568(.A(G8), .B1(new_n984), .B2(new_n985), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n987), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT62), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n950), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n988), .A2(new_n991), .B1(new_n994), .B2(new_n993), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n999), .C2(new_n987), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT124), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n999), .A2(KEYINPUT62), .A3(new_n987), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n962), .B1(new_n509), .B2(new_n510), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n952), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n980), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(G160), .A3(G40), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1004), .B1(new_n1010), .B2(G2078), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n979), .B1(new_n963), .B2(new_n967), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(G1961), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1004), .A2(G2078), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n982), .A2(new_n983), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1016), .A2(G171), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  OAI21_X1  g593(.A(G1981), .B1(new_n581), .B2(new_n584), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n581), .A2(G1981), .A3(new_n584), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT116), .B(new_n1018), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1021), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(KEYINPUT116), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(G160), .A2(G40), .A3(new_n964), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n1026), .B2(G8), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1022), .B(new_n1025), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n698), .A2(G1976), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT115), .B(G1976), .Z(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1031), .B(new_n1033), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n979), .A2(new_n965), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1026), .A2(new_n1027), .A3(G8), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1037), .A2(new_n1038), .B1(new_n698), .B2(G1976), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1030), .B(new_n1034), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1971), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n966), .B(new_n962), .C1(new_n509), .C2(new_n510), .ZN(new_n1044));
  INV_X1    g619(.A(new_n979), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n524), .A2(new_n525), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n515), .B1(new_n522), .B2(new_n523), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT55), .B(G8), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1971), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n956), .A2(new_n957), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT45), .B1(new_n1059), .B2(new_n962), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1060), .B2(new_n1008), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n968), .A2(new_n1047), .A3(new_n1045), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1036), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1056), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1017), .A2(new_n1042), .A3(new_n1057), .A4(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1002), .B1(new_n1003), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n996), .A2(new_n997), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1031), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT52), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1057), .A3(new_n1065), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1016), .A2(G171), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(KEYINPUT124), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1001), .A2(new_n1067), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT126), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1001), .A2(new_n1067), .A3(new_n1075), .A4(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1036), .B(new_n1056), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1030), .ZN(new_n1081));
  OR2_X1    g656(.A1(G288), .A2(G1976), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1023), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1080), .A2(new_n1042), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1061), .A2(new_n1048), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1064), .B1(new_n1086), .B2(G8), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1041), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(G8), .B(G168), .C1(new_n984), .C2(new_n985), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT63), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(KEYINPUT63), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1092), .A2(new_n1080), .A3(new_n1041), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1085), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT122), .B(G2078), .Z(new_n1096));
  AND4_X1   g671(.A1(KEYINPUT53), .A2(new_n975), .A3(G40), .A4(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(new_n959), .A3(new_n482), .A4(new_n1007), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1011), .A2(new_n1013), .A3(G301), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1095), .B1(new_n1073), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1072), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1011), .A2(new_n1013), .A3(new_n1098), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1011), .A2(new_n1013), .A3(G301), .A4(new_n1015), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(KEYINPUT123), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(KEYINPUT123), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT54), .B(new_n1103), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n996), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1101), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(G299), .B(KEYINPUT57), .Z(new_n1110));
  AOI21_X1  g685(.A(new_n1008), .B1(new_n952), .B2(new_n1005), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1110), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1110), .B1(new_n1117), .B2(new_n1113), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT61), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1110), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1118), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n968), .A2(new_n1045), .ZN(new_n1128));
  INV_X1    g703(.A(G2067), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1128), .A2(new_n748), .B1(new_n1129), .B2(new_n1035), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n604), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1012), .A2(G1348), .B1(G2067), .B2(new_n1026), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n612), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1134), .A2(KEYINPUT60), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT117), .B(G1996), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1111), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1026), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1138), .A2(KEYINPUT118), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT118), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT59), .B(new_n560), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n560), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1127), .A2(new_n1136), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1133), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1118), .B1(new_n1148), .B2(new_n1120), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1094), .B1(new_n1109), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1077), .A2(new_n1079), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n979), .A2(new_n959), .ZN(new_n1153));
  INV_X1    g728(.A(G1996), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n782), .B(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n741), .B(new_n1129), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n719), .B(new_n722), .Z(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(G1986), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n708), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G290), .A2(G1986), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1153), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1152), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1153), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1159), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1162), .A2(new_n1153), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1168), .B2(KEYINPUT48), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(KEYINPUT48), .B2(new_n1168), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT46), .ZN(new_n1172));
  INV_X1    g747(.A(new_n782), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1156), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1172), .B1(new_n1165), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT47), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n720), .A2(new_n722), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1157), .A2(new_n1177), .B1(G2067), .B2(new_n741), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1153), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1170), .A2(new_n1176), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1164), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g757(.A1(G401), .A2(new_n464), .A3(G227), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n682), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1186));
  XNOR2_X1  g760(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n1187), .A2(new_n870), .A3(new_n945), .ZN(G225));
  INV_X1    g762(.A(G225), .ZN(G308));
endmodule


