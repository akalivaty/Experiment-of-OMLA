//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1180, new_n1181, new_n1182;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT68), .B(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  OR2_X1    g034(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G2104), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n458), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n464), .A2(G136), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(new_n463), .B2(new_n475), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n459), .A2(KEYINPUT70), .A3(new_n462), .A4(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n466), .A2(G138), .A3(new_n475), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n459), .A2(G138), .A3(new_n462), .A4(new_n475), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n459), .A2(G126), .A3(new_n462), .A4(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n487), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(new_n490), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n496), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(KEYINPUT72), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n506), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XOR2_X1   g089(.A(new_n514), .B(KEYINPUT73), .Z(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n509), .A2(new_n508), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(G63), .A2(G651), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n506), .A2(new_n523), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT5), .B(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(new_n505), .A3(G89), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n532), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n529), .B1(new_n528), .B2(new_n534), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n534), .B1(new_n512), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT74), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n544), .A2(KEYINPUT75), .A3(new_n526), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n539), .A2(new_n545), .ZN(G168));
  INV_X1    g121(.A(new_n506), .ZN(new_n547));
  INV_X1    g122(.A(new_n512), .ZN(new_n548));
  AOI22_X1  g123(.A1(G52), .A2(new_n547), .B1(new_n548), .B2(G90), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G651), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n547), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n548), .A2(G81), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n555), .B(new_n556), .C1(new_n551), .C2(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT76), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND3_X1  g139(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(G91), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n527), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n551), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n566), .A2(new_n569), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT75), .B1(new_n544), .B2(new_n526), .ZN(new_n574));
  AOI211_X1 g149(.A(new_n538), .B(new_n525), .C1(new_n542), .C2(new_n543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n539), .A2(new_n545), .A3(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G286));
  AND2_X1   g154(.A1(new_n567), .A2(new_n568), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G87), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n527), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(G49), .A2(new_n547), .B1(new_n582), .B2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  INV_X1    g159(.A(G73), .ZN(new_n585));
  INV_X1    g160(.A(G543), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT79), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT79), .B1(new_n585), .B2(new_n586), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n517), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  INV_X1    g166(.A(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n567), .A2(new_n568), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n591), .B1(new_n592), .B2(new_n506), .C1(new_n593), .C2(new_n594), .ZN(G305));
  AND2_X1   g170(.A1(new_n527), .A2(G60), .ZN(new_n596));
  AND2_X1   g171(.A1(G72), .A2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT80), .ZN(new_n599));
  AOI22_X1  g174(.A1(G47), .A2(new_n547), .B1(new_n548), .B2(G85), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n598), .A2(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n593), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n605), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n567), .A2(G92), .A3(new_n568), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n517), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(G54), .A2(new_n547), .B1(new_n612), .B2(G651), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n607), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n604), .B1(new_n615), .B2(G868), .ZN(G321));
  NOR2_X1   g192(.A1(G299), .A2(G868), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n578), .B2(G868), .ZN(G297));
  XOR2_X1   g194(.A(G297), .B(KEYINPUT82), .Z(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n615), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n625), .B(new_n626), .C1(G868), .C2(new_n559), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n464), .A2(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n475), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n483), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT85), .B(G2096), .Z(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n471), .A2(new_n466), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT13), .B(G2100), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n636), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n661), .B2(new_n658), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n663), .B2(new_n665), .ZN(new_n667));
  INV_X1    g242(.A(new_n658), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n664), .A3(new_n660), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n659), .A2(new_n664), .A3(new_n661), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n679), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT20), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n676), .A2(new_n680), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT87), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(KEYINPUT87), .ZN(new_n686));
  AOI211_X1 g261(.A(new_n681), .B(new_n683), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  XOR2_X1   g271(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT90), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(G288), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n706), .B(new_n707), .Z(new_n708));
  MUX2_X1   g283(.A(G6), .B(G305), .S(G16), .Z(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n702), .A2(KEYINPUT90), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n703), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n715));
  INV_X1    g290(.A(new_n483), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G119), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT89), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G131), .B2(new_n464), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G25), .B2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  AND2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n698), .A2(G24), .ZN(new_n729));
  INV_X1    g304(.A(G290), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n698), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1986), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n727), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n714), .B2(KEYINPUT34), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n697), .B1(new_n715), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n736));
  INV_X1    g311(.A(new_n697), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n733), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n740), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT29), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G2090), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT96), .Z(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n748));
  OR2_X1    g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  NAND2_X1  g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G5), .A2(G16), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT95), .Z(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G301), .B2(new_n698), .ZN(new_n754));
  INV_X1    g329(.A(G1961), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n755), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n698), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n559), .B2(new_n698), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n633), .A2(new_n740), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n464), .A2(G139), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n475), .C2(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G33), .B(new_n766), .S(G29), .Z(new_n767));
  AOI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(G2072), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n698), .A2(G4), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n615), .B2(new_n698), .ZN(new_n770));
  INV_X1    g345(.A(G1348), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AND4_X1   g347(.A1(new_n757), .A2(new_n760), .A3(new_n768), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n767), .A2(G2072), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT93), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n740), .B1(KEYINPUT24), .B2(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(KEYINPUT24), .B2(G34), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n473), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n698), .A2(G20), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G299), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n775), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n740), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n740), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G2078), .Z(new_n790));
  NAND3_X1  g365(.A1(new_n773), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n740), .A2(G32), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n464), .A2(G141), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT94), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n716), .A2(G129), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT26), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n471), .A2(G105), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n794), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G168), .A2(new_n698), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n698), .B2(G21), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n804), .B1(G1966), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n809), .A2(new_n806), .B1(new_n802), .B2(new_n803), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n740), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT28), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n716), .A2(G128), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n475), .A2(G116), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n464), .A2(G140), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT92), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n808), .B(new_n810), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n743), .A2(G2090), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT97), .ZN(new_n826));
  NOR4_X1   g401(.A1(new_n745), .A2(new_n791), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n735), .A2(new_n739), .A3(new_n827), .ZN(G150));
  XNOR2_X1  g403(.A(G150), .B(KEYINPUT99), .ZN(G311));
  NAND2_X1  g404(.A1(new_n615), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n547), .A2(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n548), .A2(G93), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OAI211_X1 g409(.A(new_n832), .B(new_n833), .C1(new_n551), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n559), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n558), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n831), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n842), .ZN(new_n845));
  INV_X1    g420(.A(new_n838), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n633), .B(new_n473), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G162), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n766), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n801), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n500), .A2(new_n501), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(new_n855), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n818), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  INV_X1    g435(.A(new_n818), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n861), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n464), .A2(G142), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n475), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n716), .B2(G130), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT102), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n722), .B(new_n639), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n859), .A2(new_n862), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n859), .B2(new_n862), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n872), .B1(new_n873), .B2(KEYINPUT103), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n859), .A2(new_n862), .A3(new_n871), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n851), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n873), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n851), .A3(new_n872), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT40), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n884), .A2(new_n877), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n886), .ZN(G395));
  INV_X1    g462(.A(G868), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n846), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(G290), .B(G305), .Z(new_n890));
  XNOR2_X1  g465(.A(G303), .B(new_n705), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n893));
  NOR2_X1   g468(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n840), .B(new_n623), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  INV_X1    g472(.A(G299), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n614), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g474(.A1(G299), .A2(new_n607), .A3(new_n609), .A4(new_n613), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n897), .B1(new_n614), .B2(new_n898), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT41), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  INV_X1    g481(.A(new_n902), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n900), .A4(new_n899), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n905), .B1(new_n896), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n895), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n889), .B1(new_n912), .B2(new_n888), .ZN(G295));
  OAI21_X1  g488(.A(new_n889), .B1(new_n912), .B2(new_n888), .ZN(G331));
  NAND3_X1  g489(.A1(new_n576), .A2(G171), .A3(new_n577), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(G168), .B2(G301), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n576), .A2(new_n916), .A3(G171), .A4(new_n577), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n918), .A2(new_n840), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n840), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n920), .A2(new_n921), .A3(new_n903), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n919), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n841), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n840), .A3(new_n919), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n910), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT107), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n892), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n906), .A2(new_n909), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n920), .B2(new_n921), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n904), .A3(new_n925), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n927), .A2(new_n928), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n931), .A3(new_n892), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n935), .A2(new_n881), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT108), .B1(new_n937), .B2(KEYINPUT43), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n931), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n929), .B(new_n939), .C1(new_n920), .C2(new_n921), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n928), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n936), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n935), .A2(new_n881), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n930), .A2(new_n931), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n892), .B1(new_n947), .B2(KEYINPUT107), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n948), .B2(new_n933), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n949), .B2(new_n944), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n938), .B1(new_n950), .B2(KEYINPUT108), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n943), .A2(new_n936), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n934), .A2(new_n936), .A3(new_n944), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n920), .A2(new_n921), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n930), .A2(KEYINPUT109), .B1(new_n958), .B2(new_n904), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n892), .B1(new_n959), .B2(new_n941), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n960), .B2(new_n946), .ZN(new_n961));
  AND4_X1   g536(.A1(new_n952), .A2(new_n961), .A3(KEYINPUT44), .A4(new_n956), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n951), .A2(KEYINPUT44), .B1(new_n957), .B2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n492), .B2(new_n496), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n465), .A2(G40), .A3(new_n470), .A4(new_n472), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n818), .B(new_n821), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n801), .A2(G1996), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT112), .ZN(new_n976));
  INV_X1    g551(.A(new_n801), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT113), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n722), .B(new_n726), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n970), .B2(new_n980), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n970), .A2(G1986), .A3(G290), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT111), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n965), .A2(new_n968), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1976), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(G288), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT52), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n990), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n506), .A2(new_n592), .B1(new_n512), .B2(new_n594), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g574(.A(KEYINPUT116), .B1(new_n512), .B2(new_n594), .C1(new_n592), .C2(new_n506), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(new_n591), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G1981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT117), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1004), .A3(G1981), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n996), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n989), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1008), .A2(new_n989), .A3(KEYINPUT118), .A4(new_n1009), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n995), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT72), .B1(new_n500), .B2(new_n501), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n492), .A2(new_n487), .A3(new_n496), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n964), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT50), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  INV_X1    g599(.A(new_n968), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n964), .C1(new_n492), .C2(new_n496), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT114), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n855), .A2(new_n1029), .A3(new_n1026), .A4(new_n964), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n966), .A2(G1384), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n968), .B1(new_n855), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n701), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n988), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1014), .A2(new_n1019), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n996), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G288), .A2(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n989), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT63), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n967), .A2(new_n1025), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1033), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n497), .B2(new_n502), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n809), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1023), .A2(new_n779), .A3(new_n1025), .A4(new_n1031), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT120), .B(new_n809), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(G8), .A3(new_n578), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n968), .B1(KEYINPUT50), .B2(new_n965), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1024), .B(new_n1059), .C1(new_n1022), .C2(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n988), .B1(new_n1037), .B2(new_n1060), .ZN(new_n1061));
  OR3_X1    g636(.A1(new_n1061), .A2(KEYINPUT119), .A3(new_n1019), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1038), .A2(new_n1019), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT119), .B1(new_n1061), .B2(new_n1019), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1014), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1046), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1056), .B(KEYINPUT121), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1038), .A2(new_n1019), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n1046), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1067), .A2(new_n1063), .A3(new_n1014), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1045), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1055), .A2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G168), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1055), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1052), .A2(new_n1053), .A3(G168), .A4(new_n1054), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(G8), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT125), .B1(new_n1055), .B2(G8), .ZN(new_n1081));
  OAI211_X1 g656(.A(G8), .B(new_n1078), .C1(new_n1081), .C2(new_n1072), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(new_n1085), .A3(new_n1082), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1025), .B1(new_n1035), .B2(new_n1026), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT123), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1023), .A2(new_n1090), .A3(new_n1025), .A4(new_n1031), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n755), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G2078), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OR3_X1    g670(.A1(new_n1047), .A2(new_n1049), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1093), .B1(new_n1036), .B2(G2078), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G171), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1065), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1084), .A2(new_n1086), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1071), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1089), .A2(new_n771), .A3(new_n1091), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n987), .A2(new_n821), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(KEYINPUT60), .A3(new_n1104), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n615), .A3(new_n1108), .ZN(new_n1109));
  AOI211_X1 g684(.A(KEYINPUT50), .B(G1384), .C1(new_n497), .C2(new_n502), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1059), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n785), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(G299), .B(KEYINPUT57), .Z(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1034), .B(new_n1114), .C1(new_n1035), .C2(KEYINPUT45), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT122), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1112), .A2(new_n1119), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1034), .B(new_n974), .C1(new_n1035), .C2(KEYINPUT45), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n965), .B2(new_n968), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1125), .A2(KEYINPUT59), .A3(new_n559), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT59), .B1(new_n1125), .B2(new_n559), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1113), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1121), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1108), .A2(new_n615), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1105), .A2(new_n615), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT124), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1105), .A2(new_n1138), .A3(new_n615), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1139), .A3(new_n1131), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1109), .A2(new_n1135), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n469), .A2(KEYINPUT127), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n475), .B1(new_n469), .B2(KEYINPUT127), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(G40), .A3(new_n1094), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n465), .A2(new_n472), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(KEYINPUT126), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n855), .A2(new_n1033), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n967), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1092), .A2(new_n1097), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1099), .B1(G171), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1065), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1152), .A2(G171), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(KEYINPUT54), .C1(G171), .C2(new_n1098), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1155), .A2(new_n1156), .A3(new_n1083), .A4(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1142), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n986), .B1(new_n1102), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n976), .B(KEYINPUT46), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n971), .A2(new_n977), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n969), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT47), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n982), .B(KEYINPUT48), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n981), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n979), .A2(new_n723), .A3(new_n726), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n861), .A2(new_n821), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n970), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1161), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g748(.A(G319), .ZN(new_n1175));
  NOR3_X1   g749(.A1(G401), .A2(G227), .A3(new_n1175), .ZN(new_n1176));
  AND3_X1   g750(.A1(new_n694), .A2(new_n695), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n1177), .B1(new_n884), .B2(new_n877), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n1178), .ZN(G308));
  INV_X1    g753(.A(KEYINPUT108), .ZN(new_n1180));
  NAND2_X1  g754(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1181), .B2(new_n945), .ZN(new_n1182));
  OAI221_X1 g756(.A(new_n1177), .B1(new_n877), .B2(new_n884), .C1(new_n1182), .C2(new_n938), .ZN(G225));
endmodule


