//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  INV_X1    g000(.A(KEYINPUT2), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n189), .A2(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n196), .B2(new_n192), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G143), .B(G146), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT0), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT0), .B(G128), .Z(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n205), .A2(new_n206), .A3(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G134), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n207), .B1(new_n212), .B2(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(G134), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G137), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n215), .A3(new_n218), .A4(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT65), .B(G131), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n213), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n213), .B2(new_n220), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n204), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n213), .A2(new_n220), .A3(new_n221), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n212), .B1(G134), .B2(new_n208), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G131), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G143), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(new_n232), .C1(KEYINPUT1), .C2(new_n201), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n232), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(G128), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n226), .A2(new_n228), .A3(new_n233), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n198), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n225), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(KEYINPUT69), .B(new_n204), .C1(new_n222), .C2(new_n224), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n236), .A2(new_n233), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT70), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n246), .A3(new_n233), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n226), .A2(new_n228), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n242), .A2(KEYINPUT30), .A3(new_n243), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n240), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT31), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n254), .B(KEYINPUT27), .Z(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n255), .B(new_n256), .Z(new_n257));
  NAND4_X1  g071(.A1(new_n242), .A2(new_n198), .A3(new_n243), .A4(new_n248), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n250), .A2(new_n251), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n257), .A3(new_n258), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT31), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n257), .ZN(new_n264));
  INV_X1    g078(.A(new_n224), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n226), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n197), .B1(new_n266), .B2(new_n204), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT28), .B1(new_n267), .B2(new_n248), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n238), .A2(new_n197), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n258), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI211_X1 g088(.A(KEYINPUT72), .B(new_n270), .C1(new_n258), .C2(new_n271), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n264), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n261), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n263), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(G472), .A2(G902), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(KEYINPUT73), .A3(new_n279), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n242), .A2(new_n243), .A3(new_n248), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n197), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n258), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n269), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT76), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n274), .A2(new_n264), .A3(new_n275), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n250), .A2(new_n258), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(new_n257), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n297), .A2(KEYINPUT29), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G472), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n282), .A2(KEYINPUT75), .A3(new_n283), .A4(new_n284), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n278), .A2(KEYINPUT32), .A3(new_n279), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n287), .A2(new_n301), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G234), .ZN(new_n305));
  OAI21_X1  g119(.A(G217), .B1(new_n305), .B2(G902), .ZN(new_n306));
  XNOR2_X1  g120(.A(G125), .B(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT16), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n309), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n229), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(G146), .A3(new_n310), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(G128), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n317), .B(new_n318), .C1(G119), .C2(new_n201), .ZN(new_n319));
  XNOR2_X1  g133(.A(G119), .B(G128), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT24), .B(G110), .Z(new_n321));
  AOI22_X1  g135(.A1(new_n319), .A2(G110), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n319), .A2(G110), .B1(new_n320), .B2(new_n321), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n307), .A2(new_n229), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n313), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT22), .B(G137), .ZN(new_n328));
  INV_X1    g142(.A(G221), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n329), .A2(new_n305), .A3(G953), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT77), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n323), .A2(new_n326), .A3(new_n331), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G902), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n306), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n337), .B2(new_n336), .ZN(new_n339));
  AOI21_X1  g153(.A(G902), .B1(new_n305), .B2(G217), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n333), .B2(new_n334), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n304), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G214), .B1(G237), .B2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G107), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT79), .A3(G104), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(new_n347), .A3(KEYINPUT79), .A4(G104), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G101), .ZN(new_n354));
  INV_X1    g168(.A(G101), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n347), .A2(KEYINPUT79), .A3(G104), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n357), .B2(G107), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n355), .B(new_n352), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n354), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n353), .A2(new_n361), .A3(G101), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n197), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n357), .A2(G107), .ZN(new_n366));
  OAI21_X1  g180(.A(G101), .B1(new_n366), .B2(new_n349), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n316), .A3(G116), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G113), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n196), .B2(KEYINPUT5), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n373), .A2(KEYINPUT86), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(KEYINPUT86), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n194), .B(new_n369), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G122), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n365), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n204), .A2(new_n309), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n244), .A2(new_n309), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n253), .A2(G224), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n379), .A2(new_n380), .B1(KEYINPUT7), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n204), .A2(new_n383), .A3(new_n309), .ZN(new_n385));
  AND4_X1   g199(.A1(new_n381), .A2(new_n384), .A3(new_n385), .A4(new_n380), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n386), .B2(KEYINPUT7), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n378), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n374), .A2(new_n375), .ZN(new_n389));
  INV_X1    g203(.A(new_n194), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n368), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n194), .B1(new_n372), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n368), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n377), .B(KEYINPUT8), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(G902), .B1(new_n388), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n377), .B1(new_n365), .B2(new_n376), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n384), .A2(new_n385), .A3(new_n380), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n401), .B(new_n381), .Z(new_n402));
  NAND2_X1  g216(.A1(new_n378), .A2(KEYINPUT6), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n400), .B(new_n402), .C1(new_n403), .C2(new_n398), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G210), .B1(G237), .B2(G902), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n397), .A2(new_n404), .A3(new_n406), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n346), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  AOI211_X1 g225(.A(G953), .B(new_n411), .C1(G234), .C2(G237), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT21), .B(G898), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT94), .ZN(new_n415));
  AOI211_X1 g229(.A(new_n288), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n413), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  XOR2_X1   g234(.A(G110), .B(G140), .Z(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT78), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n253), .A2(G227), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n422), .B(new_n423), .Z(new_n424));
  NAND4_X1  g238(.A1(new_n359), .A2(new_n236), .A3(new_n233), .A4(new_n367), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT10), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n362), .A2(new_n204), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n355), .B1(new_n350), .B2(new_n352), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT80), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n360), .A2(new_n433), .A3(new_n204), .A4(new_n362), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n427), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n359), .A2(KEYINPUT10), .A3(new_n367), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n245), .A2(new_n436), .A3(new_n247), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT81), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n245), .A2(new_n436), .A3(new_n439), .A4(new_n247), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n435), .A2(new_n441), .A3(KEYINPUT84), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT84), .B1(new_n435), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n266), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n265), .A2(KEYINPUT82), .A3(new_n226), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n222), .B2(new_n224), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n435), .A2(new_n448), .A3(new_n441), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n424), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n424), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n368), .A2(new_n244), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n425), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n266), .B(new_n453), .C1(KEYINPUT83), .C2(KEYINPUT12), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n453), .B1(new_n222), .B2(new_n224), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT83), .B1(new_n222), .B2(new_n224), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n451), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n420), .B(new_n288), .C1(new_n450), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n454), .A2(new_n458), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n449), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n424), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n266), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n435), .A2(new_n441), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n435), .A2(new_n441), .A3(KEYINPUT84), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n464), .B(G469), .C1(new_n470), .C2(new_n451), .ZN(new_n471));
  NAND2_X1  g285(.A1(G469), .A2(G902), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n460), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT9), .B(G234), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n329), .B1(new_n475), .B2(new_n288), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n314), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n252), .A2(new_n253), .A3(G214), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(new_n231), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n480), .B1(new_n483), .B2(new_n221), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n485));
  INV_X1    g299(.A(new_n221), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(KEYINPUT88), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n221), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n484), .A2(new_n485), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n484), .A2(new_n487), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n479), .B(new_n489), .C1(new_n490), .C2(new_n485), .ZN(new_n491));
  XNOR2_X1  g305(.A(G113), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n357), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT18), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n483), .B1(new_n494), .B2(new_n223), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n482), .A2(KEYINPUT18), .A3(G131), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n307), .B(new_n229), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n493), .B1(new_n491), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n288), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G475), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n307), .A2(KEYINPUT89), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n505), .B(KEYINPUT19), .Z(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n229), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n507), .A3(new_n313), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(new_n498), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n499), .B1(new_n509), .B2(new_n493), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT20), .ZN(new_n511));
  NOR2_X1   g325(.A1(G475), .A2(G902), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT90), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n511), .B1(new_n510), .B2(new_n513), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n503), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G122), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G116), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT91), .Z(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(G116), .B2(new_n517), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(G107), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n231), .A2(G128), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n201), .A2(G143), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT92), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n210), .A2(new_n211), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(KEYINPUT13), .ZN(new_n530));
  MUX2_X1   g344(.A(KEYINPUT13), .B(new_n530), .S(new_n522), .Z(new_n531));
  AOI22_X1  g345(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(G134), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n521), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n347), .B1(new_n519), .B2(KEYINPUT14), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n534), .A2(new_n520), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(new_n529), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n526), .B(new_n527), .C1(new_n210), .C2(new_n211), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT93), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n520), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n535), .A2(new_n539), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n533), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G217), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n474), .A2(new_n545), .A3(G953), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n533), .A2(new_n543), .A3(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n288), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(G478), .ZN(new_n553));
  INV_X1    g367(.A(G478), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n550), .B(new_n288), .C1(KEYINPUT15), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR4_X1   g370(.A1(new_n419), .A2(new_n478), .A3(new_n516), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n344), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G101), .ZN(G3));
  AND2_X1   g373(.A1(new_n282), .A2(new_n283), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n278), .A2(new_n288), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G472), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n478), .A2(new_n342), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n550), .B(KEYINPUT33), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n554), .B1(new_n566), .B2(new_n288), .ZN(new_n567));
  INV_X1    g381(.A(new_n551), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n567), .B1(new_n554), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n516), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(new_n419), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT95), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT34), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G104), .ZN(G6));
  INV_X1    g389(.A(new_n516), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n556), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n419), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n564), .A2(new_n565), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G107), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(G9));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n332), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(new_n327), .Z(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n340), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n339), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n564), .A2(new_n557), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT37), .B(G110), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G12));
  INV_X1    g403(.A(new_n478), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n413), .B1(new_n417), .B2(G900), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n577), .A2(new_n592), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n593), .A2(new_n410), .A3(new_n586), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n304), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n304), .A2(KEYINPUT96), .A3(new_n590), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G128), .ZN(G30));
  XNOR2_X1  g414(.A(new_n591), .B(KEYINPUT39), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n590), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT40), .Z(new_n603));
  NAND2_X1  g417(.A1(new_n408), .A2(new_n409), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(KEYINPUT38), .Z(new_n605));
  NAND2_X1  g419(.A1(new_n516), .A2(new_n556), .ZN(new_n606));
  NOR4_X1   g420(.A1(new_n605), .A2(new_n346), .A3(new_n586), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n291), .A2(new_n264), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT97), .A3(new_n261), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n288), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT97), .B1(new_n608), .B2(new_n261), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n287), .A2(new_n302), .A3(new_n303), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n603), .A2(new_n607), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT98), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n231), .ZN(G45));
  INV_X1    g430(.A(new_n570), .ZN(new_n617));
  AND4_X1   g431(.A1(new_n410), .A2(new_n617), .A3(new_n586), .A4(new_n591), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n304), .A2(new_n618), .A3(new_n590), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G146), .ZN(G48));
  INV_X1    g434(.A(new_n450), .ZN(new_n621));
  INV_X1    g435(.A(new_n459), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n420), .B1(new_n623), .B2(new_n288), .ZN(new_n624));
  INV_X1    g438(.A(new_n460), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n477), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(KEYINPUT99), .A3(new_n477), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(new_n304), .A3(new_n343), .A4(new_n571), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT41), .B(G113), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G15));
  NAND4_X1  g448(.A1(new_n631), .A2(new_n304), .A3(new_n343), .A4(new_n578), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G116), .ZN(G18));
  NAND2_X1  g450(.A1(new_n623), .A2(new_n288), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G469), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n410), .A2(new_n638), .A3(new_n477), .A4(new_n460), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n626), .A2(KEYINPUT100), .A3(new_n477), .A4(new_n410), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n516), .A2(new_n556), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n418), .A3(new_n586), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n304), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G119), .ZN(G21));
  NAND2_X1  g463(.A1(new_n562), .A2(KEYINPUT101), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n293), .A2(new_n264), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n262), .A3(new_n259), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n279), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n562), .A2(KEYINPUT101), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n343), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n606), .B(KEYINPUT102), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n410), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(new_n629), .A3(new_n418), .A4(new_n630), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n517), .ZN(G24));
  INV_X1    g476(.A(new_n586), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n654), .A2(new_n663), .A3(new_n655), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n570), .A2(new_n592), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n665), .A3(new_n643), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G125), .ZN(G27));
  NOR2_X1   g481(.A1(new_n604), .A2(new_n346), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n471), .A2(KEYINPUT103), .ZN(new_n670));
  INV_X1    g484(.A(new_n451), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n444), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n672), .A2(new_n673), .A3(G469), .A4(new_n464), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n460), .A2(new_n472), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT104), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n670), .A2(new_n674), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n460), .A4(new_n472), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n477), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT105), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n681), .A2(new_n684), .A3(new_n477), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n669), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n570), .A2(KEYINPUT42), .A3(new_n592), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n344), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n684), .B1(new_n681), .B2(new_n477), .ZN(new_n689));
  AOI211_X1 g503(.A(KEYINPUT105), .B(new_n476), .C1(new_n677), .C2(new_n680), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n665), .B(new_n668), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  INV_X1    g506(.A(new_n303), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT32), .B1(new_n278), .B2(new_n279), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT32), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n280), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(KEYINPUT106), .A3(new_n303), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(new_n301), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n343), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT107), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n699), .A2(new_n702), .A3(new_n343), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n691), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n688), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n223), .ZN(G33));
  NAND4_X1  g521(.A1(new_n686), .A2(new_n304), .A3(new_n343), .A4(new_n593), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  XNOR2_X1  g523(.A(new_n516), .B(KEYINPUT109), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n569), .A3(KEYINPUT43), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n569), .A2(new_n576), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n713), .B(new_n714), .C1(KEYINPUT43), .C2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n563), .A3(new_n586), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n464), .B1(new_n470), .B2(new_n451), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n472), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n625), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT108), .B1(new_n723), .B2(new_n724), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n477), .A3(new_n601), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n717), .A2(new_n718), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n719), .A2(new_n668), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G137), .ZN(G39));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n477), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT47), .Z(new_n735));
  NAND3_X1  g549(.A1(new_n665), .A2(new_n342), .A3(new_n668), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n304), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G140), .ZN(G42));
  NAND2_X1  g553(.A1(new_n619), .A2(new_n666), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n658), .A2(new_n410), .A3(new_n663), .A4(new_n591), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n682), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n613), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT113), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n613), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n599), .A2(new_n741), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n740), .B1(new_n597), .B2(new_n598), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT114), .A3(new_n748), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(KEYINPUT52), .A3(new_n748), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n645), .A2(new_n591), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n645), .A2(new_n760), .A3(new_n591), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n668), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n586), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n304), .A3(new_n590), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n686), .A2(new_n665), .A3(new_n664), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n708), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n706), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n572), .A2(new_n579), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n558), .A2(new_n770), .A3(new_n587), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n661), .B1(new_n647), .B2(new_n304), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT116), .A3(new_n632), .A4(new_n635), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n657), .A2(new_n660), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n648), .A2(new_n776), .A3(new_n632), .A4(new_n635), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n769), .A2(new_n773), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n757), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n777), .A2(new_n771), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n769), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n752), .B2(new_n748), .ZN(new_n786));
  AND4_X1   g600(.A1(KEYINPUT114), .A2(new_n599), .A3(new_n748), .A4(new_n741), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n785), .B1(new_n788), .B2(new_n755), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n782), .B(new_n783), .C1(new_n789), .C2(KEYINPUT53), .ZN(new_n790));
  INV_X1    g604(.A(new_n785), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n757), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n751), .A2(new_n754), .A3(new_n753), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n754), .B1(new_n751), .B2(new_n753), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT115), .B1(new_n795), .B2(new_n772), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n789), .A2(new_n797), .A3(KEYINPUT53), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n792), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n790), .B1(new_n799), .B2(new_n783), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n716), .A2(new_n412), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n343), .A3(new_n656), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n605), .A2(new_n477), .A3(new_n346), .A4(new_n626), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n627), .A2(new_n669), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n343), .A3(new_n412), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n613), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n569), .A2(new_n516), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n805), .A2(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n802), .A2(new_n669), .ZN(new_n812));
  INV_X1    g626(.A(new_n626), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n477), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n735), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n801), .A2(new_n664), .A3(new_n807), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n701), .A2(new_n703), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n801), .A2(new_n820), .A3(new_n807), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(KEYINPUT48), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n821), .B(new_n823), .Z(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n822), .B2(KEYINPUT48), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(G952), .B(new_n253), .C1(new_n802), .C2(new_n644), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n617), .B2(new_n809), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n826), .B(new_n828), .C1(new_n818), .C2(new_n817), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n800), .A2(new_n829), .B1(G952), .B2(G953), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n343), .A2(new_n477), .A3(new_n345), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n605), .A2(new_n832), .A3(new_n569), .A4(new_n710), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n830), .B1(new_n613), .B2(new_n836), .ZN(G75));
  AOI21_X1  g651(.A(new_n780), .B1(new_n755), .B2(new_n756), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n795), .B2(new_n772), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n288), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(G210), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n400), .B1(new_n403), .B2(new_n398), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT118), .Z(new_n844));
  XNOR2_X1  g658(.A(new_n402), .B(KEYINPUT55), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n841), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n841), .B2(new_n842), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n253), .A2(G952), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G51));
  OAI21_X1  g664(.A(new_n782), .B1(new_n789), .B2(KEYINPUT53), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n790), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n472), .B(KEYINPUT57), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n623), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n722), .B(KEYINPUT119), .Z(new_n857));
  NAND2_X1  g671(.A1(new_n840), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n849), .B1(new_n856), .B2(new_n858), .ZN(G54));
  NAND2_X1  g673(.A1(KEYINPUT58), .A2(G475), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n788), .A2(new_n755), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n862), .B2(new_n791), .ZN(new_n863));
  OAI211_X1 g677(.A(G902), .B(new_n861), .C1(new_n863), .C2(new_n838), .ZN(new_n864));
  INV_X1    g678(.A(new_n510), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n851), .A2(G902), .A3(new_n510), .A4(new_n861), .ZN(new_n869));
  INV_X1    g683(.A(new_n849), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n864), .A2(KEYINPUT120), .A3(new_n865), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n868), .A2(new_n871), .A3(KEYINPUT121), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(G60));
  NAND2_X1  g691(.A1(G478), .A2(G902), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT59), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n566), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT122), .B1(new_n853), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n883), .B(new_n880), .C1(new_n852), .C2(new_n790), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n870), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n566), .B1(new_n800), .B2(new_n879), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(G63));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n545), .A2(new_n288), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n839), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n851), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n893), .A2(new_n335), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n870), .ZN(new_n897));
  INV_X1    g711(.A(new_n584), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n893), .B2(new_n895), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n888), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n895), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n584), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(KEYINPUT61), .A3(new_n870), .A4(new_n896), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(G66));
  NAND2_X1  g718(.A1(new_n415), .A2(G224), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n784), .B2(G953), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n844), .B1(G898), .B2(new_n253), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(G69));
  NOR2_X1   g723(.A1(new_n253), .A2(G900), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n730), .A2(new_n659), .A3(new_n820), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n738), .A2(new_n732), .A3(new_n708), .A4(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n706), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n752), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n914), .B2(new_n253), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n249), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n239), .B2(new_n238), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(new_n506), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(G953), .B1(new_n913), .B2(new_n752), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT126), .B1(new_n922), .B2(new_n910), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n669), .B(new_n602), .C1(new_n570), .C2(new_n577), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n344), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n732), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n732), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n738), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n752), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n615), .A2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n920), .B1(new_n935), .B2(G953), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n924), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n924), .B2(new_n936), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(G72));
  NAND2_X1  g755(.A1(G472), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT63), .Z(new_n943));
  INV_X1    g757(.A(new_n784), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n914), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n298), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n257), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n849), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n943), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n935), .B2(new_n784), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n257), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n799), .ZN(new_n953));
  INV_X1    g767(.A(new_n299), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n949), .B1(new_n954), .B2(new_n261), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(G57));
endmodule


