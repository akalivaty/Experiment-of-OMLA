//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT65), .Z(G319));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(KEYINPUT66), .A3(G137), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n462), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n461), .A2(new_n471), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n478), .B(new_n480), .C1(G124), .C2(new_n481), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n463), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n471), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n481), .A2(G126), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  OR2_X1    g067(.A1(KEYINPUT5), .A2(G543), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT5), .A2(G543), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n495), .A2(G62), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT68), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n496), .B2(KEYINPUT68), .ZN(new_n500));
  OAI21_X1  g075(.A(G651), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(G543), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  OR3_X1    g080(.A1(new_n504), .A2(KEYINPUT67), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT67), .B1(new_n504), .B2(new_n505), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n493), .A2(new_n494), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n506), .A2(new_n507), .B1(G88), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n501), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n495), .A2(new_n514), .A3(G89), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n518), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n515), .A2(KEYINPUT70), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT70), .B1(new_n515), .B2(new_n520), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n514), .B2(G543), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n524), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(G51), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n495), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n523), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n495), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n495), .A2(new_n514), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n504), .A2(KEYINPUT69), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n526), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n539), .B2(new_n526), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n510), .A2(G81), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT71), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(G43), .B1(new_n525), .B2(new_n527), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n510), .A2(G81), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n495), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n534), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n508), .B2(new_n509), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT5), .A2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(KEYINPUT5), .A2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n510), .B2(G91), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n564), .A2(new_n571), .ZN(G299));
  OAI21_X1  g147(.A(KEYINPUT72), .B1(new_n537), .B2(new_n540), .ZN(new_n573));
  NAND2_X1  g148(.A1(G77), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G64), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n568), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n510), .B2(G90), .ZN(new_n577));
  OAI21_X1  g152(.A(G52), .B1(new_n525), .B2(new_n527), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G301));
  INV_X1    g157(.A(KEYINPUT73), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n523), .B2(new_n531), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n539), .A2(new_n526), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G51), .B1(new_n495), .B2(new_n529), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n586), .B(KEYINPUT73), .C1(new_n522), .C2(new_n521), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G286));
  OAI21_X1  g164(.A(G651), .B1(new_n495), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n562), .A2(G49), .ZN(new_n591));
  INV_X1    g166(.A(G87), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n536), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n495), .A2(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(KEYINPUT74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n495), .A2(KEYINPUT74), .A3(G61), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n510), .A2(G86), .B1(new_n562), .B2(G48), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n585), .A2(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n568), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(new_n510), .B2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G290));
  XNOR2_X1  g182(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n536), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n510), .A2(G92), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n568), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n611), .A2(new_n612), .B1(G651), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n585), .A2(G54), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n581), .ZN(G284));
  AOI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n581), .ZN(G321));
  NOR2_X1   g196(.A1(G299), .A2(G868), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n588), .B2(G868), .ZN(G297));
  AOI21_X1  g198(.A(new_n622), .B1(new_n588), .B2(G868), .ZN(G280));
  INV_X1    g199(.A(G860), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n618), .B1(G559), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT76), .ZN(G148));
  OR2_X1    g202(.A1(new_n618), .A2(G559), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g206(.A(new_n461), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n472), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n462), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n481), .A2(G123), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n471), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G2096), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n638), .A3(new_n645), .ZN(G156));
  INV_X1    g221(.A(G14), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT78), .B(G2438), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n661), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n647), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n667));
  INV_X1    g242(.A(new_n664), .ZN(new_n668));
  INV_X1    g243(.A(new_n665), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n669), .C1(new_n662), .C2(new_n663), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n666), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(KEYINPUT81), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(new_n666), .C1(new_n670), .C2(new_n672), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G401));
  XNOR2_X1  g253(.A(G2084), .B(G2090), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT82), .Z(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2072), .B(G2078), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n683), .B(KEYINPUT17), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n683), .B(KEYINPUT84), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(new_n644), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT85), .B(G2100), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT86), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1961), .B(G1966), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT19), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT20), .Z(new_n704));
  NOR2_X1   g279(.A1(new_n697), .A2(new_n699), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n706), .A2(new_n702), .A3(new_n700), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n704), .B(new_n707), .C1(new_n702), .C2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n714), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(G229));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G22), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT88), .Z(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G303), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1971), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(G6), .A2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G305), .B2(new_n718), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT32), .B(G1981), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n721), .A2(new_n722), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n723), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n718), .A2(G23), .ZN(new_n730));
  INV_X1    g305(.A(G288), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n718), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT33), .B(G1976), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n725), .B2(new_n726), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n729), .A2(KEYINPUT34), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n718), .A2(G24), .ZN(new_n737));
  INV_X1    g312(.A(G290), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n718), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1986), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G25), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n462), .A2(G131), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT87), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n481), .A2(G119), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n471), .A2(G107), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n742), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT35), .B(G1991), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n736), .A2(new_n740), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT89), .ZN(new_n753));
  OR2_X1    g328(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT34), .B1(new_n729), .B2(new_n735), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(G164), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G27), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G34), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n762), .B2(KEYINPUT24), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(KEYINPUT24), .B2(new_n762), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n474), .B2(new_n741), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  NOR2_X1   g343(.A1(G171), .A2(new_n718), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G5), .B2(new_n718), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n761), .B(new_n767), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n768), .ZN(new_n772));
  AOI21_X1  g347(.A(KEYINPUT23), .B1(new_n718), .B2(G20), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n718), .A2(KEYINPUT23), .A3(G20), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n773), .B(new_n774), .C1(G299), .C2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT95), .B(G1956), .Z(new_n776));
  OAI22_X1  g351(.A1(new_n759), .A2(new_n760), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n772), .B(new_n777), .C1(new_n775), .C2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n741), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n741), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT29), .B(G2090), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n741), .A2(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT25), .Z(new_n785));
  INV_X1    g360(.A(G139), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n463), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n632), .A2(G127), .ZN(new_n788));
  NAND2_X1  g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n471), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n783), .B1(new_n791), .B2(new_n741), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G2072), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT30), .B(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  NAND2_X1  g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n794), .A2(new_n741), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n793), .B(new_n797), .C1(new_n741), .C2(new_n643), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n462), .A2(G140), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n481), .A2(G128), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n471), .A2(G116), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n741), .A2(G26), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT28), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT92), .B(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n792), .A2(G2072), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n782), .A2(new_n798), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G4), .A2(G16), .ZN(new_n812));
  INV_X1    g387(.A(new_n618), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT91), .B(G1348), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n771), .A2(new_n778), .A3(new_n811), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n741), .A2(G32), .ZN(new_n818));
  NAND3_X1  g393(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT26), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G129), .B2(new_n481), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n462), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n824), .B2(new_n741), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT93), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT27), .B(G1996), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n586), .B1(new_n522), .B2(new_n521), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(new_n718), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT94), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G16), .B2(G21), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n831), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G1966), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(G1966), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n828), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(G16), .A2(G19), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n555), .B2(G16), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1341), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n817), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n757), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(G311));
  INV_X1    g419(.A(G311), .ZN(G150));
  NAND2_X1  g420(.A1(G80), .A2(G543), .ZN(new_n846));
  INV_X1    g421(.A(G67), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n568), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n848), .A2(G651), .B1(new_n510), .B2(G93), .ZN(new_n849));
  OAI21_X1  g424(.A(G55), .B1(new_n525), .B2(new_n527), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G860), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT97), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n813), .A2(G559), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI211_X1 g432(.A(new_n552), .B(new_n851), .C1(new_n545), .C2(new_n549), .ZN(new_n858));
  INV_X1    g433(.A(new_n851), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n550), .B2(new_n553), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n857), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n625), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n854), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT98), .Z(G145));
  XNOR2_X1  g442(.A(new_n748), .B(new_n634), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n481), .A2(G130), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n871), .A2(new_n471), .A3(G118), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n471), .B2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n872), .B(new_n873), .C1(KEYINPUT101), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(KEYINPUT101), .B2(new_n874), .ZN(new_n876));
  AOI211_X1 g451(.A(new_n870), .B(new_n876), .C1(G142), .C2(new_n462), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n868), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n791), .B(new_n823), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(new_n803), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n803), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n491), .A2(KEYINPUT99), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n485), .A2(new_n885), .A3(new_n486), .A4(new_n490), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n881), .A2(new_n884), .A3(new_n886), .A4(new_n882), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G162), .B(new_n643), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G160), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(KEYINPUT102), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n888), .A2(new_n896), .A3(new_n889), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT103), .B1(new_n898), .B2(new_n879), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n900));
  AOI211_X1 g475(.A(new_n900), .B(new_n878), .C1(new_n895), .C2(new_n897), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n894), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n878), .B1(new_n889), .B2(new_n888), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n893), .B1(new_n891), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g482(.A1(new_n618), .A2(G299), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n618), .A2(G299), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n911), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n917), .B2(KEYINPUT104), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n861), .B(new_n628), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n908), .A2(new_n910), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n922), .B2(new_n919), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n924));
  XNOR2_X1  g499(.A(G303), .B(new_n738), .ZN(new_n925));
  XNOR2_X1  g500(.A(G305), .B(new_n731), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n924), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n924), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(G868), .B2(new_n859), .ZN(G295));
  OAI21_X1  g508(.A(new_n932), .B1(G868), .B2(new_n859), .ZN(G331));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n581), .B2(new_n829), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n584), .A2(G171), .A3(new_n587), .ZN(new_n937));
  NAND4_X1  g512(.A1(G168), .A2(KEYINPUT105), .A3(new_n573), .A4(new_n580), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n858), .A2(new_n860), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n861), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n917), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n922), .B1(new_n942), .B2(new_n861), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(new_n861), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n921), .B1(new_n939), .B2(new_n940), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n942), .A2(new_n861), .A3(new_n948), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n948), .B1(new_n942), .B2(new_n861), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n953), .B(new_n951), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n928), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n941), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  INV_X1    g534(.A(new_n911), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n915), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n913), .B1(new_n961), .B2(new_n912), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n959), .A2(new_n962), .B1(new_n943), .B2(new_n953), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n963), .B2(new_n927), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n958), .A2(new_n964), .A3(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n953), .A2(new_n943), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n942), .A2(new_n861), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n947), .B2(new_n949), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n927), .B(new_n967), .C1(new_n969), .C2(new_n918), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n903), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n959), .A2(new_n962), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n927), .B1(new_n972), .B2(new_n967), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n966), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT44), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n978), .A2(KEYINPUT107), .B1(new_n917), .B2(new_n944), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n927), .B1(new_n979), .B2(new_n956), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n980), .A2(new_n971), .A3(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n972), .A2(new_n967), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n928), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n966), .B1(new_n964), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n977), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n976), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n977), .B1(new_n965), .B2(new_n974), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n958), .A2(new_n964), .A3(new_n966), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n971), .B2(new_n973), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT44), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT108), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n987), .A2(new_n992), .ZN(G397));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n884), .A2(new_n994), .A3(new_n886), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n467), .A2(G40), .A3(new_n473), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n803), .B(G2067), .Z(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n823), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1000), .A2(G1996), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1000), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1005), .B2(new_n824), .ZN(new_n1012));
  NOR4_X1   g587(.A1(new_n1000), .A2(KEYINPUT111), .A3(G1996), .A4(new_n823), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1003), .B1(G1996), .B2(new_n823), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1012), .A2(new_n1013), .B1(new_n1000), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(KEYINPUT112), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(KEYINPUT112), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n748), .B(new_n750), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT113), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n1001), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1986), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n738), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT110), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1000), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT48), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1010), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n750), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n748), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1016), .A2(new_n1017), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n803), .A2(G2067), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1000), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2090), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n491), .A2(new_n994), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n491), .B2(new_n994), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1036), .A2(new_n998), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n994), .A4(new_n886), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n996), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n999), .A3(new_n1041), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1034), .A2(new_n1039), .B1(new_n1042), .B2(new_n722), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(G303), .B2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G166), .A2(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1051), .A3(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1035), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1047), .B1(new_n1053), .B2(new_n999), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n731), .A2(G1976), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1054), .A2(KEYINPUT116), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n1059));
  OAI211_X1 g634(.A(G8), .B(new_n1055), .C1(new_n1035), .C2(new_n998), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1057), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G305), .A2(G1981), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n599), .B2(new_n600), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n1064), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1054), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n1060), .B2(KEYINPUT52), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1060), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1063), .B(new_n1071), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1054), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1064), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1052), .A2(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1071), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1063), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1050), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1082));
  INV_X1    g657(.A(new_n996), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n491), .A2(KEYINPUT118), .A3(new_n994), .A4(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n999), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT45), .B1(new_n491), .B2(new_n994), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1086), .A2(new_n1087), .B1(new_n1035), .B2(new_n996), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1966), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1089), .A2(new_n1090), .B1(new_n1039), .B2(new_n766), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1091), .A2(new_n1047), .A3(G286), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1081), .A2(new_n1082), .A3(new_n1052), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1044), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1098), .A3(new_n1050), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1043), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1074), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1099), .A2(new_n1101), .A3(KEYINPUT63), .A4(new_n1092), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1078), .B1(new_n1095), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1047), .B1(new_n1091), .B2(G168), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1038), .A2(new_n998), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(KEYINPUT50), .B2(new_n1035), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(G2084), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1966), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n829), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT51), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  AOI211_X1 g687(.A(KEYINPUT51), .B(new_n1047), .C1(new_n1091), .C2(G168), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1082), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1040), .A2(new_n760), .A3(new_n999), .A4(new_n1041), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n768), .A2(new_n1106), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1085), .A2(new_n1088), .A3(KEYINPUT53), .A4(new_n760), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n581), .ZN(new_n1122));
  NOR4_X1   g697(.A1(new_n1116), .A2(new_n1122), .A3(new_n1074), .A4(new_n1100), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT62), .B1(new_n1125), .B2(new_n1113), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1115), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1103), .A2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1039), .A2(G1956), .ZN(new_n1129));
  NAND2_X1  g704(.A1(G299), .A2(KEYINPUT120), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT57), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1040), .A2(new_n999), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1041), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1131), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1053), .A2(new_n999), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(G2067), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n815), .B2(new_n1106), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n618), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1136), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1135), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT121), .B(G1996), .Z(new_n1147));
  NAND3_X1  g722(.A1(new_n1132), .A2(new_n1041), .A3(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n1137), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g725(.A(new_n554), .B(new_n1146), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1139), .A2(KEYINPUT60), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n813), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1154), .A2(new_n1155), .A3(new_n618), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1139), .A2(KEYINPUT60), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1145), .B(new_n1153), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1142), .A2(KEYINPUT61), .A3(new_n1135), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT123), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1141), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1119), .A2(new_n1120), .A3(G301), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1119), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n760), .A2(KEYINPUT53), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n995), .B2(new_n996), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1169), .B1(new_n1132), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1132), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1168), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(G171), .ZN(new_n1176));
  OAI211_X1 g751(.A(KEYINPUT54), .B(new_n1167), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1116), .A2(new_n1074), .A3(new_n1100), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1166), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1174), .ZN(new_n1180));
  OAI211_X1 g755(.A(G301), .B(new_n1119), .C1(new_n1180), .C2(new_n1172), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT54), .B1(new_n1122), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1179), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1128), .B1(new_n1165), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1024), .B1(new_n1022), .B2(new_n738), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1001), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1016), .A2(new_n1189), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1033), .B1(new_n1187), .B2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g766(.A1(new_n989), .A2(new_n990), .ZN(new_n1193));
  INV_X1    g767(.A(new_n456), .ZN(new_n1194));
  OR2_X1    g768(.A1(G227), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1195), .B1(new_n715), .B2(new_n716), .ZN(new_n1196));
  AND4_X1   g770(.A1(new_n677), .A2(new_n1193), .A3(new_n906), .A4(new_n1196), .ZN(G308));
  NAND4_X1  g771(.A1(new_n677), .A2(new_n906), .A3(new_n1193), .A4(new_n1196), .ZN(G225));
endmodule


