//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(KEYINPUT1), .A3(G146), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n193), .B(new_n194), .C1(G128), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT0), .B(G128), .Z(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n198), .B1(new_n203), .B2(new_n197), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n205), .A2(KEYINPUT89), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G224), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G953), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(new_n205), .ZN(new_n210));
  XOR2_X1   g024(.A(new_n207), .B(new_n210), .Z(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT3), .A3(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n215), .B2(G104), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(KEYINPUT75), .A3(G107), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n213), .A2(G107), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n215), .A2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT2), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT2), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G113), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G116), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G119), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT5), .ZN(new_n238));
  OAI21_X1  g052(.A(G113), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n233), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n226), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(G110), .B(G122), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT8), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n232), .A2(KEYINPUT5), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(KEYINPUT86), .A3(new_n245), .A4(G113), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n238), .B2(new_n239), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n248), .A3(new_n233), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n241), .B(new_n243), .C1(new_n226), .C2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n250), .A2(KEYINPUT88), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(KEYINPUT88), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n211), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G101), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT76), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n222), .A3(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n254), .B(G101), .C1(KEYINPUT76), .C2(new_n256), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n235), .A2(new_n237), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT2), .B(G113), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n233), .B2(new_n265), .ZN(new_n266));
  AOI211_X1 g080(.A(KEYINPUT68), .B(KEYINPUT69), .C1(new_n231), .C2(new_n232), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n265), .B1(new_n261), .B2(new_n262), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n233), .A2(new_n265), .A3(new_n264), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n270), .A2(new_n261), .A3(new_n271), .A4(new_n262), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n260), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n222), .A2(new_n225), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n249), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n277), .A3(new_n242), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT87), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n276), .B1(new_n260), .B2(new_n273), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT87), .A3(new_n242), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n253), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n281), .A2(new_n242), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT6), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n281), .A2(new_n242), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n281), .A2(KEYINPUT87), .A3(new_n242), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT87), .B1(new_n281), .B2(new_n242), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n290), .B2(KEYINPUT6), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n204), .B(new_n209), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n284), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n295), .B(new_n284), .C1(new_n291), .C2(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n300), .B(KEYINPUT85), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n197), .A2(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT19), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G125), .B(G140), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT19), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n189), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT16), .ZN(new_n314));
  OR3_X1    g128(.A1(new_n197), .A2(KEYINPUT16), .A3(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G146), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n307), .A2(new_n308), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n310), .A2(KEYINPUT19), .ZN(new_n319));
  AOI21_X1  g133(.A(G146), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n316), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT91), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G237), .A2(G953), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(G143), .A3(G214), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(G143), .B1(new_n323), .B2(G214), .ZN(new_n326));
  OAI21_X1  g140(.A(G131), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n324), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n317), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n310), .B(new_n189), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT18), .B(G131), .C1(new_n325), .C2(new_n326), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT18), .A2(G131), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n328), .A2(new_n324), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT93), .ZN(new_n339));
  XOR2_X1   g153(.A(G113), .B(G122), .Z(new_n340));
  XOR2_X1   g154(.A(KEYINPUT92), .B(G104), .Z(new_n341));
  XOR2_X1   g155(.A(new_n340), .B(new_n341), .Z(new_n342));
  NAND3_X1  g156(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(G475), .A2(G902), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT94), .ZN(new_n345));
  INV_X1    g159(.A(new_n342), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n332), .B2(new_n337), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n331), .A2(KEYINPUT17), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n314), .A2(new_n315), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n189), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n350), .B(new_n316), .C1(new_n327), .C2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n346), .B(new_n337), .C1(new_n348), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT93), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n343), .B(new_n345), .C1(new_n347), .C2(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n354), .A2(new_n347), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n343), .A4(new_n345), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G475), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n337), .B1(new_n348), .B2(new_n352), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n342), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n353), .ZN(new_n366));
  INV_X1    g180(.A(G902), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n191), .A3(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n191), .A2(G128), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n187), .A2(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(G134), .B(new_n372), .C1(new_n375), .C2(new_n371), .ZN(new_n376));
  XNOR2_X1  g190(.A(G116), .B(G122), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G107), .ZN(new_n378));
  INV_X1    g192(.A(G122), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n236), .A2(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n215), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n375), .A2(KEYINPUT95), .ZN(new_n385));
  XNOR2_X1  g199(.A(G128), .B(G143), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT95), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(G134), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT96), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G134), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n375), .A2(KEYINPUT95), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n383), .A2(new_n378), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT96), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .A4(new_n376), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n385), .A2(new_n388), .A3(G134), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n215), .B1(new_n380), .B2(KEYINPUT14), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n377), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT9), .B(G234), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G953), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(G217), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n398), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n398), .B2(new_n403), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT97), .B(new_n367), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G478), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(KEYINPUT15), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n411), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n370), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G952), .ZN(new_n416));
  AOI211_X1 g230(.A(G953), .B(new_n416), .C1(G234), .C2(G237), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G234), .ZN(new_n419));
  INV_X1    g233(.A(G237), .ZN(new_n420));
  OAI211_X1 g234(.A(G902), .B(G953), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT98), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n418), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n303), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n406), .A2(G227), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n226), .A2(new_n196), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n432));
  AOI21_X1  g246(.A(G128), .B1(new_n190), .B2(new_n192), .ZN(new_n433));
  INV_X1    g247(.A(new_n194), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT77), .B(new_n194), .C1(new_n195), .C2(G128), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n435), .A2(new_n193), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT78), .B1(new_n437), .B2(new_n275), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n193), .A3(new_n436), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n226), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n431), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  OR2_X1    g256(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n443));
  INV_X1    g257(.A(G137), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G134), .ZN(new_n445));
  NAND2_X1  g259(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(KEYINPUT65), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G137), .ZN(new_n450));
  AND2_X1   g264(.A1(KEYINPUT11), .A2(G134), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n444), .A2(G134), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G131), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n447), .A2(new_n452), .A3(new_n329), .A4(new_n454), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT81), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n442), .A2(KEYINPUT12), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n226), .A2(new_n439), .A3(new_n440), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n440), .B1(new_n226), .B2(new_n439), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n196), .B2(new_n226), .ZN(new_n464));
  INV_X1    g278(.A(new_n459), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n458), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n196), .A2(KEYINPUT10), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n226), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n258), .A2(new_n259), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n203), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n438), .A2(new_n441), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT80), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT80), .ZN(new_n478));
  AOI211_X1 g292(.A(new_n478), .B(new_n475), .C1(new_n438), .C2(new_n441), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n468), .B(new_n473), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n467), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n467), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n430), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n476), .B1(new_n462), .B2(new_n463), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n478), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n474), .A2(KEYINPUT80), .A3(new_n476), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n472), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT83), .B1(new_n488), .B2(new_n468), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n458), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n430), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n480), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n484), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT84), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n458), .B(new_n472), .C1(new_n486), .C2(new_n487), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT12), .B1(new_n442), .B2(new_n459), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n464), .A2(new_n461), .A3(new_n465), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT82), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n467), .A2(new_n480), .A3(new_n481), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n494), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n495), .B1(new_n492), .B2(new_n489), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n367), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT84), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(G469), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n496), .A2(new_n467), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n501), .B1(new_n489), .B2(new_n492), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n494), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n499), .A3(new_n367), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n500), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n350), .A2(new_n316), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n234), .A2(G128), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n234), .A2(G128), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n187), .A2(G119), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT24), .B(G110), .Z(new_n524));
  AOI22_X1  g338(.A1(new_n521), .A2(G110), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  OAI22_X1  g340(.A1(new_n521), .A2(G110), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n316), .C1(G146), .C2(new_n307), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT22), .B(G137), .ZN(new_n530));
  INV_X1    g344(.A(G221), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n531), .A2(new_n419), .A3(G953), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n530), .B(new_n532), .Z(new_n533));
  XNOR2_X1  g347(.A(new_n529), .B(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n534), .B(new_n367), .C1(KEYINPUT74), .C2(KEYINPUT25), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT74), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G217), .B1(new_n419), .B2(G902), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n535), .B2(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n367), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n539), .A2(new_n541), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n196), .A2(new_n457), .ZN(new_n547));
  AOI21_X1  g361(.A(G134), .B1(new_n448), .B2(new_n450), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n445), .B1(new_n548), .B2(KEYINPUT67), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT65), .B(G137), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT67), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n550), .A2(new_n551), .A3(G134), .ZN(new_n552));
  OAI21_X1  g366(.A(G131), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n453), .B1(new_n550), .B2(new_n451), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n329), .B1(new_n555), .B2(new_n447), .ZN(new_n556));
  AND4_X1   g370(.A1(new_n329), .A2(new_n447), .A3(new_n452), .A4(new_n454), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n202), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(KEYINPUT30), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n196), .A2(new_n457), .ZN(new_n560));
  INV_X1    g374(.A(new_n552), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n551), .B1(new_n550), .B2(G134), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n445), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n563), .B2(G131), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT66), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n458), .A2(KEYINPUT66), .A3(new_n202), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n273), .B(new_n559), .C1(new_n568), .C2(KEYINPUT30), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n554), .A2(new_n558), .A3(new_n272), .A4(new_n268), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT71), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n420), .A2(new_n406), .A3(G210), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT26), .B(G101), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n571), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n572), .B1(new_n571), .B2(new_n578), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n546), .B1(new_n570), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n571), .A2(new_n578), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT71), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n571), .A2(new_n578), .A3(new_n572), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(KEYINPUT31), .A3(new_n569), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT28), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n571), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n571), .ZN(new_n590));
  INV_X1    g404(.A(new_n567), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT66), .B1(new_n458), .B2(new_n202), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n554), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n593), .B2(new_n273), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n582), .A2(new_n587), .B1(new_n577), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(G472), .A2(G902), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT32), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n596), .A2(new_n577), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n586), .A2(KEYINPUT31), .A3(new_n569), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT31), .B1(new_n586), .B2(new_n569), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT32), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n598), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT29), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(new_n589), .C1(new_n594), .C2(new_n595), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n589), .A2(KEYINPUT73), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n554), .A2(new_n558), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n273), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n588), .B1(new_n613), .B2(new_n571), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n589), .A2(KEYINPUT73), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n610), .B(new_n578), .C1(new_n616), .C2(new_n609), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n569), .A2(new_n609), .A3(new_n577), .A4(new_n571), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n618), .A2(new_n367), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n608), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n545), .B1(new_n607), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n531), .B1(new_n405), .B2(new_n367), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n427), .A2(new_n516), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  AND2_X1   g440(.A1(new_n516), .A2(new_n624), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n597), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n604), .A2(new_n598), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n628), .A2(new_n629), .A3(new_n544), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n390), .A2(new_n397), .B1(new_n400), .B2(new_n402), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT99), .B1(new_n633), .B2(new_n408), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n634), .B(KEYINPUT33), .C1(new_n409), .C2(new_n410), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n398), .A2(new_n403), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n407), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n408), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n637), .B(new_n638), .C1(KEYINPUT99), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n412), .A2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n367), .B1(new_n409), .B2(new_n410), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n412), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n641), .A2(new_n644), .A3(new_n642), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n368), .B1(new_n358), .B2(new_n361), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n632), .A2(new_n425), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n631), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  NAND3_X1  g469(.A1(new_n299), .A2(new_n302), .A3(new_n425), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n359), .A2(new_n356), .A3(new_n343), .A4(new_n345), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n368), .B1(new_n358), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n414), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n631), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NAND2_X1  g477(.A1(new_n539), .A2(new_n541), .ZN(new_n664));
  INV_X1    g478(.A(new_n533), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n529), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n543), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n628), .A2(new_n629), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n672), .A2(new_n624), .A3(new_n516), .A4(new_n427), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT37), .B(G110), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  AOI21_X1  g491(.A(new_n620), .B1(new_n600), .B2(new_n606), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n418), .B1(new_n422), .B2(G900), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n658), .A2(new_n414), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n658), .A2(KEYINPUT104), .A3(new_n414), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n669), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n678), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n516), .A2(new_n686), .A3(new_n624), .A4(new_n632), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT105), .B(G128), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G30));
  XNOR2_X1  g503(.A(new_n679), .B(KEYINPUT39), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n627), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n692));
  INV_X1    g506(.A(new_n413), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n411), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n650), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n685), .A2(new_n695), .A3(new_n302), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT106), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n299), .B(KEYINPUT38), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n570), .A2(new_n581), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n578), .B1(new_n613), .B2(new_n571), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n367), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G472), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n607), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n697), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n691), .B2(KEYINPUT40), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n692), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n191), .ZN(G45));
  AND4_X1   g521(.A1(new_n370), .A2(new_n647), .A3(new_n648), .A4(new_n679), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n678), .A2(new_n709), .A3(new_n685), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n516), .A2(new_n710), .A3(new_n624), .A4(new_n632), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND2_X1  g526(.A1(new_n514), .A2(new_n367), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n714), .A2(new_n624), .A3(new_n515), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n652), .A3(new_n622), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND3_X1  g532(.A1(new_n660), .A2(new_n715), .A3(new_n622), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  AND4_X1   g534(.A1(new_n624), .A2(new_n714), .A3(new_n632), .A4(new_n515), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n678), .A2(new_n426), .A3(new_n685), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  INV_X1    g538(.A(new_n695), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n602), .A2(new_n603), .B1(new_n578), .B2(new_n616), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n598), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n628), .A2(new_n727), .A3(new_n544), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n656), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n715), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NAND3_X1  g545(.A1(new_n628), .A2(new_n669), .A3(new_n727), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n709), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n721), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G125), .ZN(G27));
  OAI21_X1  g549(.A(new_n515), .B1(new_n499), .B2(new_n498), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n623), .A2(new_n301), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n297), .A2(new_n298), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n708), .A2(new_n740), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n622), .A2(new_n736), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n509), .A2(G469), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n738), .B1(new_n743), .B2(new_n515), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n597), .A2(KEYINPUT32), .A3(new_n599), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n605), .B1(new_n604), .B2(new_n598), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n600), .A2(KEYINPUT107), .A3(new_n606), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n621), .A3(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n744), .A2(new_n750), .A3(new_n544), .A4(new_n708), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n742), .B1(KEYINPUT42), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  INV_X1    g567(.A(new_n684), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n622), .A2(new_n736), .A3(new_n739), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n507), .B2(new_n508), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n484), .A2(KEYINPUT45), .A3(new_n497), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(G469), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(G469), .A2(G902), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT108), .B1(new_n762), .B2(KEYINPUT46), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(KEYINPUT46), .A3(new_n761), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n515), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT46), .B1(new_n760), .B2(new_n761), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n763), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n647), .A2(new_n650), .A3(new_n648), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT43), .B1(new_n650), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n770), .B(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n685), .B1(new_n628), .B2(new_n629), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT44), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT44), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n297), .A2(new_n302), .A3(new_n298), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n769), .A2(new_n624), .A3(new_n690), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  INV_X1    g594(.A(new_n678), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n781), .A2(new_n777), .A3(new_n709), .A4(new_n544), .ZN(new_n782));
  INV_X1    g596(.A(new_n768), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n515), .B(new_n764), .C1(new_n766), .C2(new_n767), .ZN(new_n784));
  OAI211_X1 g598(.A(KEYINPUT47), .B(new_n624), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT47), .B1(new_n769), .B2(new_n624), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  AND3_X1   g603(.A1(new_n734), .A2(new_n711), .A3(new_n687), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n303), .A2(new_n725), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n685), .A2(new_n624), .A3(new_n679), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n703), .A3(new_n736), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n687), .A2(new_n734), .A3(new_n711), .A4(new_n794), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n733), .A2(new_n736), .A3(new_n739), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n755), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n750), .A2(new_n544), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n736), .A2(new_n739), .A3(new_n708), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT42), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n742), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n658), .A2(new_n694), .A3(new_n679), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n297), .A2(new_n298), .A3(new_n302), .A4(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n678), .A3(new_n685), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n516), .A3(new_n624), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n730), .A2(new_n719), .A3(new_n723), .A4(new_n716), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n415), .B1(new_n370), .B2(new_n649), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n656), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n516), .A3(new_n624), .A4(new_n630), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n673), .A2(new_n815), .A3(new_n625), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT113), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n809), .A2(new_n810), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n798), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n807), .A2(new_n624), .A3(new_n516), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n755), .A2(new_n799), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n622), .A2(new_n624), .A3(new_n515), .A4(new_n714), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n828), .A2(new_n652), .B1(new_n729), .B2(new_n715), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n828), .A2(new_n660), .B1(new_n721), .B2(new_n722), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n827), .A2(new_n752), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n816), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n791), .B1(new_n734), .B2(new_n687), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n822), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n798), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n823), .A2(new_n824), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n821), .B1(new_n822), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n823), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n836), .B1(new_n840), .B2(new_n824), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n773), .A2(new_n417), .ZN(new_n843));
  INV_X1    g657(.A(new_n728), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n777), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n786), .A2(new_n787), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n714), .A2(new_n515), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n623), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n849), .B2(KEYINPUT114), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n848), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n698), .A2(new_n302), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n845), .A2(new_n715), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT50), .Z(new_n857));
  AND3_X1   g671(.A1(new_n851), .A2(new_n417), .A3(new_n739), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n607), .A2(new_n858), .A3(new_n544), .A4(new_n702), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n650), .A3(new_n649), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n773), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n857), .B(new_n860), .C1(new_n732), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n842), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n406), .A2(KEYINPUT115), .A3(G952), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(KEYINPUT115), .B2(new_n406), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n859), .B2(new_n651), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n861), .A2(new_n801), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(KEYINPUT116), .A3(KEYINPUT48), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n845), .A2(new_n721), .ZN(new_n869));
  XOR2_X1   g683(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n861), .B2(new_n801), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n866), .A2(new_n868), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n862), .A2(new_n842), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n847), .B1(new_n849), .B2(new_n852), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n863), .A2(new_n875), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n841), .A2(new_n876), .B1(G952), .B2(G953), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n770), .A2(new_n545), .A3(new_n623), .A4(new_n301), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT110), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT49), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n851), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT111), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n703), .B(new_n698), .C1(new_n880), .C2(new_n851), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT112), .Z(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n885), .ZN(G75));
  NAND2_X1  g700(.A1(new_n795), .A2(new_n797), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n819), .B1(new_n831), .B2(new_n816), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n803), .A2(new_n800), .A3(new_n804), .A4(new_n808), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n716), .A2(new_n730), .A3(new_n719), .A4(new_n723), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(KEYINPUT113), .A3(new_n817), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n887), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n835), .B1(new_n892), .B2(KEYINPUT53), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(G210), .A3(G902), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n291), .B(new_n292), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT55), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n894), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n406), .A2(G952), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(new_n761), .B(KEYINPUT117), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT57), .ZN(new_n903));
  INV_X1    g717(.A(new_n836), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n824), .B1(new_n823), .B2(new_n835), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n514), .ZN(new_n907));
  INV_X1    g721(.A(new_n760), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n893), .A2(G902), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n900), .B1(new_n907), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n359), .A2(new_n343), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n900), .ZN(G60));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n641), .B1(new_n841), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n641), .B(new_n918), .C1(new_n904), .C2(new_n905), .ZN(new_n920));
  INV_X1    g734(.A(new_n900), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n922), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT60), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n823), .B2(new_n835), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n924), .B(new_n921), .C1(new_n927), .C2(new_n534), .ZN(new_n928));
  INV_X1    g742(.A(new_n926), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n534), .B1(new_n893), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT118), .B1(new_n930), .B2(new_n900), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n667), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n930), .A2(KEYINPUT119), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n930), .A2(KEYINPUT119), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n900), .A2(new_n934), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n936), .A2(new_n932), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n935), .A2(new_n939), .ZN(G66));
  NAND2_X1  g754(.A1(new_n890), .A2(new_n817), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n406), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n423), .B2(new_n208), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n291), .B1(G898), .B2(new_n406), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G69));
  INV_X1    g760(.A(new_n790), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT62), .B1(new_n706), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n813), .A2(new_n777), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n627), .A2(new_n622), .A3(new_n690), .A4(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n779), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n952), .B(new_n790), .C1(new_n692), .C2(new_n705), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n948), .A2(new_n788), .A3(new_n951), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n406), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n559), .B1(new_n568), .B2(KEYINPUT30), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT120), .Z(new_n957));
  NOR2_X1   g771(.A1(new_n309), .A2(new_n311), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(new_n959));
  NAND2_X1  g773(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n779), .A2(new_n790), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n803), .A2(new_n804), .A3(new_n755), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n752), .A2(new_n964), .A3(new_n755), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n788), .A2(new_n961), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n801), .A2(new_n303), .A3(new_n725), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n769), .A2(new_n624), .A3(new_n690), .A4(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n406), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n406), .A2(G900), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT122), .Z(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(KEYINPUT125), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n959), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT125), .B1(new_n972), .B2(new_n974), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n960), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT121), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n977), .B2(new_n978), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n406), .B1(G227), .B2(G900), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  OAI221_X1 g798(.A(new_n960), .B1(new_n980), .B2(new_n982), .C1(new_n977), .C2(new_n978), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OR2_X1    g802(.A1(new_n967), .A2(new_n971), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n941), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n570), .A2(new_n590), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n577), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n988), .B1(new_n954), .B2(new_n941), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n991), .A2(new_n577), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n900), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n840), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n991), .A2(new_n578), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n988), .B1(new_n998), .B2(new_n699), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n997), .A2(KEYINPUT127), .A3(new_n1000), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(G57));
endmodule


