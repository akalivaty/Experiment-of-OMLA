//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n642, new_n643, new_n644,
    new_n647, new_n649, new_n650, new_n651, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n469), .B(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G101), .A3(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n478), .A2(KEYINPUT70), .A3(G101), .A4(G2104), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n477), .A2(G137), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OAI21_X1  g060(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G112), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(G136), .B2(new_n477), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  OAI211_X1 g074(.A(G138), .B(new_n478), .C1(new_n464), .C2(new_n465), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n488), .A2(new_n502), .A3(G138), .A4(new_n478), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n478), .A2(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(G114), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n508), .A2(new_n510), .A3(new_n511), .A4(G2104), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n478), .B1(new_n475), .B2(new_n476), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n507), .A2(new_n512), .B1(new_n513), .B2(G126), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n504), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n522), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n536), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(KEYINPUT6), .A2(G651), .ZN(new_n539));
  NOR2_X1   g114(.A1(KEYINPUT6), .A2(G651), .ZN(new_n540));
  OAI211_X1 g115(.A(G51), .B(G543), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G89), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n524), .B2(new_n525), .ZN(new_n544));
  NAND2_X1  g119(.A1(G63), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n519), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G168));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n517), .B2(new_n518), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(KEYINPUT5), .A2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT5), .A2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g133(.A(KEYINPUT73), .B(new_n553), .C1(new_n558), .C2(new_n551), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(G651), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n519), .A2(new_n529), .A3(G90), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n529), .A2(G52), .A3(G543), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n563), .B1(new_n561), .B2(new_n562), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(G301));
  INV_X1    g141(.A(G301), .ZN(G171));
  AOI22_X1  g142(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n521), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n526), .A2(G43), .ZN(new_n570));
  INV_X1    g145(.A(G81), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n530), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(G188));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT76), .B(new_n579), .C1(new_n558), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n519), .A2(G65), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT76), .B1(new_n583), .B2(new_n579), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT77), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n580), .B1(new_n517), .B2(new_n518), .ZN(new_n587));
  INV_X1    g162(.A(new_n579), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n589), .A2(new_n581), .A3(new_n590), .A4(G651), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n526), .B2(G53), .ZN(new_n594));
  OAI211_X1 g169(.A(G53), .B(G543), .C1(new_n539), .C2(new_n540), .ZN(new_n595));
  INV_X1    g170(.A(new_n593), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G91), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n594), .A2(new_n597), .B1(new_n598), .B2(new_n530), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT78), .B1(new_n592), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n602));
  AOI211_X1 g177(.A(new_n602), .B(new_n599), .C1(new_n585), .C2(new_n591), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n601), .A2(new_n603), .ZN(G299));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n542), .A2(new_n547), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(G89), .B1(new_n539), .B2(new_n540), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n558), .B1(new_n607), .B2(new_n545), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n538), .A2(new_n541), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT79), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(G286));
  INV_X1    g187(.A(new_n530), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G87), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n526), .A2(G49), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(G288));
  INV_X1    g192(.A(G86), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n530), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT80), .ZN(new_n620));
  NAND2_X1  g195(.A1(G73), .A2(G543), .ZN(new_n621));
  INV_X1    g196(.A(G61), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n558), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n623), .A2(G651), .B1(G48), .B2(new_n526), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n530), .B2(new_n618), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n624), .A3(new_n626), .ZN(G305));
  AOI22_X1  g202(.A1(new_n613), .A2(G85), .B1(G47), .B2(new_n526), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n521), .B2(new_n629), .ZN(G290));
  NAND2_X1  g205(.A1(G301), .A2(G868), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n519), .A2(new_n529), .A3(G92), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g208(.A1(G79), .A2(G543), .ZN(new_n634));
  INV_X1    g209(.A(G66), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n558), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n636), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n631), .B1(new_n639), .B2(G868), .ZN(G321));
  XNOR2_X1  g215(.A(G321), .B(KEYINPUT81), .ZN(G284));
  INV_X1    g216(.A(G868), .ZN(new_n642));
  NOR2_X1   g217(.A1(G286), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G299), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n642), .ZN(G280));
  XOR2_X1   g220(.A(G280), .B(KEYINPUT82), .Z(G297));
  INV_X1    g221(.A(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n639), .B1(new_n647), .B2(G860), .ZN(G148));
  OR2_X1    g223(.A1(new_n569), .A2(new_n572), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(new_n642), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n638), .A2(G559), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n651), .B2(new_n642), .ZN(G323));
  XOR2_X1   g227(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n653));
  XNOR2_X1  g228(.A(G323), .B(new_n653), .ZN(G282));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  INV_X1    g230(.A(G111), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n655), .B1(new_n656), .B2(G2105), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(G135), .B2(new_n477), .ZN(new_n658));
  INV_X1    g233(.A(G123), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n491), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT85), .B(G2096), .Z(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT12), .Z(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT13), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n667), .A3(new_n668), .ZN(G156));
  XNOR2_X1  g244(.A(G2427), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2430), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(KEYINPUT14), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1341), .B(G1348), .Z(new_n676));
  XNOR2_X1  g251(.A(G2443), .B(G2446), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2451), .B(G2454), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n682), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n683), .A2(G14), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(G401));
  INV_X1    g261(.A(KEYINPUT18), .ZN(new_n687));
  XOR2_X1   g262(.A(G2084), .B(G2090), .Z(new_n688));
  XNOR2_X1  g263(.A(G2067), .B(G2678), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT17), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n687), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G2100), .ZN(new_n694));
  XOR2_X1   g269(.A(G2072), .B(G2078), .Z(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n690), .B2(KEYINPUT18), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G2096), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(G227));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(new_n709), .B(new_n708), .S(new_n701), .Z(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(G1991), .B(G1996), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1981), .B(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(G229));
  NOR2_X1   g292(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT91), .ZN(new_n722));
  INV_X1    g297(.A(G1971), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n719), .A2(G23), .ZN(new_n725));
  INV_X1    g300(.A(G288), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT33), .ZN(new_n728));
  INV_X1    g303(.A(G1976), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT34), .ZN(new_n732));
  MUX2_X1   g307(.A(G6), .B(G305), .S(G16), .Z(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT32), .B(G1981), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n731), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n487), .A2(new_n490), .A3(G119), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n742));
  INV_X1    g317(.A(G107), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G2105), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G131), .B2(new_n477), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT35), .B(G1991), .Z(new_n749));
  XOR2_X1   g324(.A(new_n748), .B(new_n749), .Z(new_n750));
  MUX2_X1   g325(.A(G24), .B(G290), .S(G16), .Z(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT88), .B(G1986), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n750), .B(new_n753), .C1(KEYINPUT92), .C2(KEYINPUT36), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n738), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n732), .B1(new_n731), .B2(new_n737), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n718), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n756), .ZN(new_n758));
  INV_X1    g333(.A(new_n718), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n758), .A2(new_n759), .A3(new_n738), .A4(new_n754), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n719), .A2(G4), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n639), .B2(new_n719), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT93), .B(G1348), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n762), .B(new_n763), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n739), .A2(G32), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND3_X1  g342(.A1(new_n478), .A2(G105), .A3(G2104), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n478), .A2(KEYINPUT97), .A3(G105), .A4(G2104), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n477), .A2(G141), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G129), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n767), .B(new_n772), .C1(new_n491), .C2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n765), .B1(new_n775), .B2(new_n739), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT27), .ZN(new_n777));
  INV_X1    g352(.A(G1996), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n548), .A2(new_n719), .ZN(new_n781));
  MUX2_X1   g356(.A(new_n780), .B(KEYINPUT98), .S(new_n781), .Z(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n777), .A2(new_n778), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n764), .A2(new_n779), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n739), .A2(G26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT28), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n487), .A2(new_n490), .A3(G128), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n790));
  INV_X1    g365(.A(G116), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(G2105), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G140), .B2(new_n477), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n794), .A2(KEYINPUT95), .A3(G29), .ZN(new_n795));
  AOI21_X1  g370(.A(KEYINPUT95), .B1(new_n794), .B2(G29), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n788), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(G171), .A2(new_n719), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G5), .B2(new_n719), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(G1961), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(G1961), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n739), .A2(G35), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G162), .B2(new_n739), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT29), .B(G2090), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n803), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(G164), .A2(G29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G27), .B2(G29), .ZN(new_n811));
  INV_X1    g386(.A(G2078), .ZN(new_n812));
  INV_X1    g387(.A(G2072), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n739), .A2(G33), .ZN(new_n814));
  NAND2_X1  g389(.A1(G115), .A2(G2104), .ZN(new_n815));
  INV_X1    g390(.A(G127), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n466), .B2(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n817), .A2(G2105), .B1(G139), .B2(new_n477), .ZN(new_n818));
  NAND2_X1  g393(.A1(G103), .A2(G2104), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT96), .B1(new_n819), .B2(G2105), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n821), .A2(new_n478), .A3(G103), .A4(G2104), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n820), .A2(KEYINPUT25), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT25), .B1(new_n820), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n814), .B1(new_n826), .B2(G29), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n827), .ZN(new_n828));
  OAI221_X1 g403(.A(new_n828), .B1(new_n739), .B2(new_n661), .C1(new_n813), .C2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(G160), .A2(G29), .ZN(new_n830));
  INV_X1    g405(.A(G34), .ZN(new_n831));
  AOI21_X1  g406(.A(G29), .B1(new_n831), .B2(KEYINPUT24), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(KEYINPUT24), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G2084), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n830), .A2(G2084), .A3(new_n833), .ZN(new_n837));
  NOR2_X1   g412(.A1(G16), .A2(G19), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n573), .B2(G16), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT94), .B(G1341), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n836), .B(new_n837), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n811), .A2(new_n812), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  NOR2_X1   g418(.A1(KEYINPUT31), .A2(G11), .ZN(new_n844));
  AND2_X1   g419(.A1(KEYINPUT31), .A2(G11), .ZN(new_n845));
  INV_X1    g420(.A(G28), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT30), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT30), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n739), .B1(new_n848), .B2(G28), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n843), .B1(new_n844), .B2(new_n845), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  NOR4_X1   g425(.A1(new_n829), .A2(new_n841), .A3(new_n842), .A4(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n786), .A2(new_n799), .A3(new_n809), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n719), .A2(G20), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT23), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n644), .B2(new_n719), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G1956), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n757), .A2(new_n760), .A3(new_n857), .ZN(G150));
  INV_X1    g433(.A(G150), .ZN(G311));
  AND2_X1   g434(.A1(G80), .A2(G543), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n519), .B2(G67), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(new_n521), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n526), .A2(G55), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n613), .A2(G93), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n649), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT99), .A4(new_n863), .ZN(new_n870));
  INV_X1    g445(.A(G93), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n863), .B1(new_n871), .B2(new_n530), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n861), .A2(new_n521), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n874), .A3(new_n573), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n639), .A2(G559), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT100), .Z(new_n882));
  INV_X1    g457(.A(G860), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n879), .B2(new_n880), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n867), .B1(new_n882), .B2(new_n884), .ZN(G145));
  NAND2_X1  g460(.A1(new_n661), .A2(G162), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n661), .A2(G162), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n484), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n661), .A2(G162), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(G160), .A3(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n826), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n515), .A2(new_n794), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n504), .A2(new_n789), .A3(new_n514), .A4(new_n793), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n895), .A2(new_n774), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n774), .B1(new_n895), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n896), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n504), .A2(new_n514), .B1(new_n789), .B2(new_n793), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n775), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n774), .A3(new_n896), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n818), .A2(new_n825), .A3(KEYINPUT101), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  INV_X1    g482(.A(G130), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n491), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT103), .A4(G130), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  INV_X1    g487(.A(G118), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(G2105), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n477), .A2(G142), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT102), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n477), .A2(new_n917), .A3(G142), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n911), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n746), .A2(new_n665), .ZN(new_n921));
  INV_X1    g496(.A(new_n665), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(new_n741), .A3(new_n745), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n911), .A2(new_n921), .A3(new_n919), .A4(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n899), .A2(new_n906), .A3(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n892), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n899), .A2(new_n906), .ZN(new_n930));
  INV_X1    g505(.A(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(KEYINPUT104), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n932), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(KEYINPUT104), .A3(new_n931), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n892), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n934), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g515(.A(KEYINPUT105), .B(new_n892), .C1(new_n936), .C2(new_n937), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n933), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT106), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(new_n933), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n943), .A2(KEYINPUT40), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT40), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(G395));
  XNOR2_X1  g523(.A(new_n876), .B(new_n651), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n638), .B1(new_n601), .B2(new_n603), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n588), .B1(new_n519), .B2(G65), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n521), .B1(new_n951), .B2(KEYINPUT76), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n590), .B1(new_n952), .B2(new_n589), .ZN(new_n953));
  INV_X1    g528(.A(new_n591), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n600), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n602), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n592), .A2(KEYINPUT78), .A3(new_n600), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(new_n957), .A3(new_n639), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n950), .A2(new_n958), .A3(KEYINPUT41), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT41), .B1(new_n950), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n949), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(KEYINPUT107), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n950), .A2(new_n958), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n961), .B(KEYINPUT107), .C1(new_n964), .C2(new_n949), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n965), .A3(KEYINPUT108), .ZN(new_n967));
  XOR2_X1   g542(.A(G290), .B(G305), .Z(new_n968));
  XNOR2_X1  g543(.A(new_n726), .B(G303), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT42), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n966), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n962), .A2(new_n965), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(new_n971), .ZN(new_n975));
  OAI21_X1  g550(.A(G868), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n865), .A2(new_n642), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(G295));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n977), .ZN(G331));
  NAND2_X1  g554(.A1(new_n561), .A2(new_n562), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT74), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n611), .A2(new_n983), .A3(new_n560), .ZN(new_n984));
  NAND2_X1  g559(.A1(G301), .A2(new_n548), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n984), .B2(new_n985), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n876), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n985), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT110), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n869), .A2(new_n875), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n964), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n994), .A2(KEYINPUT111), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n959), .A2(new_n960), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G37), .B1(new_n1002), .B2(new_n970), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n995), .B1(new_n959), .B2(new_n960), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n995), .B(KEYINPUT112), .C1(new_n959), .C2(new_n960), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n998), .A2(new_n963), .A3(new_n999), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n970), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1003), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n989), .B2(new_n994), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n994), .A2(KEYINPUT111), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1014), .A2(new_n1015), .B1(new_n960), .B2(new_n959), .ZN(new_n1016));
  INV_X1    g591(.A(new_n996), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n970), .ZN(new_n1018));
  INV_X1    g593(.A(G37), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n970), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT43), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT43), .B1(new_n1026), .B2(new_n1020), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1003), .B(new_n1012), .C1(new_n970), .C2(new_n1002), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(KEYINPUT44), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1029), .ZN(G397));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n501), .A2(new_n503), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n507), .A2(new_n512), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n513), .A2(G126), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n504), .B2(new_n514), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n472), .A2(G40), .A3(new_n483), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n746), .B(new_n749), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT114), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n794), .B(new_n798), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n774), .B(new_n778), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(G290), .B(G1986), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1044), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1036), .A2(KEYINPUT116), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1043), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1039), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n726), .A2(G1976), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(G8), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT52), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n623), .A2(G651), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n526), .A2(G48), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(G1981), .B1(new_n1062), .B2(new_n619), .ZN(new_n1063));
  INV_X1    g638(.A(G1981), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n620), .A2(new_n624), .A3(new_n1064), .A4(new_n626), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1065), .A3(KEYINPUT49), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n1056), .A3(G8), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1059), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n729), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1056), .A2(G8), .A3(new_n1057), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n515), .A2(KEYINPUT45), .A3(new_n1031), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1053), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1039), .A2(KEYINPUT45), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n723), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT50), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n515), .A2(new_n1082), .A3(new_n1031), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1039), .A2(KEYINPUT120), .A3(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1054), .B1(new_n515), .B2(new_n1031), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT116), .B(G1384), .C1(new_n504), .C2(new_n514), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT50), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1090), .A3(new_n1053), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1081), .B1(new_n1091), .B2(G2090), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G303), .A2(G8), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1081), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1052), .A2(new_n1082), .A3(new_n1055), .ZN(new_n1101));
  INV_X1    g676(.A(G2090), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1036), .A2(KEYINPUT50), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1053), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1043), .B1(new_n1039), .B2(KEYINPUT45), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(KEYINPUT45), .B2(new_n1039), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(KEYINPUT115), .A3(new_n723), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(new_n1104), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(G8), .A3(new_n1096), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT121), .B(G2084), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1043), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1101), .A2(new_n1103), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1038), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1966), .B1(new_n1113), .B2(new_n1105), .ZN(new_n1114));
  OAI211_X1 g689(.A(G8), .B(new_n611), .C1(new_n1112), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1077), .A2(new_n1098), .A3(new_n1109), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1108), .A2(G8), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1097), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1076), .A2(new_n1075), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1059), .A2(new_n1070), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1109), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1120), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1096), .B1(new_n1108), .B2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT45), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n783), .B1(new_n1130), .B2(new_n1079), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1101), .A2(new_n1103), .A3(new_n1111), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(KEYINPUT63), .A3(G8), .A4(new_n611), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(KEYINPUT122), .A3(new_n1109), .A4(new_n1077), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1119), .A2(new_n1128), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1070), .A2(new_n729), .A3(new_n726), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1065), .ZN(new_n1139));
  OAI211_X1 g714(.A(G8), .B(new_n1056), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1075), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1126), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1143), .B2(new_n1109), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT119), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1140), .B(new_n1146), .C1(new_n1143), .C2(new_n1109), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(KEYINPUT51), .ZN(new_n1150));
  INV_X1    g725(.A(G8), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1152));
  NOR2_X1   g727(.A1(G168), .A2(new_n1151), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1149), .B2(KEYINPUT51), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1150), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(G8), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1150), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1133), .A2(new_n1153), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT62), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1077), .A2(new_n1098), .A3(new_n1109), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1113), .A2(new_n812), .A3(new_n1105), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT124), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1113), .A2(new_n1166), .A3(new_n812), .A4(new_n1105), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(KEYINPUT53), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1101), .A2(new_n1053), .A3(new_n1103), .ZN(new_n1169));
  XOR2_X1   g744(.A(KEYINPUT125), .B(G1961), .Z(new_n1170));
  INV_X1    g745(.A(KEYINPUT53), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1105), .B(new_n812), .C1(KEYINPUT45), .C2(new_n1039), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1169), .A2(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(G301), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1156), .A2(new_n1159), .A3(new_n1175), .A4(new_n1160), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1162), .A2(new_n1163), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1137), .A2(new_n1148), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(G1956), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1091), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT57), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n955), .B(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT56), .B(G2072), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1180), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1056), .A2(G2067), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n763), .B2(new_n1169), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1188), .A2(new_n638), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1182), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1043), .B1(new_n1191), .B2(KEYINPUT50), .ZN(new_n1192));
  AOI21_X1  g767(.A(G1956), .B1(new_n1192), .B2(new_n1087), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1185), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1190), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1186), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1182), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1186), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1180), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1200));
  AOI21_X1  g775(.A(KEYINPUT61), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1169), .A2(new_n763), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1187), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1203), .A2(new_n1204), .A3(KEYINPUT60), .A4(new_n638), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT59), .ZN(new_n1206));
  XOR2_X1   g781(.A(KEYINPUT58), .B(G1341), .Z(new_n1207));
  AOI22_X1  g782(.A1(new_n1183), .A2(new_n778), .B1(new_n1056), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1208), .B2(new_n649), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n1056), .A2(new_n1207), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1106), .A2(G1996), .ZN(new_n1211));
  OAI211_X1 g786(.A(KEYINPUT59), .B(new_n573), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1205), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1188), .A2(KEYINPUT60), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n638), .B1(new_n1188), .B2(KEYINPUT60), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1213), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1196), .B1(new_n1202), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT54), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1171), .A2(G2078), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1105), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1219), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  NAND4_X1  g798(.A1(new_n1042), .A2(KEYINPUT126), .A3(new_n1105), .A4(new_n1221), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AND3_X1   g800(.A1(new_n1225), .A2(new_n1173), .A3(G301), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1218), .B1(new_n1174), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1168), .A2(G301), .A3(new_n1173), .ZN(new_n1228));
  AND2_X1   g803(.A1(new_n1225), .A2(new_n1173), .ZN(new_n1229));
  OAI211_X1 g804(.A(new_n1228), .B(KEYINPUT54), .C1(new_n1229), .C2(G301), .ZN(new_n1230));
  NAND4_X1  g805(.A1(new_n1163), .A2(new_n1227), .A3(new_n1230), .A4(new_n1161), .ZN(new_n1231));
  NOR2_X1   g806(.A1(new_n1217), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1051), .B1(new_n1178), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1049), .A2(new_n1044), .ZN(new_n1234));
  NOR2_X1   g809(.A1(G290), .A2(G1986), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1044), .A2(new_n1235), .ZN(new_n1236));
  XOR2_X1   g811(.A(new_n1236), .B(KEYINPUT127), .Z(new_n1237));
  OAI21_X1  g812(.A(new_n1234), .B1(new_n1237), .B2(KEYINPUT48), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1238), .B1(KEYINPUT48), .B2(new_n1237), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1044), .A2(new_n778), .ZN(new_n1240));
  OR2_X1    g815(.A1(new_n1240), .A2(KEYINPUT46), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1240), .A2(KEYINPUT46), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1047), .A2(new_n775), .ZN(new_n1243));
  AOI22_X1  g818(.A1(new_n1241), .A2(new_n1242), .B1(new_n1044), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g819(.A(new_n1244), .B(KEYINPUT47), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1048), .A2(new_n1047), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n747), .A2(new_n749), .ZN(new_n1247));
  OAI22_X1  g822(.A1(new_n1246), .A2(new_n1247), .B1(G2067), .B2(new_n794), .ZN(new_n1248));
  AND2_X1   g823(.A1(new_n1248), .A2(new_n1044), .ZN(new_n1249));
  NOR3_X1   g824(.A1(new_n1239), .A2(new_n1245), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1233), .A2(new_n1250), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g826(.A1(new_n943), .A2(new_n945), .ZN(new_n1253));
  NOR4_X1   g827(.A1(G229), .A2(new_n462), .A3(new_n685), .A4(G227), .ZN(new_n1254));
  AND3_X1   g828(.A1(new_n1023), .A2(new_n1253), .A3(new_n1254), .ZN(G308));
  NAND3_X1  g829(.A1(new_n1023), .A2(new_n1253), .A3(new_n1254), .ZN(G225));
endmodule


