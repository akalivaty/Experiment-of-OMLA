

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n728), .A2(n752), .ZN(n730) );
  XOR2_X1 U556 ( .A(n719), .B(n718), .Z(n523) );
  OR2_X1 U557 ( .A1(n732), .A2(G301), .ZN(n524) );
  XOR2_X1 U558 ( .A(n735), .B(KEYINPUT31), .Z(n525) );
  INV_X1 U559 ( .A(KEYINPUT30), .ZN(n729) );
  XNOR2_X1 U560 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U561 ( .A1(n523), .A2(n524), .ZN(n736) );
  NOR2_X1 U562 ( .A1(n739), .A2(G2084), .ZN(n725) );
  NAND2_X1 U563 ( .A1(n736), .A2(n525), .ZN(n750) );
  AND2_X1 U564 ( .A1(n746), .A2(n745), .ZN(n748) );
  INV_X1 U565 ( .A(KEYINPUT105), .ZN(n758) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n784) );
  XNOR2_X1 U567 ( .A(KEYINPUT65), .B(G2104), .ZN(n529) );
  NOR2_X2 U568 ( .A1(G2105), .A2(n529), .ZN(n897) );
  NOR2_X1 U569 ( .A1(n541), .A2(n540), .ZN(G160) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XOR2_X1 U571 ( .A(KEYINPUT17), .B(n526), .Z(n896) );
  NAND2_X1 U572 ( .A1(G138), .A2(n896), .ZN(n528) );
  NAND2_X1 U573 ( .A1(G102), .A2(n897), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n534) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NAND2_X1 U576 ( .A1(G114), .A2(n892), .ZN(n532) );
  NAND2_X1 U577 ( .A1(n529), .A2(G2105), .ZN(n530) );
  XOR2_X2 U578 ( .A(KEYINPUT66), .B(n530), .Z(n893) );
  NAND2_X1 U579 ( .A1(G126), .A2(n893), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U581 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U582 ( .A1(n892), .A2(G113), .ZN(n536) );
  NAND2_X1 U583 ( .A1(n896), .A2(G137), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U585 ( .A1(G125), .A2(n893), .ZN(n539) );
  NAND2_X1 U586 ( .A1(G101), .A2(n897), .ZN(n537) );
  XOR2_X1 U587 ( .A(KEYINPUT23), .B(n537), .Z(n538) );
  NAND2_X1 U588 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U589 ( .A(G2443), .B(G2446), .Z(n543) );
  XNOR2_X1 U590 ( .A(G2427), .B(G2451), .ZN(n542) );
  XNOR2_X1 U591 ( .A(n543), .B(n542), .ZN(n549) );
  XOR2_X1 U592 ( .A(G2430), .B(G2454), .Z(n545) );
  XNOR2_X1 U593 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U594 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U595 ( .A(G2435), .B(G2438), .Z(n546) );
  XNOR2_X1 U596 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U597 ( .A(n549), .B(n548), .Z(n550) );
  AND2_X1 U598 ( .A1(G14), .A2(n550), .ZN(G401) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U600 ( .A(G57), .ZN(G237) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U603 ( .A(G651), .B(KEYINPUT67), .ZN(n553) );
  NOR2_X1 U604 ( .A1(G543), .A2(n553), .ZN(n551) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n551), .Z(n663) );
  NAND2_X1 U606 ( .A1(n663), .A2(G64), .ZN(n552) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(n552), .ZN(n562) );
  XNOR2_X1 U608 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n557) );
  XOR2_X1 U609 ( .A(KEYINPUT0), .B(G543), .Z(n651) );
  NOR2_X1 U610 ( .A1(n651), .A2(n553), .ZN(n657) );
  NAND2_X1 U611 ( .A1(G77), .A2(n657), .ZN(n555) );
  NOR2_X1 U612 ( .A1(G651), .A2(G543), .ZN(n658) );
  NAND2_X1 U613 ( .A1(G90), .A2(n658), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n557), .B(n556), .ZN(n560) );
  NOR2_X1 U616 ( .A1(G651), .A2(n651), .ZN(n558) );
  XNOR2_X1 U617 ( .A(KEYINPUT64), .B(n558), .ZN(n662) );
  NAND2_X1 U618 ( .A1(G52), .A2(n662), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U620 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U621 ( .A1(G89), .A2(n658), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT4), .B(n563), .Z(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT75), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G76), .A2(n657), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G63), .A2(n663), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G51), .A2(n662), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U632 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U635 ( .A(n574), .B(KEYINPUT10), .ZN(n575) );
  XNOR2_X1 U636 ( .A(KEYINPUT72), .B(n575), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n839) );
  NAND2_X1 U638 ( .A1(n839), .A2(G567), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n663), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n577), .Z(n585) );
  NAND2_X1 U642 ( .A1(n657), .A2(G68), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT74), .B(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT73), .B(KEYINPUT12), .Z(n580) );
  NAND2_X1 U645 ( .A1(G81), .A2(n658), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n583), .Z(n584) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G43), .A2(n662), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n959) );
  INV_X1 U652 ( .A(G860), .ZN(n627) );
  OR2_X1 U653 ( .A1(n959), .A2(n627), .ZN(G153) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U656 ( .A1(G79), .A2(n657), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G66), .A2(n663), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U659 ( .A1(G92), .A2(n658), .ZN(n591) );
  NAND2_X1 U660 ( .A1(G54), .A2(n662), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n594), .Z(n953) );
  OR2_X1 U664 ( .A1(n953), .A2(G868), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G65), .A2(n663), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G53), .A2(n662), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G78), .A2(n657), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G91), .A2(n658), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n954) );
  XNOR2_X1 U673 ( .A(n954), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U674 ( .A1(G286), .A2(G868), .ZN(n605) );
  INV_X1 U675 ( .A(G868), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G299), .A2(n603), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n627), .A2(G559), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n606), .A2(n953), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT16), .ZN(n608) );
  XNOR2_X1 U681 ( .A(KEYINPUT76), .B(n608), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n959), .ZN(n609) );
  XOR2_X1 U683 ( .A(KEYINPUT77), .B(n609), .Z(n612) );
  NAND2_X1 U684 ( .A1(G868), .A2(n953), .ZN(n610) );
  NOR2_X1 U685 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U687 ( .A(KEYINPUT78), .B(n613), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G123), .A2(n893), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G135), .A2(n896), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT79), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G111), .A2(n892), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n897), .A2(G99), .ZN(n620) );
  XOR2_X1 U696 ( .A(KEYINPUT80), .B(n620), .Z(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n1011) );
  XNOR2_X1 U698 ( .A(n1011), .B(G2096), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT81), .ZN(n624) );
  NOR2_X1 U700 ( .A1(G2100), .A2(n624), .ZN(n625) );
  XOR2_X1 U701 ( .A(KEYINPUT82), .B(n625), .Z(G156) );
  NAND2_X1 U702 ( .A1(G559), .A2(n953), .ZN(n626) );
  XOR2_X1 U703 ( .A(n959), .B(n626), .Z(n673) );
  NAND2_X1 U704 ( .A1(n627), .A2(n673), .ZN(n634) );
  NAND2_X1 U705 ( .A1(G67), .A2(n663), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G55), .A2(n662), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G80), .A2(n657), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G93), .A2(n658), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n675) );
  XOR2_X1 U712 ( .A(n634), .B(n675), .Z(G145) );
  NAND2_X1 U713 ( .A1(n662), .A2(G50), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G75), .A2(n657), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G88), .A2(n658), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n663), .A2(G62), .ZN(n637) );
  XOR2_X1 U718 ( .A(KEYINPUT84), .B(n637), .Z(n638) );
  NOR2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(KEYINPUT85), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G86), .A2(n658), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G48), .A2(n662), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U725 ( .A1(G73), .A2(n657), .ZN(n645) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n645), .Z(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n663), .A2(G61), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U730 ( .A(KEYINPUT83), .B(n650), .Z(G305) );
  NAND2_X1 U731 ( .A1(G87), .A2(n651), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U734 ( .A1(n663), .A2(n654), .ZN(n656) );
  NAND2_X1 U735 ( .A1(G49), .A2(n662), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(G288) );
  NAND2_X1 U737 ( .A1(G72), .A2(n657), .ZN(n660) );
  NAND2_X1 U738 ( .A1(G85), .A2(n658), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U740 ( .A(KEYINPUT68), .B(n661), .Z(n667) );
  NAND2_X1 U741 ( .A1(n662), .A2(G47), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G60), .A2(n663), .ZN(n664) );
  AND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n667), .A2(n666), .ZN(G290) );
  XNOR2_X1 U745 ( .A(G166), .B(G299), .ZN(n672) );
  XNOR2_X1 U746 ( .A(KEYINPUT19), .B(G305), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n668), .B(G288), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n675), .B(n669), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n670), .B(G290), .ZN(n671) );
  XNOR2_X1 U750 ( .A(n672), .B(n671), .ZN(n911) );
  XNOR2_X1 U751 ( .A(n673), .B(n911), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n674), .A2(G868), .ZN(n677) );
  OR2_X1 U753 ( .A1(G868), .A2(n675), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n678) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n679), .ZN(n681) );
  XNOR2_X1 U758 ( .A(KEYINPUT86), .B(KEYINPUT21), .ZN(n680) );
  XNOR2_X1 U759 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U760 ( .A1(n682), .A2(G2072), .ZN(n683) );
  XOR2_X1 U761 ( .A(KEYINPUT87), .B(n683), .Z(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U765 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U766 ( .A1(G96), .A2(n686), .ZN(n845) );
  NAND2_X1 U767 ( .A1(n845), .A2(G2106), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G69), .A2(G120), .ZN(n687) );
  NOR2_X1 U769 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U770 ( .A1(G108), .A2(n688), .ZN(n844) );
  NAND2_X1 U771 ( .A1(n844), .A2(G567), .ZN(n689) );
  NAND2_X1 U772 ( .A1(n690), .A2(n689), .ZN(n847) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U774 ( .A1(n847), .A2(n691), .ZN(n841) );
  NAND2_X1 U775 ( .A1(n841), .A2(G36), .ZN(G176) );
  XOR2_X1 U776 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  NOR2_X1 U777 ( .A1(G303), .A2(G1971), .ZN(n692) );
  NOR2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n947) );
  NOR2_X1 U779 ( .A1(n692), .A2(n947), .ZN(n757) );
  NAND2_X1 U780 ( .A1(G160), .A2(G40), .ZN(n783) );
  INV_X1 U781 ( .A(n783), .ZN(n699) );
  AND2_X1 U782 ( .A1(n784), .A2(G1996), .ZN(n693) );
  AND2_X1 U783 ( .A1(n699), .A2(n693), .ZN(n694) );
  XOR2_X1 U784 ( .A(n694), .B(KEYINPUT26), .Z(n697) );
  NAND2_X2 U785 ( .A1(n699), .A2(n784), .ZN(n739) );
  AND2_X1 U786 ( .A1(n739), .A2(G1341), .ZN(n695) );
  NOR2_X1 U787 ( .A1(n695), .A2(n959), .ZN(n696) );
  AND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n708) );
  NOR2_X1 U789 ( .A1(n708), .A2(n953), .ZN(n704) );
  AND2_X1 U790 ( .A1(G1348), .A2(n739), .ZN(n698) );
  XNOR2_X1 U791 ( .A(n698), .B(KEYINPUT99), .ZN(n701) );
  AND2_X1 U792 ( .A1(n699), .A2(n784), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n720), .A2(G2067), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U795 ( .A(n702), .B(KEYINPUT100), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n712) );
  NAND2_X1 U797 ( .A1(n720), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  AND2_X1 U799 ( .A1(G1956), .A2(n739), .ZN(n706) );
  NOR2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n714) );
  NAND2_X1 U801 ( .A1(n714), .A2(n954), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n708), .A2(n953), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U805 ( .A(n713), .B(KEYINPUT101), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n954), .A2(n714), .ZN(n715) );
  XOR2_X1 U807 ( .A(KEYINPUT28), .B(n715), .Z(n716) );
  NAND2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U809 ( .A(KEYINPUT102), .B(KEYINPUT29), .ZN(n718) );
  NOR2_X1 U810 ( .A1(n720), .A2(G1961), .ZN(n721) );
  XNOR2_X1 U811 ( .A(n721), .B(KEYINPUT98), .ZN(n723) );
  XOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .Z(n926) );
  NOR2_X1 U813 ( .A1(n739), .A2(n926), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n732) );
  INV_X1 U815 ( .A(KEYINPUT97), .ZN(n724) );
  XNOR2_X1 U816 ( .A(n725), .B(n724), .ZN(n749) );
  INV_X1 U817 ( .A(n749), .ZN(n726) );
  NAND2_X1 U818 ( .A1(G8), .A2(n726), .ZN(n728) );
  NAND2_X1 U819 ( .A1(n739), .A2(G8), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(KEYINPUT94), .ZN(n827) );
  NOR2_X1 U821 ( .A1(n827), .A2(G1966), .ZN(n752) );
  NOR2_X1 U822 ( .A1(G168), .A2(n731), .ZN(n734) );
  AND2_X1 U823 ( .A1(G301), .A2(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n750), .A2(n737), .ZN(n746) );
  INV_X1 U827 ( .A(G8), .ZN(n744) );
  NOR2_X1 U828 ( .A1(n827), .A2(G1971), .ZN(n738) );
  XOR2_X1 U829 ( .A(KEYINPUT103), .B(n738), .Z(n741) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(G303), .A2(n742), .ZN(n743) );
  OR2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U834 ( .A(KEYINPUT104), .B(KEYINPUT32), .ZN(n747) );
  XNOR2_X1 U835 ( .A(n748), .B(n747), .ZN(n756) );
  NAND2_X1 U836 ( .A1(n749), .A2(G8), .ZN(n754) );
  INV_X1 U837 ( .A(n750), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n756), .A2(n755), .ZN(n821) );
  NAND2_X1 U841 ( .A1(n757), .A2(n821), .ZN(n759) );
  XNOR2_X1 U842 ( .A(n759), .B(n758), .ZN(n760) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n948) );
  NAND2_X1 U844 ( .A1(n760), .A2(n948), .ZN(n761) );
  XNOR2_X1 U845 ( .A(KEYINPUT106), .B(n761), .ZN(n763) );
  OR2_X1 U846 ( .A1(n827), .A2(KEYINPUT107), .ZN(n762) );
  NOR2_X1 U847 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n764), .ZN(n771) );
  INV_X1 U849 ( .A(KEYINPUT107), .ZN(n766) );
  NAND2_X1 U850 ( .A1(n947), .A2(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n947), .A2(KEYINPUT107), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U854 ( .A1(n827), .A2(n769), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n807) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n944) );
  XNOR2_X1 U857 ( .A(G2067), .B(KEYINPUT37), .ZN(n815) );
  NAND2_X1 U858 ( .A1(n896), .A2(G140), .ZN(n772) );
  XNOR2_X1 U859 ( .A(n772), .B(KEYINPUT90), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G104), .A2(n897), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n776) );
  XOR2_X1 U862 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n775) );
  XNOR2_X1 U863 ( .A(n776), .B(n775), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G116), .A2(n892), .ZN(n778) );
  NAND2_X1 U865 ( .A1(G128), .A2(n893), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT35), .B(n779), .Z(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(KEYINPUT36), .B(n782), .ZN(n889) );
  NOR2_X1 U870 ( .A1(n815), .A2(n889), .ZN(n1014) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n818) );
  NAND2_X1 U872 ( .A1(n1014), .A2(n818), .ZN(n813) );
  XNOR2_X1 U873 ( .A(G1986), .B(G290), .ZN(n956) );
  NAND2_X1 U874 ( .A1(n956), .A2(n818), .ZN(n785) );
  XOR2_X1 U875 ( .A(KEYINPUT89), .B(n785), .Z(n786) );
  NAND2_X1 U876 ( .A1(n813), .A2(n786), .ZN(n831) );
  INV_X1 U877 ( .A(n831), .ZN(n787) );
  AND2_X1 U878 ( .A1(n944), .A2(n787), .ZN(n805) );
  NAND2_X1 U879 ( .A1(n897), .A2(G95), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G119), .A2(n893), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G131), .A2(n896), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G107), .A2(n892), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n877) );
  NAND2_X1 U886 ( .A1(G1991), .A2(n877), .ZN(n794) );
  XNOR2_X1 U887 ( .A(n794), .B(KEYINPUT92), .ZN(n804) );
  NAND2_X1 U888 ( .A1(G105), .A2(n897), .ZN(n795) );
  XNOR2_X1 U889 ( .A(n795), .B(KEYINPUT38), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G117), .A2(n892), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G129), .A2(n893), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U893 ( .A1(G141), .A2(n896), .ZN(n798) );
  XNOR2_X1 U894 ( .A(KEYINPUT93), .B(n798), .ZN(n799) );
  NOR2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n903) );
  NAND2_X1 U897 ( .A1(G1996), .A2(n903), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n1010) );
  NAND2_X1 U899 ( .A1(n818), .A2(n1010), .ZN(n808) );
  AND2_X1 U900 ( .A1(n805), .A2(n808), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n837) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n903), .ZN(n1004) );
  INV_X1 U903 ( .A(n808), .ZN(n833) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n877), .ZN(n1009) );
  NOR2_X1 U906 ( .A1(n809), .A2(n1009), .ZN(n810) );
  NOR2_X1 U907 ( .A1(n833), .A2(n810), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n1004), .A2(n811), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n815), .A2(n889), .ZN(n1018) );
  NAND2_X1 U912 ( .A1(n816), .A2(n1018), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n835) );
  NOR2_X1 U914 ( .A1(G2090), .A2(G303), .ZN(n819) );
  NAND2_X1 U915 ( .A1(G8), .A2(n819), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n827), .A2(n822), .ZN(n829) );
  NOR2_X1 U918 ( .A1(G1981), .A2(G305), .ZN(n825) );
  XOR2_X1 U919 ( .A(KEYINPUT24), .B(KEYINPUT96), .Z(n823) );
  XNOR2_X1 U920 ( .A(KEYINPUT95), .B(n823), .ZN(n824) );
  XOR2_X1 U921 ( .A(n825), .B(n824), .Z(n826) );
  OR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  AND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  OR2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  OR2_X1 U925 ( .A1(n833), .A2(n832), .ZN(n834) );
  AND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U928 ( .A(n838), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n839), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U931 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G1), .A2(G3), .ZN(n842) );
  NAND2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U934 ( .A(n843), .B(KEYINPUT108), .ZN(G188) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U940 ( .A(n846), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U941 ( .A(G261), .ZN(G325) );
  INV_X1 U942 ( .A(n847), .ZN(G319) );
  XOR2_X1 U943 ( .A(G2678), .B(G2096), .Z(n849) );
  XNOR2_X1 U944 ( .A(KEYINPUT110), .B(G2100), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U946 ( .A(n850), .B(KEYINPUT43), .Z(n852) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(KEYINPUT111), .Z(n854) );
  XNOR2_X1 U950 ( .A(G2090), .B(KEYINPUT112), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U952 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(G227) );
  XOR2_X1 U955 ( .A(G1966), .B(G1956), .Z(n860) );
  XNOR2_X1 U956 ( .A(G1971), .B(G1961), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U958 ( .A(n861), .B(KEYINPUT41), .Z(n863) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U961 ( .A(G2474), .B(G1986), .Z(n865) );
  XNOR2_X1 U962 ( .A(G1981), .B(G1976), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G112), .A2(n892), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G100), .A2(n897), .ZN(n868) );
  NAND2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U968 ( .A1(G136), .A2(n896), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n870), .B(KEYINPUT114), .ZN(n874) );
  XOR2_X1 U970 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n872) );
  NAND2_X1 U971 ( .A1(G124), .A2(n893), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U974 ( .A1(n876), .A2(n875), .ZN(G162) );
  XNOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n877), .B(KEYINPUT115), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(G162), .B(n880), .ZN(n891) );
  NAND2_X1 U979 ( .A1(G139), .A2(n896), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G103), .A2(n897), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G115), .A2(n892), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G127), .A2(n893), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT116), .B(n888), .Z(n998) );
  XNOR2_X1 U988 ( .A(n889), .B(n998), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n906) );
  NAND2_X1 U990 ( .A1(G118), .A2(n892), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U993 ( .A1(G142), .A2(n896), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G106), .A2(n897), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(n900), .B(KEYINPUT45), .Z(n901) );
  NOR2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U999 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U1000 ( .A(G160), .B(G164), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1002 ( .A(n1011), .B(n909), .Z(n910) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(G171), .B(n953), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1006 ( .A(n959), .B(G286), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(n918), .B(KEYINPUT118), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n921), .ZN(n922) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n922), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1019 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n1028) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n1022) );
  XNOR2_X1 U1021 ( .A(G2090), .B(G35), .ZN(n935) );
  XOR2_X1 U1022 ( .A(G1991), .B(G25), .Z(n923) );
  NAND2_X1 U1023 ( .A1(n923), .A2(G28), .ZN(n932) );
  XNOR2_X1 U1024 ( .A(G1996), .B(G32), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G33), .B(G2072), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n926), .B(G27), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(G2067), .B(G26), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT53), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1034 ( .A(G2084), .B(G34), .Z(n936) );
  XNOR2_X1 U1035 ( .A(KEYINPUT54), .B(n936), .ZN(n937) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(n1022), .B(n939), .ZN(n941) );
  INV_X1 U1038 ( .A(G29), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(G11), .A2(n942), .ZN(n997) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .ZN(n969) );
  XOR2_X1 U1042 ( .A(G168), .B(G1966), .Z(n943) );
  XNOR2_X1 U1043 ( .A(KEYINPUT121), .B(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(n946), .B(KEYINPUT57), .ZN(n967) );
  INV_X1 U1046 ( .A(n947), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(n950), .B(KEYINPUT122), .ZN(n952) );
  XOR2_X1 U1049 ( .A(G1961), .B(G171), .Z(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(n953), .B(G1348), .ZN(n958) );
  XOR2_X1 U1052 ( .A(n954), .B(G1956), .Z(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G1341), .B(n959), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G303), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n995) );
  INV_X1 U1062 ( .A(G16), .ZN(n993) );
  XOR2_X1 U1063 ( .A(G1986), .B(G24), .Z(n971) );
  XOR2_X1 U1064 ( .A(G1971), .B(G22), .Z(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(G23), .B(G1976), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1068 ( .A(KEYINPUT58), .B(n974), .Z(n990) );
  XOR2_X1 U1069 ( .A(G1961), .B(G5), .Z(n985) );
  XNOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(n975), .B(G4), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(G1956), .B(G20), .ZN(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1076 ( .A(KEYINPUT123), .B(G1341), .Z(n980) );
  XNOR2_X1 U1077 ( .A(G19), .B(n980), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT60), .B(n983), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(G21), .B(G1966), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1083 ( .A(KEYINPUT124), .B(n988), .Z(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(KEYINPUT61), .B(n991), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1026) );
  XNOR2_X1 U1089 ( .A(G2072), .B(n998), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(n999), .B(KEYINPUT120), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(G2078), .B(G164), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1002), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT51), .B(n1005), .Z(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1020) );
  XOR2_X1 U1098 ( .A(G2084), .B(G160), .Z(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT119), .B(n1016), .Z(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(n1028), .B(n1027), .ZN(n1029) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1029), .ZN(G150) );
  INV_X1 U1112 ( .A(G150), .ZN(G311) );
endmodule

