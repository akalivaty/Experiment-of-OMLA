//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n187), .A2(KEYINPUT67), .A3(G119), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n194));
  INV_X1    g008(.A(new_n188), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n194), .B(G113), .C1(KEYINPUT5), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G107), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n200), .A2(KEYINPUT3), .A3(G104), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT3), .B1(new_n200), .B2(G104), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n197), .B(new_n199), .C1(new_n201), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n199), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n198), .A2(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n208));
  INV_X1    g022(.A(G113), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT2), .A3(G113), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n210), .A2(new_n212), .B1(new_n208), .B2(new_n209), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT68), .A3(new_n193), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT68), .B1(new_n213), .B2(new_n193), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n196), .B(new_n207), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n198), .B2(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n200), .A2(KEYINPUT3), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n197), .B1(new_n222), .B2(new_n199), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT77), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT4), .A4(new_n203), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n213), .A2(new_n193), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n213), .A2(new_n193), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n232), .B1(new_n235), .B2(new_n214), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n217), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT79), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(KEYINPUT79), .B(new_n217), .C1(new_n231), .C2(new_n236), .ZN(new_n240));
  XOR2_X1   g054(.A(G110), .B(G122), .Z(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT6), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n239), .A2(KEYINPUT6), .A3(new_n240), .A4(new_n241), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n237), .A2(new_n241), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT64), .A2(G143), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT64), .A2(G143), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT64), .A2(G143), .ZN(new_n259));
  OAI21_X1  g073(.A(G146), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n251), .A2(G146), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n260), .A2(G128), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n257), .B1(new_n263), .B2(KEYINPUT0), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n255), .A2(new_n256), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  OAI21_X1  g083(.A(G128), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n260), .A2(new_n269), .A3(G128), .A4(new_n262), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G125), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G224), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n276), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n248), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(KEYINPUT7), .ZN(new_n283));
  OR3_X1    g097(.A1(new_n266), .A2(new_n274), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n285), .B(new_n283), .C1(new_n266), .C2(new_n274), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n276), .A2(new_n283), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT80), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n196), .B1(new_n215), .B2(new_n216), .ZN(new_n290));
  INV_X1    g104(.A(new_n207), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n217), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n241), .B(KEYINPUT8), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n247), .A2(new_n287), .A3(new_n289), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n282), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n300), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n246), .B1(new_n242), .B2(new_n243), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n280), .B1(new_n303), .B2(new_n245), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n304), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G221), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT9), .B(G234), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n309), .B1(new_n311), .B2(new_n297), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  INV_X1    g128(.A(G128), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(new_n255), .B2(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n252), .A2(new_n254), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n261), .B1(new_n317), .B2(G146), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n272), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n207), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT10), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(KEYINPUT78), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n224), .A2(new_n228), .A3(new_n264), .A4(new_n230), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n273), .A2(KEYINPUT10), .A3(new_n207), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G137), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(G137), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(KEYINPUT11), .ZN(new_n333));
  NAND2_X1  g147(.A1(KEYINPUT11), .A2(G134), .ZN(new_n334));
  INV_X1    g148(.A(G137), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT65), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT65), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G137), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G131), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT11), .B1(new_n335), .B2(G134), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n335), .A2(G134), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G131), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n336), .A2(new_n338), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n334), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n326), .A2(new_n329), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n319), .A2(new_n207), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n273), .A2(new_n207), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT12), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT12), .B(new_n347), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G110), .B(G140), .ZN(new_n357));
  INV_X1    g171(.A(G953), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(G227), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n357), .B(new_n359), .Z(new_n360));
  AND3_X1   g174(.A1(new_n349), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT78), .B1(new_n320), .B2(new_n321), .ZN(new_n362));
  AOI211_X1 g176(.A(new_n323), .B(KEYINPUT10), .C1(new_n319), .C2(new_n207), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n327), .A2(new_n328), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n347), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n360), .B1(new_n366), .B2(new_n349), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n314), .B(new_n297), .C1(new_n361), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n349), .A2(new_n356), .ZN(new_n370));
  INV_X1    g184(.A(new_n360), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n349), .A3(new_n360), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(G469), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(G469), .A2(G902), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n313), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n308), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G472), .ZN(new_n379));
  INV_X1    g193(.A(G237), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n358), .A3(G210), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(new_n197), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n382), .B(new_n383), .Z(new_n384));
  AND3_X1   g198(.A1(new_n336), .A2(new_n338), .A3(new_n330), .ZN(new_n385));
  OAI21_X1  g199(.A(G131), .B1(new_n385), .B2(new_n332), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n273), .A2(new_n346), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT69), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n264), .A2(new_n388), .A3(new_n347), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n264), .B2(new_n347), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n236), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n264), .A2(new_n347), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n387), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT30), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n395), .B2(KEYINPUT30), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n384), .B(new_n391), .C1(new_n396), .C2(new_n236), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT31), .ZN(new_n398));
  INV_X1    g212(.A(new_n393), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n387), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(KEYINPUT69), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n264), .A2(new_n347), .A3(new_n388), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n401), .B1(new_n405), .B2(new_n400), .ZN(new_n406));
  INV_X1    g220(.A(new_n236), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT31), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n384), .A4(new_n391), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT28), .B1(new_n399), .B2(new_n236), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n393), .A2(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n391), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT28), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n415), .B2(KEYINPUT70), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT28), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n391), .B2(new_n413), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT70), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n384), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n379), .B(new_n297), .C1(new_n411), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n384), .ZN(new_n425));
  INV_X1    g239(.A(new_n420), .ZN(new_n426));
  INV_X1    g240(.A(new_n412), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n418), .B2(new_n419), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n398), .A3(new_n410), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT32), .A3(new_n379), .A4(new_n297), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n395), .A2(new_n407), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n417), .B1(new_n432), .B2(new_n391), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n412), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT29), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n426), .A2(new_n428), .A3(new_n425), .ZN(new_n438));
  INV_X1    g252(.A(new_n391), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n406), .B2(new_n407), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n435), .B1(new_n440), .B2(new_n384), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n437), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G472), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n424), .A2(new_n431), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n315), .A2(G119), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n315), .A2(G119), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT71), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n315), .A2(KEYINPUT71), .A3(G119), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT24), .B(G110), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT23), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n446), .B1(new_n453), .B2(new_n445), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n190), .A2(G128), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n455), .A2(KEYINPUT72), .A3(KEYINPUT23), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT72), .B1(new_n455), .B2(KEYINPUT23), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n452), .B1(new_n458), .B2(G110), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n265), .A2(G140), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT16), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT74), .ZN(new_n462));
  INV_X1    g276(.A(G140), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(G125), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT74), .B1(new_n265), .B2(G140), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n464), .B1(new_n465), .B2(new_n460), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n461), .B1(new_n466), .B2(KEYINPUT16), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(new_n253), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(G125), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n265), .A2(G140), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n469), .A2(new_n470), .A3(new_n253), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n459), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G110), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(KEYINPUT73), .B2(new_n458), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n467), .A2(new_n253), .ZN(new_n478));
  AOI211_X1 g292(.A(G146), .B(new_n461), .C1(new_n466), .C2(KEYINPUT16), .ZN(new_n479));
  OAI22_X1  g293(.A1(new_n478), .A2(new_n479), .B1(new_n450), .B2(new_n451), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n473), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT75), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n473), .B(KEYINPUT75), .C1(new_n477), .C2(new_n480), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT22), .B(G137), .ZN(new_n485));
  INV_X1    g299(.A(G234), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n309), .A2(new_n486), .A3(G953), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n485), .B(new_n487), .Z(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(new_n482), .A3(new_n488), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G217), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(G234), .B2(new_n297), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(G902), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n492), .A2(KEYINPUT76), .A3(new_n495), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n490), .B2(new_n491), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n494), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI211_X1 g316(.A(KEYINPUT25), .B(G902), .C1(new_n490), .C2(new_n491), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n498), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n198), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT19), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n469), .A2(new_n470), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n466), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n253), .B(new_n511), .C1(new_n512), .C2(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n468), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n258), .A2(new_n259), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n380), .A2(new_n358), .A3(G214), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT81), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT81), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n380), .A2(new_n358), .A3(G214), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n317), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT82), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n516), .A2(new_n521), .A3(G143), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT82), .B1(new_n519), .B2(new_n251), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n517), .A2(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(new_n344), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n344), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n520), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n522), .A2(new_n523), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT18), .A3(G131), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n471), .B1(G146), .B2(new_n466), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT18), .A2(G131), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n509), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n508), .B(KEYINPUT83), .ZN(new_n539));
  INV_X1    g353(.A(new_n527), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n540), .A2(new_n525), .A3(KEYINPUT17), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n478), .A2(new_n479), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n531), .A2(KEYINPUT17), .A3(G131), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n536), .B(new_n539), .C1(new_n541), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G475), .A2(G902), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n506), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n547), .ZN(new_n549));
  AOI211_X1 g363(.A(KEYINPUT20), .B(new_n549), .C1(new_n538), .C2(new_n545), .ZN(new_n550));
  INV_X1    g364(.A(G475), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n536), .B1(new_n541), .B2(new_n544), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n509), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n553), .B2(new_n545), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n548), .A2(new_n550), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n310), .A2(new_n493), .A3(G953), .ZN(new_n557));
  INV_X1    g371(.A(G122), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G116), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n200), .B1(new_n559), .B2(KEYINPUT14), .ZN(new_n560));
  XNOR2_X1  g374(.A(G116), .B(G122), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n317), .A2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n315), .A2(G143), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n563), .A2(new_n330), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n330), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT86), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n562), .B(KEYINPUT86), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT84), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n561), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n200), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n561), .B(KEYINPUT84), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G107), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n563), .A2(new_n330), .A3(new_n564), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n515), .A2(new_n315), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT85), .B1(new_n579), .B2(KEYINPUT13), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT85), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n563), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(KEYINPUT13), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n580), .A2(new_n564), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n578), .B1(G134), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n557), .B1(new_n571), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(G134), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n588), .A2(new_n577), .A3(new_n574), .A4(new_n576), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n569), .A2(new_n570), .ZN(new_n590));
  INV_X1    g404(.A(new_n557), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n587), .A2(new_n297), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT15), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n595), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n587), .A2(new_n297), .A3(new_n592), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n556), .A2(new_n600), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n297), .B(new_n358), .C1(G234), .C2(G237), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT21), .B(G898), .Z(new_n604));
  OR2_X1    g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(KEYINPUT87), .A2(G952), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(KEYINPUT87), .A2(G952), .ZN(new_n608));
  AOI21_X1  g422(.A(G953), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n486), .B2(new_n380), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n601), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n378), .A2(new_n444), .A3(new_n505), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n557), .B2(KEYINPUT89), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT88), .ZN(new_n617));
  INV_X1    g431(.A(new_n592), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n591), .B1(new_n589), .B2(new_n590), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n617), .B1(KEYINPUT88), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n587), .A2(new_n592), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n594), .A2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n593), .A2(new_n594), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n555), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n306), .A2(new_n629), .A3(new_n307), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n611), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n297), .B1(new_n411), .B2(new_n421), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n422), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(new_n504), .A3(new_n377), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  XNOR2_X1  g453(.A(new_n611), .B(KEYINPUT90), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n555), .A2(new_n600), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n306), .A2(new_n641), .A3(new_n307), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  INV_X1    g459(.A(new_n307), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n301), .B2(new_n305), .ZN(new_n647));
  INV_X1    g461(.A(new_n376), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n312), .B1(new_n648), .B2(new_n368), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n481), .B(KEYINPUT91), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n489), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n495), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n653), .B1(new_n503), .B2(new_n502), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n647), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n635), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n613), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT92), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G12));
  AND2_X1   g474(.A1(new_n655), .A2(new_n444), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n556), .A2(new_n599), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n610), .B1(G900), .B2(new_n603), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XNOR2_X1  g481(.A(new_n663), .B(KEYINPUT39), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT40), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n306), .B(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n556), .A2(new_n600), .ZN(new_n674));
  INV_X1    g488(.A(new_n502), .ZN(new_n675));
  INV_X1    g489(.A(new_n503), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n675), .A2(new_n676), .B1(new_n495), .B2(new_n652), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n677), .A3(new_n307), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n670), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n440), .A2(new_n425), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n432), .A2(new_n425), .A3(new_n391), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n297), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n424), .A2(new_n431), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(KEYINPUT94), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(KEYINPUT94), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n679), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n515), .ZN(G45));
  NOR2_X1   g503(.A1(new_n628), .A2(new_n664), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n661), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  OAI21_X1  g506(.A(new_n297), .B1(new_n361), .B2(new_n367), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n313), .A3(new_n368), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT95), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT95), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n694), .A2(new_n697), .A3(new_n313), .A4(new_n368), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n444), .A2(new_n505), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT96), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n632), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT96), .B1(new_n700), .B2(new_n631), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT41), .B(G113), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT97), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n444), .A2(new_n642), .A3(new_n505), .A4(new_n699), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  INV_X1    g524(.A(KEYINPUT99), .ZN(new_n711));
  INV_X1    g525(.A(new_n695), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n647), .A2(new_n712), .A3(KEYINPUT98), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT98), .B1(new_n647), .B2(new_n712), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n677), .A2(new_n601), .A3(new_n612), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n444), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n711), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n715), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(KEYINPUT99), .A3(new_n444), .A4(new_n717), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  OAI21_X1  g538(.A(new_n425), .B1(new_n433), .B2(new_n412), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n398), .A2(new_n410), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(G472), .A2(G902), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n633), .A2(G472), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT100), .B1(new_n728), .B2(new_n505), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n379), .B1(new_n430), .B2(new_n297), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n726), .A2(new_n727), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n504), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n674), .A2(new_n306), .A3(new_n307), .ZN(new_n735));
  INV_X1    g549(.A(new_n640), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n699), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT101), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n735), .A2(new_n736), .A3(new_n699), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n726), .A2(new_n727), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n634), .A2(new_n505), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n732), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n728), .A2(KEYINPUT100), .A3(new_n505), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT101), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n739), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  AND3_X1   g562(.A1(new_n728), .A2(new_n654), .A3(new_n690), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n714), .B2(new_n715), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  NAND3_X1  g565(.A1(new_n301), .A2(new_n305), .A3(new_n307), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n377), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n444), .A2(new_n505), .A3(new_n753), .A4(new_n690), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT102), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n444), .A2(new_n505), .A3(new_n690), .A4(new_n753), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT42), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT102), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n754), .A2(new_n755), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n444), .A2(new_n505), .A3(new_n753), .A4(new_n665), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  AND2_X1   g581(.A1(new_n625), .A2(new_n626), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n555), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT43), .Z(new_n770));
  OR3_X1    g584(.A1(new_n770), .A2(new_n656), .A3(new_n677), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n752), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n372), .A2(new_n373), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n314), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n775), .B2(new_n774), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n375), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n368), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT46), .B1(new_n777), .B2(new_n375), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n313), .B(new_n668), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n773), .B(new_n782), .C1(new_n772), .C2(new_n771), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT103), .B(G137), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT104), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n783), .B(new_n785), .ZN(G39));
  OAI21_X1  g600(.A(new_n313), .B1(new_n779), .B2(new_n780), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n690), .A2(new_n504), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n444), .A2(new_n790), .A3(new_n752), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT106), .B(G140), .Z(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G42));
  NOR3_X1   g608(.A1(new_n734), .A2(new_n610), .A3(new_n770), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n672), .A2(new_n307), .A3(new_n695), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT50), .Z(new_n798));
  NOR2_X1   g612(.A1(new_n752), .A2(new_n695), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT112), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n770), .A2(new_n610), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT113), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(new_n654), .A3(new_n728), .ZN(new_n804));
  INV_X1    g618(.A(new_n752), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n694), .A2(new_n368), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n313), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n805), .B(new_n795), .C1(new_n789), .C2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n798), .A2(new_n804), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n504), .B1(new_n686), .B2(new_n687), .ZN(new_n812));
  INV_X1    g626(.A(new_n610), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n800), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n812), .A2(new_n814), .A3(new_n556), .A4(new_n768), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n811), .A2(new_n816), .B1(KEYINPUT115), .B2(new_n809), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n814), .A3(new_n629), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n795), .A2(new_n721), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n609), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n444), .A2(new_n505), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n803), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT48), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(KEYINPUT48), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n811), .A2(new_n816), .A3(KEYINPUT115), .A4(new_n809), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n655), .B(new_n444), .C1(new_n665), .C2(new_n690), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n377), .A2(new_n654), .A3(new_n664), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n735), .A2(new_n831), .A3(new_n684), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n750), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n750), .A2(new_n830), .A3(new_n835), .A4(new_n832), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(KEYINPUT53), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n614), .A2(new_n657), .A3(new_n709), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n738), .B2(new_n746), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n647), .A2(new_n641), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n630), .A2(new_n736), .B1(new_n841), .B2(KEYINPUT107), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n841), .A2(KEYINPUT107), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n636), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n840), .A2(new_n705), .A3(new_n723), .A4(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n677), .A2(new_n601), .A3(new_n664), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n444), .A3(new_n753), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT108), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n749), .A2(new_n753), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n847), .A2(new_n444), .A3(KEYINPUT108), .A4(new_n753), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n850), .A2(new_n766), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT102), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n838), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n614), .A2(new_n657), .A3(new_n709), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n734), .A2(new_n737), .A3(KEYINPUT101), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n745), .B1(new_n739), .B2(new_n744), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n845), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n853), .B1(new_n758), .B2(new_n763), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n719), .A2(new_n722), .B1(new_n703), .B2(new_n704), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT109), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n837), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n834), .A2(new_n836), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n858), .B2(new_n866), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n829), .A2(new_n867), .B1(new_n869), .B2(KEYINPUT53), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n867), .A2(new_n829), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n756), .A2(new_n757), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n853), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n865), .A3(new_n845), .A4(new_n840), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT111), .B1(new_n875), .B2(new_n837), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n723), .A2(new_n705), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n862), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT111), .ZN(new_n879));
  INV_X1    g693(.A(new_n837), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n874), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n882), .B(new_n883), .C1(KEYINPUT53), .C2(new_n869), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n828), .A2(new_n872), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n769), .A2(new_n307), .A3(new_n313), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n806), .A2(KEYINPUT49), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n806), .A2(KEYINPUT49), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n812), .A2(new_n673), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n358), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n882), .B1(KEYINPUT53), .B2(new_n869), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(G210), .A3(G902), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n248), .A2(new_n281), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n304), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT116), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT55), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(KEYINPUT117), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(KEYINPUT55), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n894), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n898), .B2(new_n906), .ZN(G51));
  NAND2_X1  g722(.A1(new_n858), .A2(new_n866), .ZN(new_n909));
  INV_X1    g723(.A(new_n868), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT53), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n876), .A2(new_n881), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n884), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n911), .A2(new_n912), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n916), .A2(KEYINPUT118), .A3(new_n883), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n375), .B(KEYINPUT57), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n361), .A2(new_n367), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n916), .A2(new_n297), .A3(new_n777), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n893), .B1(new_n921), .B2(new_n922), .ZN(G54));
  NAND4_X1  g737(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  INV_X1    g739(.A(new_n546), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n894), .B1(new_n924), .B2(new_n926), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G60));
  AND2_X1   g744(.A1(new_n620), .A2(new_n623), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT59), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n915), .A2(new_n917), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n872), .B2(new_n884), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n936), .B(new_n894), .C1(new_n937), .C2(new_n931), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT121), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n652), .B(new_n942), .C1(new_n911), .C2(new_n912), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n894), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n492), .B1(new_n895), .B2(new_n942), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT120), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT120), .B(new_n947), .C1(new_n944), .C2(new_n945), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(G66));
  AOI21_X1  g765(.A(new_n358), .B1(new_n604), .B2(G224), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n846), .B2(new_n358), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n303), .B(new_n245), .C1(G898), .C2(new_n358), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(G69));
  OAI21_X1  g769(.A(new_n511), .B1(new_n512), .B2(new_n510), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n406), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n782), .A2(new_n821), .A3(new_n735), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n750), .A2(new_n830), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n766), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n783), .A2(new_n792), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n961), .B2(new_n764), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n358), .A2(G900), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT123), .B1(new_n962), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n957), .A2(new_n358), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n688), .A2(new_n959), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  AOI21_X1  g785(.A(new_n669), .B1(new_n628), .B2(new_n662), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n821), .A2(new_n972), .A3(new_n805), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n783), .A2(new_n792), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n969), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n358), .B1(G227), .B2(G900), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n975), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n968), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n976), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G72));
  NAND3_X1  g797(.A1(new_n961), .A2(new_n764), .A3(new_n878), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT125), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n425), .A3(new_n440), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n894), .ZN(new_n990));
  INV_X1    g804(.A(new_n680), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n971), .A2(new_n878), .A3(new_n974), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n987), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n870), .A2(new_n871), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n440), .A2(new_n384), .ZN(new_n996));
  INV_X1    g810(.A(new_n397), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n986), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(KEYINPUT126), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n990), .A2(new_n993), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1001), .B(new_n1002), .C1(new_n995), .C2(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1000), .A2(new_n1003), .ZN(G57));
endmodule


