//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  INV_X1    g0004(.A(G238), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n211), .C1(G107), .C2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  AND2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n203), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT0), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(G58), .A2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n231), .A2(new_n233), .A3(G50), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n226), .A2(new_n227), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n228), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n224), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(KEYINPUT65), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n221), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n242), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G68), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G107), .B(G116), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n256), .B(new_n258), .C1(new_n259), .C2(new_n257), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n260), .B(new_n263), .C1(G77), .C2(new_n256), .ZN(new_n264));
  OR2_X1    g0064(.A1(G41), .A2(G45), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n266), .A3(G274), .ZN(new_n267));
  AND2_X1   g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n265), .A2(new_n266), .B1(new_n268), .B2(new_n261), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G226), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n264), .A2(G190), .A3(new_n267), .A4(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(new_n267), .A3(new_n270), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G200), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n277), .A2(new_n229), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G1), .B2(new_n230), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n229), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n230), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR3_X1   g0085(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n230), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n286), .A2(new_n230), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n282), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n276), .B(new_n281), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n271), .B(new_n273), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n295), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n299), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT10), .B1(new_n301), .B2(new_n296), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n272), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G179), .B2(new_n272), .ZN(new_n306));
  INV_X1    g0106(.A(new_n294), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT71), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n274), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n217), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n280), .A2(KEYINPUT71), .A3(G77), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT70), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n314));
  INV_X1    g0114(.A(new_n288), .ZN(new_n315));
  OR2_X1    g0115(.A1(KEYINPUT8), .A2(G58), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g0117(.A1(KEYINPUT8), .A2(G58), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT15), .B(G87), .Z(new_n321));
  INV_X1    g0121(.A(new_n284), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(new_n322), .B1(G20), .B2(G77), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n313), .B1(new_n324), .B2(new_n282), .ZN(new_n325));
  AOI211_X1 g0125(.A(KEYINPUT70), .B(new_n278), .C1(new_n320), .C2(new_n323), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n311), .B(new_n312), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n329));
  INV_X1    g0129(.A(G274), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n262), .A2(new_n329), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n218), .ZN(new_n333));
  AND2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  NOR2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT68), .B1(new_n336), .B2(new_n205), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G1698), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(G107), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT68), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n336), .B2(new_n221), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n256), .A2(KEYINPUT68), .A3(G232), .A4(new_n257), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  AOI211_X1 g0143(.A(new_n331), .B(new_n333), .C1(new_n343), .C2(new_n263), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G190), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n263), .ZN(new_n346));
  INV_X1    g0146(.A(new_n333), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n267), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G200), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n328), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT72), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n346), .A2(new_n352), .A3(new_n267), .A4(new_n347), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n327), .B(new_n353), .C1(new_n344), .C2(G169), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n350), .B2(new_n354), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n303), .B(new_n308), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n259), .A2(new_n257), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n216), .A2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n334), .C2(new_n335), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G33), .A2(G87), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n263), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n331), .B1(new_n269), .B2(G232), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n262), .B1(new_n361), .B2(new_n362), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n267), .B1(new_n332), .B2(new_n221), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT77), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(G200), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n368), .A2(new_n369), .A3(G190), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n287), .ZN(new_n376));
  NAND2_X1  g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n230), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n376), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n377), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n204), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n220), .A2(new_n204), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n232), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n315), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n374), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n336), .B2(new_n230), .ZN(new_n388));
  INV_X1    g0188(.A(new_n381), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n386), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(new_n392), .A3(new_n282), .ZN(new_n393));
  MUX2_X1   g0193(.A(new_n279), .B(new_n274), .S(new_n283), .Z(new_n394));
  NAND4_X1  g0194(.A1(new_n373), .A2(KEYINPUT17), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(new_n394), .C1(new_n371), .C2(new_n372), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n394), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n368), .A2(new_n369), .A3(G179), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n367), .A2(new_n370), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n304), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(KEYINPUT18), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT78), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n400), .A2(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n405), .A3(new_n408), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n399), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n358), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(G226), .B(new_n257), .C1(new_n334), .C2(new_n335), .ZN(new_n414));
  OAI211_X1 g0214(.A(G232), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(new_n287), .C2(new_n209), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n263), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n269), .A2(G238), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n267), .ZN(new_n419));
  OR2_X1    g0219(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(KEYINPUT76), .A2(G169), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n331), .B1(new_n416), .B2(new_n263), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n424), .A2(KEYINPUT74), .A3(KEYINPUT13), .A4(new_n418), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT14), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT13), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(KEYINPUT75), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n429), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n424), .A2(new_n431), .A3(new_n418), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(G179), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n422), .A2(new_n434), .A3(new_n423), .A4(new_n425), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n274), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(KEYINPUT12), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT12), .B1(new_n279), .B2(new_n309), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(G68), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n310), .A2(KEYINPUT12), .A3(new_n204), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n284), .A2(new_n217), .B1(new_n230), .B2(G68), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n288), .A2(new_n215), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n282), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n444), .A2(KEYINPUT11), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(KEYINPUT11), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n440), .B(new_n441), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n422), .A2(G200), .A3(new_n425), .ZN(new_n449));
  INV_X1    g0249(.A(new_n447), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n430), .A2(G190), .A3(new_n432), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n448), .B(new_n453), .C1(new_n357), .C2(KEYINPUT73), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n274), .A2(new_n309), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n274), .A2(new_n309), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n278), .B(G116), .C1(G1), .C2(new_n287), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(new_n310), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(G20), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n282), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT84), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT84), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n282), .A2(new_n465), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n230), .C1(G33), .C2(new_n209), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT20), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AOI221_X4 g0270(.A(KEYINPUT84), .B1(new_n455), .B2(G20), .C1(new_n277), .C2(new_n229), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n465), .B1(new_n282), .B2(new_n462), .ZN(new_n472));
  OAI211_X1 g0272(.A(KEYINPUT20), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n461), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n257), .A2(G257), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G264), .A2(G1698), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n477), .C1(new_n334), .C2(new_n335), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT83), .B(G303), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n263), .C1(new_n256), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  INV_X1    g0281(.A(G45), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G270), .A3(new_n262), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(G274), .A3(new_n483), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G169), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n475), .A2(KEYINPUT21), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT21), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n460), .B1(new_n494), .B2(new_n473), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n491), .B1(new_n495), .B2(new_n488), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n487), .A2(new_n352), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n475), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n230), .B(G87), .C1(new_n334), .C2(new_n335), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT85), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(KEYINPUT22), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n256), .A2(new_n230), .A3(G87), .A4(new_n502), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(KEYINPUT22), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  INV_X1    g0308(.A(G107), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(G20), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G20), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n508), .A2(new_n509), .A3(G20), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT87), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(new_n508), .A3(new_n509), .A4(G20), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n513), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n507), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n507), .A2(KEYINPUT24), .A3(new_n511), .A4(new_n518), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n282), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n278), .B(new_n274), .C1(G1), .C2(new_n287), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G107), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n274), .A2(G107), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n527), .B(KEYINPUT25), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n523), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n208), .A2(new_n257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n210), .A2(G1698), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(new_n334), .C2(new_n335), .ZN(new_n532));
  INV_X1    g0332(.A(G294), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n287), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n262), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n481), .A2(new_n483), .B1(new_n268), .B2(new_n261), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n536), .A2(KEYINPUT88), .B1(G264), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT88), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n376), .A2(new_n377), .B1(new_n210), .B2(G1698), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n534), .B1(new_n540), .B2(new_n530), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n262), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n538), .A2(new_n542), .A3(new_n486), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n484), .A2(G264), .A3(new_n262), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(new_n486), .C1(new_n541), .C2(new_n262), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n543), .A2(new_n304), .B1(new_n352), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n529), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(G190), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n538), .A2(new_n542), .A3(new_n548), .A4(new_n486), .ZN(new_n549));
  INV_X1    g0349(.A(G200), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n523), .A2(new_n552), .A3(new_n526), .A4(new_n528), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n487), .A2(new_n548), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(G200), .B2(new_n487), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n495), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n499), .A2(new_n547), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n266), .A2(G45), .A3(G274), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT80), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(G1698), .C1(new_n334), .C2(new_n335), .ZN(new_n560));
  OAI211_X1 g0360(.A(G238), .B(new_n257), .C1(new_n334), .C2(new_n335), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(new_n512), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n559), .B1(new_n562), .B2(new_n263), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n262), .B(G250), .C1(G1), .C2(new_n482), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n304), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n263), .ZN(new_n567));
  INV_X1    g0367(.A(new_n559), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n567), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n352), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT82), .ZN(new_n571));
  NAND3_X1  g0371(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n230), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n207), .A2(new_n209), .A3(new_n509), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT81), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n256), .A2(new_n230), .A3(G68), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n284), .B2(new_n209), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(new_n580), .A3(new_n574), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n576), .A2(new_n577), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n282), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n437), .A2(KEYINPUT71), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n274), .A2(new_n309), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n321), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n525), .A2(new_n321), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n571), .A2(new_n583), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n582), .B2(new_n282), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n571), .B1(new_n590), .B2(new_n588), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n566), .B(new_n570), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n274), .A2(G97), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n524), .A2(new_n209), .ZN(new_n594));
  OAI21_X1  g0394(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n209), .A2(new_n509), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n509), .A2(KEYINPUT6), .A3(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G20), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n288), .A2(new_n217), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n595), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n593), .B(new_n594), .C1(new_n605), .C2(new_n282), .ZN(new_n606));
  OAI211_X1 g0406(.A(G244), .B(new_n257), .C1(new_n334), .C2(new_n335), .ZN(new_n607));
  NOR2_X1   g0407(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n608), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n256), .A2(G244), .A3(new_n257), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n609), .A2(new_n611), .A3(new_n468), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n263), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n537), .A2(G257), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n486), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n613), .A2(new_n263), .B1(G257), .B2(new_n537), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(G190), .A3(new_n486), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n606), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n563), .A2(G190), .A3(new_n564), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n550), .B1(new_n563), .B2(new_n564), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n525), .A2(G87), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n590), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n616), .A2(new_n304), .ZN(new_n626));
  INV_X1    g0426(.A(new_n593), .ZN(new_n627));
  INV_X1    g0427(.A(new_n594), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n509), .B1(new_n380), .B2(new_n381), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n230), .B1(new_n599), .B2(new_n600), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n629), .A2(new_n630), .A3(new_n603), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n627), .B(new_n628), .C1(new_n631), .C2(new_n278), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n618), .A2(new_n352), .A3(new_n486), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n626), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n592), .A2(new_n620), .A3(new_n625), .A4(new_n634), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n413), .A2(new_n454), .A3(new_n557), .A4(new_n635), .ZN(G372));
  NOR2_X1   g0436(.A1(new_n413), .A2(new_n454), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n590), .A2(KEYINPUT89), .A3(new_n624), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT89), .B1(new_n590), .B2(new_n624), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n623), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n592), .A2(new_n553), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n499), .A2(new_n547), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n620), .A2(new_n634), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT90), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n626), .A2(new_n632), .A3(new_n646), .A4(new_n633), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n569), .A2(G169), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT82), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n590), .A2(new_n571), .A3(new_n588), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n583), .A2(new_n587), .A3(new_n624), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT89), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n590), .A2(KEYINPUT89), .A3(new_n624), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n653), .A2(new_n570), .B1(new_n658), .B2(new_n623), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n648), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n634), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n592), .A3(new_n625), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n644), .A2(new_n592), .A3(new_n661), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n637), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n308), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n409), .A2(new_n404), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n448), .ZN(new_n670));
  INV_X1    g0470(.A(new_n354), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n453), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n669), .B1(new_n672), .B2(new_n399), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n303), .B(KEYINPUT91), .Z(new_n674));
  AOI21_X1  g0474(.A(new_n667), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n666), .A2(new_n675), .ZN(G369));
  NAND3_X1  g0476(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n677));
  INV_X1    g0477(.A(G13), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G20), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n266), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n495), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n677), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n499), .A2(new_n556), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT92), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT92), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n547), .A2(new_n553), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n529), .A2(new_n685), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n529), .A2(new_n546), .A3(new_n685), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n691), .A2(G330), .A3(new_n692), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n499), .A2(new_n685), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n529), .A2(new_n546), .A3(new_n686), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n225), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G1), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n598), .A2(new_n207), .A3(new_n455), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n233), .A2(G50), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n708), .A2(new_n709), .B1(new_n710), .B2(new_n707), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n545), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n618), .B2(new_n486), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT93), .ZN(new_n716));
  AOI21_X1  g0516(.A(G179), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n616), .A2(new_n545), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(KEYINPUT93), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n720), .A3(new_n565), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n497), .A2(new_n569), .A3(new_n618), .A4(new_n714), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT30), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n686), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n557), .A2(new_n635), .A3(new_n685), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n722), .A2(new_n729), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n487), .B(new_n565), .C1(new_n715), .C2(new_n716), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n352), .B1(new_n719), .B2(KEYINPUT93), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n713), .B1(new_n728), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n665), .A2(new_n686), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT94), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n665), .A2(new_n740), .A3(new_n686), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n644), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n592), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n648), .A2(new_n659), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(KEYINPUT26), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n620), .A2(new_n634), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n547), .B2(new_n499), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(KEYINPUT95), .A3(new_n641), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n744), .A2(new_n747), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(KEYINPUT29), .A3(new_n686), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n736), .B1(new_n742), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n712), .B1(new_n754), .B2(G1), .ZN(G364));
  AOI21_X1  g0555(.A(new_n708), .B1(G45), .B2(new_n679), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n229), .B1(G20), .B2(new_n304), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n251), .A2(new_n482), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n705), .A2(new_n256), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(G45), .B2(new_n710), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n763), .A2(new_n765), .B1(G116), .B2(new_n225), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n705), .A2(new_n336), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(G355), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n230), .A2(G190), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(G179), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n230), .A2(new_n352), .A3(new_n548), .A4(new_n550), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G68), .A2(new_n771), .B1(new_n772), .B2(G50), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT32), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n230), .B1(new_n775), .B2(G190), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n773), .B1(new_n774), .B2(new_n778), .C1(new_n209), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n550), .A2(G179), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT97), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n230), .A2(new_n548), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n256), .B1(new_n784), .B2(new_n207), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT98), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n782), .A2(new_n769), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G107), .ZN(new_n789));
  OAI211_X1 g0589(.A(KEYINPUT98), .B(new_n256), .C1(new_n784), .C2(new_n207), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT99), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n783), .A2(G179), .A3(new_n550), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n780), .B(new_n792), .C1(G58), .C2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n769), .A2(G179), .A3(new_n550), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G77), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n778), .A2(new_n774), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n795), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT100), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n770), .A2(new_n803), .B1(new_n793), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  INV_X1    g0606(.A(new_n776), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G326), .A2(new_n772), .B1(new_n807), .B2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(new_n788), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n336), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n806), .B(new_n811), .C1(G311), .C2(new_n797), .ZN(new_n812));
  INV_X1    g0612(.A(G303), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n533), .B2(new_n779), .C1(new_n813), .C2(new_n784), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n800), .A2(new_n801), .ZN(new_n815));
  AND3_X1   g0615(.A1(new_n802), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n760), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n756), .B1(new_n762), .B2(new_n768), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT102), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n691), .A2(new_n692), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n818), .A2(KEYINPUT102), .B1(new_n820), .B2(new_n759), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n713), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n691), .A2(G330), .A3(new_n692), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT96), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n756), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n819), .A2(new_n821), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NOR2_X1   g0629(.A1(new_n354), .A2(new_n685), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n350), .B1(new_n328), .B2(new_n686), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(new_n354), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n738), .A2(new_n741), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n665), .A2(new_n686), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(new_n736), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n826), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n788), .A2(G87), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n776), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT104), .Z(new_n842));
  XOR2_X1   g0642(.A(KEYINPUT103), .B(G283), .Z(new_n843));
  AOI211_X1 g0643(.A(new_n256), .B(new_n842), .C1(new_n771), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n509), .B2(new_n784), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n796), .A2(new_n455), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n793), .A2(new_n533), .ZN(new_n847));
  INV_X1    g0647(.A(new_n772), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n848), .A2(new_n813), .B1(new_n779), .B2(new_n209), .ZN(new_n849));
  NOR4_X1   g0649(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G143), .A2(new_n794), .B1(new_n771), .B2(G150), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n852), .B2(new_n848), .C1(new_n777), .C2(new_n796), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT34), .Z(new_n854));
  NOR2_X1   g0654(.A1(new_n779), .A2(new_n220), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n788), .A2(G68), .ZN(new_n856));
  INV_X1    g0656(.A(G132), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n776), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n256), .B1(new_n784), .B2(new_n215), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n854), .A2(new_n855), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n760), .B1(new_n850), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n760), .A2(new_n757), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n217), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n833), .A2(new_n757), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n861), .A2(new_n756), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n838), .A2(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n448), .A2(new_n685), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n683), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n400), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n407), .A2(new_n870), .A3(new_n396), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n407), .A2(new_n870), .A3(new_n873), .A4(new_n396), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n412), .B2(new_n870), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT38), .B(new_n875), .C1(new_n412), .C2(new_n870), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(KEYINPUT106), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n876), .A2(new_n881), .A3(new_n877), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n870), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n668), .B2(new_n399), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n885), .B2(new_n875), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n410), .A2(new_n411), .ZN(new_n887));
  INV_X1    g0687(.A(new_n399), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n889), .A2(new_n884), .B1(new_n872), .B2(new_n874), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n890), .B2(KEYINPUT38), .ZN(new_n891));
  XOR2_X1   g0691(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n868), .B1(new_n883), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n830), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n835), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n450), .A2(new_n686), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n898), .B(new_n452), .C1(new_n436), .C2(new_n447), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n448), .A2(new_n686), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n880), .A2(new_n897), .A3(new_n901), .A4(new_n882), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n668), .A2(new_n683), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n742), .A2(new_n637), .A3(new_n753), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n675), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n832), .B1(new_n899), .B2(new_n900), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n735), .A2(KEYINPUT108), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT108), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n724), .A2(new_n912), .A3(KEYINPUT31), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n910), .B1(new_n915), .B2(new_n728), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n916), .A2(new_n880), .A3(new_n917), .A4(new_n882), .ZN(new_n918));
  INV_X1    g0718(.A(new_n635), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n677), .B1(new_n495), .B2(new_n555), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(new_n693), .A3(new_n920), .A4(new_n686), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n724), .B1(new_n921), .B2(KEYINPUT31), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n901), .B(new_n832), .C1(new_n922), .C2(new_n914), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT40), .B1(new_n923), .B2(new_n891), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n918), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(G330), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n915), .A2(new_n728), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n637), .A2(G330), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n637), .A3(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n909), .B(new_n931), .Z(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n266), .B2(new_n679), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n601), .B(KEYINPUT105), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n455), .B1(new_n934), .B2(KEYINPUT35), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n231), .C1(KEYINPUT35), .C2(new_n934), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  OAI21_X1  g0737(.A(G77), .B1(new_n220), .B2(new_n204), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n710), .A2(new_n938), .B1(G50), .B2(new_n204), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(G1), .A3(new_n678), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n937), .A3(new_n940), .ZN(G367));
  INV_X1    g0741(.A(new_n764), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n242), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n321), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n761), .B1(new_n225), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n784), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(G58), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n788), .A2(G77), .ZN(new_n948));
  INV_X1    g0748(.A(new_n779), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n797), .A2(G50), .B1(new_n949), .B2(G68), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G143), .A2(new_n772), .B1(new_n807), .B2(G137), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n336), .B(new_n952), .C1(G159), .C2(new_n771), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n794), .A2(G150), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n772), .A2(G311), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n946), .A2(KEYINPUT46), .A3(G116), .ZN(new_n956));
  INV_X1    g0756(.A(G317), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n957), .B2(new_n776), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n788), .A2(G97), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n771), .A2(G294), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n794), .A2(new_n479), .B1(new_n949), .B2(G107), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n256), .B1(new_n797), .B2(new_n843), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT46), .B1(new_n946), .B2(G116), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n958), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n756), .B1(new_n943), .B2(new_n945), .C1(new_n967), .C2(new_n817), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT114), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n658), .A2(new_n686), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  MUX2_X1   g0771(.A(new_n745), .B(new_n659), .S(new_n971), .Z(new_n972));
  OR3_X1    g0772(.A1(new_n972), .A2(G20), .A3(new_n758), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n266), .B1(new_n679), .B2(G45), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n643), .B1(new_n606), .B2(new_n686), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n662), .A2(new_n685), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n702), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT44), .ZN(new_n982));
  XOR2_X1   g0782(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n979), .B2(new_n702), .ZN(new_n985));
  INV_X1    g0785(.A(new_n979), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n986), .A2(new_n703), .A3(new_n983), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n981), .A2(new_n982), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT113), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n698), .ZN(new_n990));
  INV_X1    g0790(.A(new_n698), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(KEYINPUT113), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n700), .B1(new_n697), .B2(new_n699), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n823), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n825), .B2(new_n994), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n754), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n754), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n706), .B(KEYINPUT41), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n976), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n698), .A2(KEYINPUT110), .A3(new_n979), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT110), .B1(new_n698), .B2(new_n979), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n750), .A2(new_n693), .A3(new_n699), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT42), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n634), .B1(new_n977), .B2(new_n547), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n686), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1007), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n974), .B1(new_n1000), .B2(new_n1018), .ZN(G387));
  NAND2_X1  g0819(.A1(new_n996), .A2(new_n976), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n314), .A2(new_n319), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(G50), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT50), .Z(new_n1023));
  NOR2_X1   g0823(.A1(new_n204), .A2(new_n217), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1023), .A2(G45), .A3(new_n1024), .A4(new_n709), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n942), .B1(new_n246), .B2(G45), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n709), .B2(new_n767), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1025), .A2(new_n1027), .B1(G107), .B2(new_n225), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1028), .A2(new_n761), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G317), .A2(new_n794), .B1(new_n771), .B2(G311), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n804), .B2(new_n848), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n479), .B2(new_n797), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT48), .Z(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n533), .B2(new_n784), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n949), .B2(new_n843), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT49), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n256), .B1(new_n807), .B2(G326), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n809), .B2(new_n455), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n946), .A2(G77), .B1(G159), .B2(new_n772), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n215), .B2(new_n793), .C1(new_n289), .C2(new_n776), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n959), .B1(new_n204), .B2(new_n796), .C1(new_n283), .C2(new_n770), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n944), .A2(new_n779), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n336), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n760), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n695), .A2(new_n696), .A3(new_n759), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n756), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n997), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n706), .B1(new_n996), .B2(new_n754), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1020), .B1(new_n1029), .B2(new_n1047), .C1(new_n1048), .C2(new_n1049), .ZN(G393));
  NOR2_X1   g0850(.A1(new_n993), .A2(new_n997), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT115), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n988), .B(new_n991), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n997), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1051), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n997), .A2(new_n1053), .A3(KEYINPUT115), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n706), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1053), .A2(new_n975), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n779), .A2(new_n455), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n848), .A2(new_n957), .B1(new_n840), .B2(new_n793), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT52), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n256), .B1(new_n946), .B2(new_n843), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1063), .A2(new_n789), .A3(new_n1064), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n533), .B2(new_n796), .C1(new_n804), .C2(new_n776), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1061), .B(new_n1066), .C1(new_n479), .C2(new_n771), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n848), .A2(new_n289), .B1(new_n777), .B2(new_n793), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n256), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n771), .A2(G50), .B1(new_n949), .B2(G77), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n839), .B(new_n1071), .C1(new_n204), .C2(new_n784), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1021), .A2(new_n796), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n807), .A2(G143), .ZN(new_n1074));
  NOR4_X1   g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n760), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n761), .B1(new_n209), .B2(new_n225), .C1(new_n254), .C2(new_n942), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n979), .A2(new_n759), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1076), .A2(new_n756), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1059), .A2(new_n1060), .A3(new_n1079), .ZN(G390));
  NAND3_X1  g0880(.A1(new_n883), .A2(new_n757), .A3(new_n893), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n862), .A2(new_n283), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n336), .B1(new_n784), .B2(new_n207), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT118), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1084), .A2(new_n856), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n209), .B2(new_n796), .C1(new_n509), .C2(new_n770), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n776), .A2(new_n533), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n793), .A2(new_n455), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n848), .A2(new_n810), .B1(new_n779), .B2(new_n217), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n784), .A2(new_n289), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT53), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT54), .B(G143), .Z(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n256), .C1(new_n796), .C2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(G128), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n848), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n770), .A2(new_n852), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G125), .A2(new_n807), .B1(new_n949), .B2(G159), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n857), .B2(new_n793), .C1(new_n809), .C2(new_n215), .ZN(new_n1100));
  NOR4_X1   g0900(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n760), .B1(new_n1090), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1081), .A2(new_n756), .A3(new_n1082), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n883), .A2(new_n893), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n867), .B1(new_n897), .B2(new_n901), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n899), .A2(new_n900), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n831), .A2(new_n354), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n752), .A2(new_n686), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1106), .B1(new_n1108), .B2(new_n896), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n891), .A2(new_n867), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1104), .A2(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n910), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(G330), .C1(new_n922), .C2(new_n914), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n897), .A2(new_n901), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n868), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n883), .A3(new_n893), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n891), .A2(new_n867), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1108), .A2(new_n896), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n1106), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n736), .A2(new_n832), .A3(new_n901), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1115), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1103), .B1(new_n1124), .B2(new_n975), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n907), .A2(new_n675), .A3(new_n928), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n735), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n832), .C1(new_n922), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1106), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1113), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n897), .ZN(new_n1132));
  OAI211_X1 g0932(.A(G330), .B(new_n832), .C1(new_n922), .C2(new_n914), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1106), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1120), .A2(new_n1122), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1127), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT116), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n907), .A2(new_n675), .A3(new_n928), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT116), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1138), .A2(new_n1142), .B1(new_n1123), .B2(new_n1115), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n1115), .A3(new_n1123), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n706), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1143), .A2(new_n1145), .A3(KEYINPUT117), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT117), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1113), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n707), .B1(new_n1150), .B2(new_n1136), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n897), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1130), .B2(new_n1113), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1122), .A2(new_n1134), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n1120), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1155), .A2(KEYINPUT116), .A3(new_n1127), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1137), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1124), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1147), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1126), .B1(new_n1146), .B2(new_n1159), .ZN(G378));
  NAND3_X1  g0960(.A1(new_n926), .A2(new_n895), .A3(new_n905), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n674), .A2(new_n308), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n294), .A2(new_n869), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1162), .B(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n713), .B1(new_n918), .B2(new_n924), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n904), .B2(new_n894), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1161), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1166), .B1(new_n1161), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n862), .A2(new_n215), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1166), .B2(new_n758), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n788), .A2(G58), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT119), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n797), .A2(new_n321), .B1(new_n949), .B2(G68), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n256), .B1(new_n771), .B2(G97), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n794), .A2(G107), .B1(new_n807), .B2(G283), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n455), .B2(new_n848), .C1(new_n784), .C2(new_n217), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1178), .A2(G41), .A3(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT58), .Z(new_n1182));
  OAI21_X1  g0982(.A(new_n215), .B1(new_n334), .B2(G41), .ZN(new_n1183));
  INV_X1    g0983(.A(G124), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n287), .B1(new_n776), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n779), .A2(new_n289), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n793), .A2(new_n1096), .B1(new_n770), .B2(new_n857), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(G125), .C2(new_n772), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n852), .B2(new_n796), .C1(new_n784), .C2(new_n1094), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G41), .B(new_n1185), .C1(new_n1189), .C2(KEYINPUT59), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(KEYINPUT59), .B2(new_n1189), .C1(new_n777), .C2(new_n809), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1182), .A2(new_n1183), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1173), .B1(new_n760), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1171), .A2(new_n976), .B1(new_n756), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT120), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1127), .B(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1144), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1161), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1166), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1168), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1167), .A2(new_n894), .A3(new_n904), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1197), .A2(KEYINPUT57), .A3(new_n1198), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n706), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1197), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1194), .B1(new_n1204), .B2(new_n1205), .ZN(G375));
  INV_X1    g1006(.A(KEYINPUT121), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1155), .B2(new_n975), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1106), .A2(new_n757), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n862), .A2(new_n204), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1175), .B1(new_n857), .B2(new_n848), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n776), .A2(new_n1096), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1094), .A2(new_n770), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n794), .A2(G137), .B1(new_n949), .B2(G50), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n336), .B1(new_n797), .B2(G150), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n784), .C2(new_n777), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n946), .A2(G97), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1043), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n797), .A2(G107), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1218), .A2(new_n948), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n848), .A2(new_n533), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n770), .A2(new_n455), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n336), .B1(new_n776), .B2(new_n813), .C1(new_n793), .C2(new_n810), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n760), .B1(new_n1217), .B2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1209), .A2(new_n756), .A3(new_n1210), .A4(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1139), .A2(KEYINPUT121), .A3(new_n976), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1208), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT122), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT122), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1208), .A2(new_n1231), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n999), .B1(new_n1140), .B2(new_n1139), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(G381));
  INV_X1    g1035(.A(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1202), .A2(new_n1198), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1127), .B(KEYINPUT120), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1150), .B2(new_n1136), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1236), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n706), .A3(new_n1203), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1125), .B1(new_n1151), .B2(new_n1158), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1241), .A2(new_n1194), .A3(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G390), .A2(G387), .ZN(new_n1244));
  OR2_X1    g1044(.A1(G396), .A2(G393), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G381), .A2(G384), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .A4(new_n1247), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n684), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G407), .A2(G213), .A3(new_n1249), .ZN(G409));
  AND3_X1   g1050(.A1(new_n1171), .A2(new_n999), .A3(new_n1197), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1193), .A2(new_n756), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1237), .B2(new_n975), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1242), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT117), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1151), .A2(new_n1158), .A3(new_n1147), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1125), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1254), .B1(G375), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n684), .A2(G213), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT60), .B1(new_n1155), .B2(new_n1127), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT123), .B1(new_n1260), .B2(new_n1136), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n707), .B1(new_n1262), .B2(KEYINPUT60), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT123), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1141), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1261), .A2(new_n1263), .A3(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1233), .A2(G384), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1233), .B2(new_n1268), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1258), .A2(new_n1259), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1269), .A2(new_n1270), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT121), .B1(new_n1139), .B2(new_n976), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1207), .B(new_n975), .C1(new_n1132), .C2(new_n1135), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1231), .B1(new_n1280), .B2(new_n1227), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1232), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1268), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1233), .A2(G384), .A3(new_n1268), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1275), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1277), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1274), .A2(new_n1288), .ZN(new_n1289));
  XOR2_X1   g1089(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1258), .A2(new_n1291), .A3(new_n1259), .A4(new_n1271), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1273), .A2(new_n1289), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(G387), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT124), .B1(new_n1294), .B2(G390), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n828), .B(G393), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1079), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(G387), .A2(new_n1298), .A3(new_n1060), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G387), .B1(new_n1298), .B2(new_n1060), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n1295), .A2(new_n1296), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1296), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1294), .A2(G390), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(KEYINPUT124), .A4(new_n1299), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1302), .A2(KEYINPUT126), .A3(new_n1305), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1293), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(G378), .A2(new_n1194), .A3(new_n1241), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1312), .A2(new_n1254), .B1(G213), .B2(new_n684), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1276), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1285), .A2(new_n1286), .A3(new_n1275), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT63), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1272), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1259), .A4(new_n1271), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1319), .A2(new_n1320), .A3(new_n1306), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1311), .A2(new_n1322), .ZN(G405));
  INV_X1    g1123(.A(new_n1271), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(G375), .A2(new_n1325), .A3(new_n1242), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(G375), .B2(new_n1242), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1324), .B1(new_n1329), .B2(new_n1312), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1242), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT127), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1312), .A3(new_n1326), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1333), .A2(new_n1271), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1310), .B1(new_n1330), .B2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1329), .A2(new_n1312), .A3(new_n1324), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1333), .A2(new_n1271), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1336), .A2(new_n1337), .A3(new_n1309), .A4(new_n1308), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1335), .A2(new_n1338), .ZN(G402));
endmodule


