

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G543), .A2(G651), .ZN(n796) );
  NAND2_X1 U550 ( .A1(n655), .A2(n656), .ZN(n694) );
  XNOR2_X1 U551 ( .A(KEYINPUT89), .B(n589), .ZN(n656) );
  NOR2_X1 U552 ( .A1(G651), .A2(n567), .ZN(n799) );
  XOR2_X1 U553 ( .A(KEYINPUT1), .B(n528), .Z(n803) );
  XNOR2_X1 U554 ( .A(KEYINPUT103), .B(KEYINPUT40), .ZN(n757) );
  XNOR2_X1 U555 ( .A(n758), .B(n757), .ZN(G329) );
  INV_X1 U556 ( .A(G2104), .ZN(n517) );
  NOR2_X1 U557 ( .A1(G2105), .A2(n517), .ZN(n967) );
  NAND2_X1 U558 ( .A1(n967), .A2(G102), .ZN(n512) );
  XNOR2_X1 U559 ( .A(n512), .B(KEYINPUT88), .ZN(n516) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n513) );
  XOR2_X1 U561 ( .A(KEYINPUT17), .B(n513), .Z(n514) );
  XNOR2_X2 U562 ( .A(KEYINPUT64), .B(n514), .ZN(n968) );
  NAND2_X1 U563 ( .A1(G138), .A2(n968), .ZN(n515) );
  NAND2_X1 U564 ( .A1(n516), .A2(n515), .ZN(n521) );
  AND2_X1 U565 ( .A1(n517), .A2(G2105), .ZN(n963) );
  NAND2_X1 U566 ( .A1(G126), .A2(n963), .ZN(n519) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n964) );
  NAND2_X1 U568 ( .A1(G114), .A2(n964), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U570 ( .A1(n521), .A2(n520), .ZN(G164) );
  XOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .Z(n567) );
  XOR2_X1 U572 ( .A(KEYINPUT66), .B(G651), .Z(n527) );
  OR2_X1 U573 ( .A1(n567), .A2(n527), .ZN(n522) );
  XNOR2_X1 U574 ( .A(n522), .B(KEYINPUT67), .ZN(n795) );
  AND2_X1 U575 ( .A1(n795), .A2(G72), .ZN(n526) );
  NAND2_X1 U576 ( .A1(G47), .A2(n799), .ZN(n524) );
  NAND2_X1 U577 ( .A1(G85), .A2(n796), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G543), .A2(n527), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n803), .A2(G60), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(G290) );
  NAND2_X1 U583 ( .A1(G52), .A2(n799), .ZN(n532) );
  NAND2_X1 U584 ( .A1(G64), .A2(n803), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n537) );
  NAND2_X1 U586 ( .A1(G77), .A2(n795), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G90), .A2(n796), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U589 ( .A(KEYINPUT9), .B(n535), .Z(n536) );
  NOR2_X1 U590 ( .A1(n537), .A2(n536), .ZN(G171) );
  INV_X1 U591 ( .A(G171), .ZN(G301) );
  NAND2_X1 U592 ( .A1(G65), .A2(n803), .ZN(n538) );
  XNOR2_X1 U593 ( .A(n538), .B(KEYINPUT68), .ZN(n545) );
  NAND2_X1 U594 ( .A1(G78), .A2(n795), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G91), .A2(n796), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G53), .A2(n799), .ZN(n541) );
  XNOR2_X1 U598 ( .A(KEYINPUT69), .B(n541), .ZN(n542) );
  NOR2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U601 ( .A(KEYINPUT70), .B(n546), .ZN(G299) );
  NAND2_X1 U602 ( .A1(G51), .A2(n799), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G63), .A2(n803), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U605 ( .A(KEYINPUT6), .B(n549), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n796), .A2(G89), .ZN(n550) );
  XNOR2_X1 U607 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G76), .A2(n795), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U610 ( .A(n553), .B(KEYINPUT5), .Z(n554) );
  NOR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT78), .B(n556), .Z(n557) );
  XNOR2_X1 U613 ( .A(KEYINPUT7), .B(n557), .ZN(G168) );
  NAND2_X1 U614 ( .A1(n803), .A2(G62), .ZN(n558) );
  XOR2_X1 U615 ( .A(KEYINPUT81), .B(n558), .Z(n560) );
  NAND2_X1 U616 ( .A1(n799), .A2(G50), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U618 ( .A(KEYINPUT82), .B(n561), .ZN(n564) );
  NAND2_X1 U619 ( .A1(G75), .A2(n795), .ZN(n562) );
  XNOR2_X1 U620 ( .A(KEYINPUT83), .B(n562), .ZN(n563) );
  NOR2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n796), .A2(G88), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n566), .A2(n565), .ZN(G303) );
  XOR2_X1 U624 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U625 ( .A1(G87), .A2(n567), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G74), .A2(G651), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U628 ( .A1(n803), .A2(n570), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n799), .A2(G49), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(G288) );
  XOR2_X1 U631 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n574) );
  NAND2_X1 U632 ( .A1(G73), .A2(n795), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n574), .B(n573), .ZN(n578) );
  NAND2_X1 U634 ( .A1(G48), .A2(n799), .ZN(n576) );
  NAND2_X1 U635 ( .A1(G86), .A2(n796), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U637 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U638 ( .A1(n803), .A2(G61), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n580), .A2(n579), .ZN(G305) );
  NOR2_X1 U640 ( .A1(G164), .A2(G1384), .ZN(n655) );
  NAND2_X1 U641 ( .A1(n968), .A2(G137), .ZN(n581) );
  XOR2_X1 U642 ( .A(n581), .B(KEYINPUT65), .Z(n584) );
  NAND2_X1 U643 ( .A1(G101), .A2(n967), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT23), .B(n582), .Z(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n771) );
  NAND2_X1 U646 ( .A1(G125), .A2(n963), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G113), .A2(n964), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n770) );
  INV_X1 U649 ( .A(n770), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G40), .A2(n587), .ZN(n588) );
  OR2_X1 U651 ( .A1(n771), .A2(n588), .ZN(n589) );
  INV_X1 U652 ( .A(n656), .ZN(n590) );
  NOR2_X1 U653 ( .A1(n655), .A2(n590), .ZN(n591) );
  XOR2_X1 U654 ( .A(KEYINPUT90), .B(n591), .Z(n748) );
  NAND2_X1 U655 ( .A1(n963), .A2(G128), .ZN(n592) );
  XNOR2_X1 U656 ( .A(KEYINPUT92), .B(n592), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n964), .A2(G116), .ZN(n593) );
  XOR2_X1 U658 ( .A(KEYINPUT93), .B(n593), .Z(n594) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(n596), .B(KEYINPUT35), .ZN(n602) );
  XNOR2_X1 U661 ( .A(KEYINPUT91), .B(KEYINPUT34), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G104), .A2(n967), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G140), .A2(n968), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U665 ( .A(n600), .B(n599), .ZN(n601) );
  NAND2_X1 U666 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U667 ( .A(KEYINPUT36), .B(n603), .ZN(n988) );
  XOR2_X1 U668 ( .A(G2067), .B(KEYINPUT37), .Z(n604) );
  NOR2_X1 U669 ( .A1(n988), .A2(n604), .ZN(n898) );
  NAND2_X1 U670 ( .A1(n988), .A2(n604), .ZN(n874) );
  NOR2_X1 U671 ( .A1(n748), .A2(n874), .ZN(n746) );
  NAND2_X1 U672 ( .A1(G129), .A2(n963), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G141), .A2(n968), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n967), .A2(G105), .ZN(n607) );
  XOR2_X1 U676 ( .A(KEYINPUT38), .B(n607), .Z(n608) );
  NOR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n964), .A2(G117), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n979) );
  NOR2_X1 U680 ( .A1(G1996), .A2(n979), .ZN(n880) );
  NAND2_X1 U681 ( .A1(G107), .A2(n964), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n612), .B(KEYINPUT94), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n968), .A2(G131), .ZN(n613) );
  XOR2_X1 U684 ( .A(KEYINPUT95), .B(n613), .Z(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U686 ( .A1(G95), .A2(n967), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G119), .A2(n963), .ZN(n616) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n984) );
  INV_X1 U690 ( .A(G1991), .ZN(n622) );
  NOR2_X1 U691 ( .A1(n984), .A2(n622), .ZN(n621) );
  AND2_X1 U692 ( .A1(G1996), .A2(n979), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n875) );
  NOR2_X1 U694 ( .A1(n748), .A2(n875), .ZN(n745) );
  AND2_X1 U695 ( .A1(n622), .A2(n984), .ZN(n871) );
  NOR2_X1 U696 ( .A1(G1986), .A2(G290), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n871), .A2(n623), .ZN(n624) );
  NOR2_X1 U698 ( .A1(n745), .A2(n624), .ZN(n625) );
  NOR2_X1 U699 ( .A1(n880), .A2(n625), .ZN(n626) );
  XOR2_X1 U700 ( .A(KEYINPUT39), .B(n626), .Z(n627) );
  NOR2_X1 U701 ( .A1(n746), .A2(n627), .ZN(n628) );
  NOR2_X1 U702 ( .A1(n898), .A2(n628), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n748), .A2(n629), .ZN(n756) );
  NAND2_X1 U704 ( .A1(G1961), .A2(n694), .ZN(n632) );
  AND2_X1 U705 ( .A1(n655), .A2(n656), .ZN(n671) );
  XOR2_X1 U706 ( .A(G2078), .B(KEYINPUT25), .Z(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT98), .B(n630), .ZN(n857) );
  NAND2_X1 U708 ( .A1(n671), .A2(n857), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n688) );
  OR2_X1 U710 ( .A1(G301), .A2(n688), .ZN(n683) );
  NAND2_X1 U711 ( .A1(G54), .A2(n799), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G79), .A2(n795), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G92), .A2(n796), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G66), .A2(n803), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U717 ( .A(KEYINPUT77), .B(n637), .Z(n638) );
  NOR2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U719 ( .A(KEYINPUT15), .B(n640), .Z(n991) );
  NAND2_X1 U720 ( .A1(n799), .A2(G43), .ZN(n641) );
  XNOR2_X1 U721 ( .A(KEYINPUT76), .B(n641), .ZN(n654) );
  NAND2_X1 U722 ( .A1(G68), .A2(n795), .ZN(n646) );
  XOR2_X1 U723 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n643) );
  NAND2_X1 U724 ( .A1(G81), .A2(n796), .ZN(n642) );
  XNOR2_X1 U725 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U726 ( .A(KEYINPUT72), .B(n644), .ZN(n645) );
  NAND2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U728 ( .A(n647), .B(KEYINPUT74), .ZN(n648) );
  XNOR2_X1 U729 ( .A(KEYINPUT13), .B(n648), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n803), .A2(G56), .ZN(n649) );
  XNOR2_X1 U731 ( .A(KEYINPUT14), .B(n649), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U733 ( .A(KEYINPUT75), .B(n652), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n994) );
  AND2_X1 U735 ( .A1(n655), .A2(G1996), .ZN(n657) );
  AND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U737 ( .A(n658), .B(KEYINPUT26), .Z(n660) );
  NAND2_X1 U738 ( .A1(n694), .A2(G1341), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n994), .A2(n661), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n991), .A2(n667), .ZN(n665) );
  NOR2_X1 U742 ( .A1(G2067), .A2(n694), .ZN(n663) );
  NOR2_X1 U743 ( .A1(n671), .A2(G1348), .ZN(n662) );
  NOR2_X1 U744 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U746 ( .A(KEYINPUT99), .B(n666), .Z(n669) );
  OR2_X1 U747 ( .A1(n667), .A2(n991), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n675) );
  NAND2_X1 U749 ( .A1(n671), .A2(G2072), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n670), .B(KEYINPUT27), .ZN(n673) );
  INV_X1 U751 ( .A(G1956), .ZN(n911) );
  NOR2_X1 U752 ( .A1(n911), .A2(n671), .ZN(n672) );
  NOR2_X1 U753 ( .A1(n673), .A2(n672), .ZN(n677) );
  INV_X1 U754 ( .A(G299), .ZN(n676) );
  NAND2_X1 U755 ( .A1(n677), .A2(n676), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n675), .A2(n674), .ZN(n680) );
  NOR2_X1 U757 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U758 ( .A(n678), .B(KEYINPUT28), .Z(n679) );
  NAND2_X1 U759 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U760 ( .A(n681), .B(KEYINPUT29), .Z(n682) );
  NAND2_X1 U761 ( .A1(n683), .A2(n682), .ZN(n709) );
  NOR2_X1 U762 ( .A1(G2084), .A2(n694), .ZN(n707) );
  NAND2_X1 U763 ( .A1(G8), .A2(n694), .ZN(n739) );
  NOR2_X1 U764 ( .A1(n739), .A2(G1966), .ZN(n684) );
  XNOR2_X1 U765 ( .A(n684), .B(KEYINPUT97), .ZN(n711) );
  NAND2_X1 U766 ( .A1(n711), .A2(G8), .ZN(n685) );
  NOR2_X1 U767 ( .A1(n707), .A2(n685), .ZN(n686) );
  XOR2_X1 U768 ( .A(KEYINPUT30), .B(n686), .Z(n687) );
  NOR2_X1 U769 ( .A1(G168), .A2(n687), .ZN(n691) );
  NAND2_X1 U770 ( .A1(G301), .A2(n688), .ZN(n689) );
  XOR2_X1 U771 ( .A(KEYINPUT100), .B(n689), .Z(n690) );
  NOR2_X1 U772 ( .A1(n691), .A2(n690), .ZN(n693) );
  XNOR2_X1 U773 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n692) );
  XNOR2_X1 U774 ( .A(n693), .B(n692), .ZN(n708) );
  INV_X1 U775 ( .A(G8), .ZN(n699) );
  NOR2_X1 U776 ( .A1(G1971), .A2(n739), .ZN(n696) );
  NOR2_X1 U777 ( .A1(G2090), .A2(n694), .ZN(n695) );
  NOR2_X1 U778 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U779 ( .A1(n697), .A2(G303), .ZN(n698) );
  OR2_X1 U780 ( .A1(n699), .A2(n698), .ZN(n701) );
  AND2_X1 U781 ( .A1(n708), .A2(n701), .ZN(n700) );
  NAND2_X1 U782 ( .A1(n709), .A2(n700), .ZN(n705) );
  INV_X1 U783 ( .A(n701), .ZN(n703) );
  AND2_X1 U784 ( .A1(G286), .A2(G8), .ZN(n702) );
  OR2_X1 U785 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U787 ( .A(n706), .B(KEYINPUT32), .ZN(n731) );
  NAND2_X1 U788 ( .A1(G8), .A2(n707), .ZN(n713) );
  NAND2_X1 U789 ( .A1(n709), .A2(n708), .ZN(n710) );
  AND2_X1 U790 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U791 ( .A1(n713), .A2(n712), .ZN(n730) );
  NOR2_X1 U792 ( .A1(G1976), .A2(G288), .ZN(n912) );
  NAND2_X1 U793 ( .A1(n912), .A2(KEYINPUT33), .ZN(n714) );
  NOR2_X1 U794 ( .A1(n714), .A2(n739), .ZN(n716) );
  INV_X1 U795 ( .A(n716), .ZN(n715) );
  AND2_X1 U796 ( .A1(n715), .A2(KEYINPUT33), .ZN(n722) );
  NOR2_X1 U797 ( .A1(n739), .A2(n716), .ZN(n717) );
  NAND2_X1 U798 ( .A1(G1976), .A2(G288), .ZN(n913) );
  AND2_X1 U799 ( .A1(n717), .A2(n913), .ZN(n718) );
  OR2_X1 U800 ( .A1(n722), .A2(n718), .ZN(n720) );
  AND2_X1 U801 ( .A1(n730), .A2(n720), .ZN(n719) );
  NAND2_X1 U802 ( .A1(n731), .A2(n719), .ZN(n728) );
  INV_X1 U803 ( .A(n720), .ZN(n726) );
  NOR2_X1 U804 ( .A1(G1971), .A2(G303), .ZN(n721) );
  NOR2_X1 U805 ( .A1(n912), .A2(n721), .ZN(n724) );
  INV_X1 U806 ( .A(n722), .ZN(n723) );
  AND2_X1 U807 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U808 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U809 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U810 ( .A(G1981), .B(G305), .Z(n908) );
  NAND2_X1 U811 ( .A1(n729), .A2(n908), .ZN(n744) );
  NAND2_X1 U812 ( .A1(n731), .A2(n730), .ZN(n737) );
  NOR2_X1 U813 ( .A1(G2090), .A2(G303), .ZN(n732) );
  NAND2_X1 U814 ( .A1(G8), .A2(n732), .ZN(n735) );
  NOR2_X1 U815 ( .A1(G1981), .A2(G305), .ZN(n733) );
  XOR2_X1 U816 ( .A(n733), .B(KEYINPUT24), .Z(n734) );
  OR2_X1 U817 ( .A1(n739), .A2(n734), .ZN(n738) );
  AND2_X1 U818 ( .A1(n735), .A2(n738), .ZN(n736) );
  NAND2_X1 U819 ( .A1(n737), .A2(n736), .ZN(n742) );
  INV_X1 U820 ( .A(n738), .ZN(n740) );
  OR2_X1 U821 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U822 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U823 ( .A1(n744), .A2(n743), .ZN(n753) );
  OR2_X1 U824 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U825 ( .A(KEYINPUT96), .B(n747), .Z(n751) );
  INV_X1 U826 ( .A(n748), .ZN(n749) );
  XNOR2_X1 U827 ( .A(G1986), .B(G290), .ZN(n916) );
  NAND2_X1 U828 ( .A1(n749), .A2(n916), .ZN(n750) );
  AND2_X1 U829 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U830 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U831 ( .A(n754), .B(KEYINPUT102), .ZN(n755) );
  NOR2_X1 U832 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U833 ( .A(G1341), .B(G2427), .ZN(n768) );
  XOR2_X1 U834 ( .A(G2451), .B(G2430), .Z(n760) );
  XNOR2_X1 U835 ( .A(G1348), .B(G2443), .ZN(n759) );
  XNOR2_X1 U836 ( .A(n760), .B(n759), .ZN(n764) );
  XOR2_X1 U837 ( .A(KEYINPUT105), .B(G2435), .Z(n762) );
  XNOR2_X1 U838 ( .A(G2454), .B(G2438), .ZN(n761) );
  XNOR2_X1 U839 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U840 ( .A(n764), .B(n763), .Z(n766) );
  XNOR2_X1 U841 ( .A(G2446), .B(KEYINPUT104), .ZN(n765) );
  XNOR2_X1 U842 ( .A(n766), .B(n765), .ZN(n767) );
  XNOR2_X1 U843 ( .A(n768), .B(n767), .ZN(n769) );
  AND2_X1 U844 ( .A1(n769), .A2(G14), .ZN(G401) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U846 ( .A(G120), .ZN(G236) );
  INV_X1 U847 ( .A(G57), .ZN(G237) );
  NOR2_X1 U848 ( .A1(n771), .A2(n770), .ZN(G160) );
  XOR2_X1 U849 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n773) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n772) );
  XNOR2_X1 U851 ( .A(n773), .B(n772), .ZN(G223) );
  INV_X1 U852 ( .A(G223), .ZN(n834) );
  NAND2_X1 U853 ( .A1(n834), .A2(G567), .ZN(n774) );
  XOR2_X1 U854 ( .A(KEYINPUT11), .B(n774), .Z(G234) );
  INV_X1 U855 ( .A(G860), .ZN(n794) );
  OR2_X1 U856 ( .A1(n994), .A2(n794), .ZN(G153) );
  NAND2_X1 U857 ( .A1(G868), .A2(G301), .ZN(n776) );
  OR2_X1 U858 ( .A1(n991), .A2(G868), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(G284) );
  NAND2_X1 U860 ( .A1(G868), .A2(G286), .ZN(n778) );
  INV_X1 U861 ( .A(G868), .ZN(n816) );
  NAND2_X1 U862 ( .A1(G299), .A2(n816), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n794), .A2(G559), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n779), .A2(n991), .ZN(n780) );
  XNOR2_X1 U866 ( .A(n780), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n994), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G868), .A2(n991), .ZN(n781) );
  NOR2_X1 U869 ( .A1(G559), .A2(n781), .ZN(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G123), .A2(n963), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n967), .A2(G99), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n964), .A2(G111), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G135), .A2(n968), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n961) );
  XNOR2_X1 U879 ( .A(n961), .B(G2096), .ZN(n792) );
  INV_X1 U880 ( .A(G2100), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(G156) );
  NAND2_X1 U882 ( .A1(G559), .A2(n991), .ZN(n793) );
  XOR2_X1 U883 ( .A(n994), .B(n793), .Z(n813) );
  NAND2_X1 U884 ( .A1(n794), .A2(n813), .ZN(n806) );
  NAND2_X1 U885 ( .A1(G80), .A2(n795), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G93), .A2(n796), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G55), .A2(n799), .ZN(n800) );
  XNOR2_X1 U889 ( .A(KEYINPUT79), .B(n800), .ZN(n801) );
  NOR2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n803), .A2(G67), .ZN(n804) );
  NAND2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n815) );
  XNOR2_X1 U893 ( .A(n806), .B(n815), .ZN(G145) );
  INV_X1 U894 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U895 ( .A(G166), .B(G290), .ZN(n807) );
  XNOR2_X1 U896 ( .A(n807), .B(n815), .ZN(n810) );
  XNOR2_X1 U897 ( .A(KEYINPUT19), .B(G305), .ZN(n808) );
  XNOR2_X1 U898 ( .A(n808), .B(G288), .ZN(n809) );
  XOR2_X1 U899 ( .A(n810), .B(n809), .Z(n812) );
  XNOR2_X1 U900 ( .A(G299), .B(KEYINPUT84), .ZN(n811) );
  XNOR2_X1 U901 ( .A(n812), .B(n811), .ZN(n990) );
  XNOR2_X1 U902 ( .A(n813), .B(n990), .ZN(n814) );
  NAND2_X1 U903 ( .A1(n814), .A2(G868), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U905 ( .A1(n818), .A2(n817), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n819) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n819), .Z(n820) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n820), .ZN(n821) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G237), .A2(G236), .ZN(n823) );
  NAND2_X1 U913 ( .A1(G69), .A2(n823), .ZN(n824) );
  XNOR2_X1 U914 ( .A(KEYINPUT87), .B(n824), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G108), .ZN(n840) );
  NAND2_X1 U916 ( .A1(n840), .A2(G567), .ZN(n832) );
  XOR2_X1 U917 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n827) );
  NAND2_X1 U918 ( .A1(G132), .A2(G82), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n827), .B(n826), .ZN(n828) );
  NOR2_X1 U920 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G96), .A2(n829), .ZN(n830) );
  XNOR2_X1 U922 ( .A(KEYINPUT86), .B(n830), .ZN(n841) );
  NAND2_X1 U923 ( .A1(n841), .A2(G2106), .ZN(n831) );
  NAND2_X1 U924 ( .A1(n832), .A2(n831), .ZN(n960) );
  NAND2_X1 U925 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U926 ( .A1(n960), .A2(n833), .ZN(n839) );
  NAND2_X1 U927 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  INV_X1 U929 ( .A(G661), .ZN(n836) );
  NAND2_X1 U930 ( .A1(G2), .A2(G15), .ZN(n835) );
  NOR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U932 ( .A(KEYINPUT106), .B(n837), .Z(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U935 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n841), .A2(n840), .ZN(G325) );
  XOR2_X1 U937 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  XNOR2_X1 U938 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  NAND2_X1 U940 ( .A1(G124), .A2(n963), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n842), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n967), .A2(G100), .ZN(n843) );
  NAND2_X1 U943 ( .A1(n844), .A2(n843), .ZN(n848) );
  NAND2_X1 U944 ( .A1(n964), .A2(G112), .ZN(n846) );
  NAND2_X1 U945 ( .A1(G136), .A2(n968), .ZN(n845) );
  NAND2_X1 U946 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U947 ( .A1(n848), .A2(n847), .ZN(G162) );
  XOR2_X1 U948 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n867) );
  XNOR2_X1 U949 ( .A(G2090), .B(G35), .ZN(n862) );
  XNOR2_X1 U950 ( .A(G1996), .B(G32), .ZN(n850) );
  XNOR2_X1 U951 ( .A(G33), .B(G2072), .ZN(n849) );
  NOR2_X1 U952 ( .A1(n850), .A2(n849), .ZN(n856) );
  XOR2_X1 U953 ( .A(G2067), .B(G26), .Z(n851) );
  NAND2_X1 U954 ( .A1(n851), .A2(G28), .ZN(n854) );
  XOR2_X1 U955 ( .A(G25), .B(G1991), .Z(n852) );
  XNOR2_X1 U956 ( .A(KEYINPUT119), .B(n852), .ZN(n853) );
  NOR2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n859) );
  XNOR2_X1 U959 ( .A(G27), .B(n857), .ZN(n858) );
  NOR2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT53), .B(n860), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n865) );
  XOR2_X1 U963 ( .A(G2084), .B(G34), .Z(n863) );
  XNOR2_X1 U964 ( .A(KEYINPUT54), .B(n863), .ZN(n864) );
  NAND2_X1 U965 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n869) );
  INV_X1 U967 ( .A(G29), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G11), .A2(n870), .ZN(n905) );
  XNOR2_X1 U970 ( .A(G160), .B(G2084), .ZN(n873) );
  NOR2_X1 U971 ( .A1(n871), .A2(n961), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(KEYINPUT116), .B(n878), .Z(n883) );
  XOR2_X1 U976 ( .A(G2090), .B(G162), .Z(n879) );
  NOR2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U978 ( .A(KEYINPUT51), .B(n881), .ZN(n882) );
  NOR2_X1 U979 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U980 ( .A(KEYINPUT117), .B(n884), .Z(n896) );
  NAND2_X1 U981 ( .A1(G103), .A2(n967), .ZN(n886) );
  NAND2_X1 U982 ( .A1(G139), .A2(n968), .ZN(n885) );
  NAND2_X1 U983 ( .A1(n886), .A2(n885), .ZN(n891) );
  NAND2_X1 U984 ( .A1(G127), .A2(n963), .ZN(n888) );
  NAND2_X1 U985 ( .A1(G115), .A2(n964), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n962) );
  XOR2_X1 U989 ( .A(G2072), .B(n962), .Z(n893) );
  XOR2_X1 U990 ( .A(G164), .B(G2078), .Z(n892) );
  NOR2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U992 ( .A(KEYINPUT50), .B(n894), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n899), .B(KEYINPUT52), .ZN(n901) );
  INV_X1 U996 ( .A(KEYINPUT55), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n902), .A2(G29), .ZN(n903) );
  XOR2_X1 U999 ( .A(KEYINPUT118), .B(n903), .Z(n904) );
  NOR2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n931) );
  XOR2_X1 U1001 ( .A(n994), .B(G1341), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G166), .B(G1971), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n926) );
  XNOR2_X1 U1004 ( .A(G1966), .B(G168), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(KEYINPUT57), .B(n910), .ZN(n924) );
  XNOR2_X1 U1007 ( .A(G299), .B(n911), .ZN(n918) );
  XNOR2_X1 U1008 ( .A(KEYINPUT121), .B(n912), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n922) );
  XNOR2_X1 U1012 ( .A(n991), .B(G1348), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(G171), .B(G1961), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1016 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1017 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1018 ( .A(KEYINPUT122), .B(n927), .Z(n929) );
  XNOR2_X1 U1019 ( .A(KEYINPUT56), .B(G16), .ZN(n928) );
  NAND2_X1 U1020 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1021 ( .A1(n931), .A2(n930), .ZN(n958) );
  XOR2_X1 U1022 ( .A(G1976), .B(G23), .Z(n933) );
  XOR2_X1 U1023 ( .A(G1971), .B(G22), .Z(n932) );
  NAND2_X1 U1024 ( .A1(n933), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1025 ( .A(G24), .B(G1986), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1027 ( .A(KEYINPUT58), .B(n936), .Z(n953) );
  XOR2_X1 U1028 ( .A(G1961), .B(G5), .Z(n947) );
  XNOR2_X1 U1029 ( .A(G1348), .B(KEYINPUT59), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(n937), .B(G4), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(G1341), .B(G19), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G1956), .B(G20), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n944) );
  XOR2_X1 U1035 ( .A(KEYINPUT123), .B(G1981), .Z(n942) );
  XNOR2_X1 U1036 ( .A(G6), .B(n942), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT60), .B(n945), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(G21), .B(G1966), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(KEYINPUT124), .B(n948), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT125), .B(n951), .ZN(n952) );
  NOR2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1045 ( .A(n954), .B(KEYINPUT61), .Z(n955) );
  XNOR2_X1 U1046 ( .A(KEYINPUT126), .B(n955), .ZN(n956) );
  NOR2_X1 U1047 ( .A1(G16), .A2(n956), .ZN(n957) );
  NOR2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(n959), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1050 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1051 ( .A(G132), .ZN(G219) );
  INV_X1 U1052 ( .A(G96), .ZN(G221) );
  INV_X1 U1053 ( .A(G82), .ZN(G220) );
  INV_X1 U1054 ( .A(n960), .ZN(G319) );
  XNOR2_X1 U1055 ( .A(n962), .B(n961), .ZN(n975) );
  NAND2_X1 U1056 ( .A1(G130), .A2(n963), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(G118), .A2(n964), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n973) );
  NAND2_X1 U1059 ( .A1(G106), .A2(n967), .ZN(n970) );
  NAND2_X1 U1060 ( .A1(G142), .A2(n968), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1062 ( .A(KEYINPUT45), .B(n971), .Z(n972) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n975), .B(n974), .ZN(n983) );
  XOR2_X1 U1065 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n977) );
  XNOR2_X1 U1066 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n977), .B(n976), .ZN(n978) );
  XOR2_X1 U1068 ( .A(n978), .B(G162), .Z(n981) );
  XOR2_X1 U1069 ( .A(G164), .B(n979), .Z(n980) );
  XNOR2_X1 U1070 ( .A(n981), .B(n980), .ZN(n982) );
  XOR2_X1 U1071 ( .A(n983), .B(n982), .Z(n986) );
  XNOR2_X1 U1072 ( .A(G160), .B(n984), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(n986), .B(n985), .ZN(n987) );
  XOR2_X1 U1074 ( .A(n988), .B(n987), .Z(n989) );
  NOR2_X1 U1075 ( .A1(G37), .A2(n989), .ZN(G395) );
  XNOR2_X1 U1076 ( .A(G286), .B(n990), .ZN(n993) );
  XNOR2_X1 U1077 ( .A(G171), .B(n991), .ZN(n992) );
  XNOR2_X1 U1078 ( .A(n993), .B(n992), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(n995), .B(n994), .ZN(n996) );
  NOR2_X1 U1080 ( .A1(G37), .A2(n996), .ZN(G397) );
  XOR2_X1 U1081 ( .A(G1981), .B(G1971), .Z(n998) );
  XNOR2_X1 U1082 ( .A(G1996), .B(G1966), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n998), .B(n997), .ZN(n1002) );
  XOR2_X1 U1084 ( .A(KEYINPUT111), .B(G2474), .Z(n1000) );
  XNOR2_X1 U1085 ( .A(G1991), .B(G1956), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(n1000), .B(n999), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(n1002), .B(n1001), .Z(n1004) );
  XNOR2_X1 U1088 ( .A(G1976), .B(KEYINPUT41), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(n1004), .B(n1003), .ZN(n1006) );
  XOR2_X1 U1090 ( .A(G1986), .B(G1961), .Z(n1005) );
  XNOR2_X1 U1091 ( .A(n1006), .B(n1005), .ZN(G229) );
  XOR2_X1 U1092 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n1008) );
  XNOR2_X1 U1093 ( .A(G2072), .B(G2090), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1008), .B(n1007), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(KEYINPUT43), .B(G2678), .Z(n1010) );
  XNOR2_X1 U1096 ( .A(G2067), .B(KEYINPUT42), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1010), .B(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(n1012), .B(n1011), .Z(n1014) );
  XNOR2_X1 U1099 ( .A(G2096), .B(G2100), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1014), .B(n1013), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(G2078), .B(G2084), .Z(n1015) );
  XNOR2_X1 U1102 ( .A(n1016), .B(n1015), .ZN(G227) );
  NOR2_X1 U1103 ( .A1(G395), .A2(G397), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(n1017), .B(KEYINPUT114), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(G319), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(G401), .A2(n1019), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(G229), .A2(G227), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT49), .B(n1020), .Z(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(G225) );
  INV_X1 U1110 ( .A(G225), .ZN(G308) );
endmodule

