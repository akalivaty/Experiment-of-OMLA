//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(KEYINPUT88), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n203), .A2(new_n207), .A3(new_n208), .A4(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n213), .B(new_n212), .C1(new_n205), .C2(new_n206), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G43gat), .ZN(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G50gat), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT15), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n216), .A2(KEYINPUT89), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT89), .B1(new_n216), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n215), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n226), .B(new_n215), .C1(new_n222), .C2(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT90), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n230), .A3(G1gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G8gat), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n233), .A2(new_n239), .A3(new_n234), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT91), .B1(new_n228), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244));
  AOI211_X1 g043(.A(new_n244), .B(new_n241), .C1(new_n225), .C2(new_n227), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n224), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n246), .A2(KEYINPUT18), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n216), .A2(new_n221), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT89), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n216), .A2(KEYINPUT89), .A3(new_n221), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n226), .B1(new_n254), .B2(new_n215), .ZN(new_n255));
  INV_X1    g054(.A(new_n227), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n242), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n244), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n228), .A2(KEYINPUT91), .A3(new_n242), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n258), .A2(new_n247), .A3(new_n248), .A4(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n241), .A2(new_n224), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n263), .A2(new_n247), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n248), .B(KEYINPUT13), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G113gat), .B(G141gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(G197gat), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT11), .B(G169gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT87), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT12), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n249), .A2(new_n262), .A3(new_n273), .A4(new_n266), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G57gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT67), .ZN(new_n284));
  INV_X1    g083(.A(G127gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(G134gat), .A3(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(G127gat), .A2(G134gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n288), .B(new_n289), .C1(KEYINPUT1), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT68), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  INV_X1    g092(.A(G113gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G120gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(G120gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n289), .A4(new_n288), .ZN(new_n300));
  AND2_X1   g099(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n302));
  OAI21_X1  g101(.A(G113gat), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G127gat), .A2(G134gat), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n303), .A2(new_n295), .B1(new_n289), .B2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n306));
  AOI22_X1  g105(.A1(new_n292), .A2(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G141gat), .ZN(new_n309));
  XOR2_X1   g108(.A(KEYINPUT79), .B(G141gat), .Z(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n315), .B2(KEYINPUT2), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n319), .A2(new_n321), .B1(new_n313), .B2(new_n314), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n312), .B(new_n320), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n311), .A2(new_n316), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n307), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT81), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n292), .A2(new_n300), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n306), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n324), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n307), .A2(KEYINPUT81), .A3(new_n324), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n325), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT5), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n324), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n329), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI221_X4 g139(.A(KEYINPUT71), .B1(new_n305), .B2(new_n306), .C1(new_n292), .C2(new_n300), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n327), .B2(new_n328), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n324), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n347), .A3(new_n332), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n340), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n335), .B1(new_n349), .B2(new_n334), .ZN(new_n350));
  INV_X1    g149(.A(new_n334), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT5), .ZN(new_n352));
  INV_X1    g151(.A(new_n345), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n324), .B(new_n353), .C1(new_n341), .C2(new_n343), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n347), .B1(new_n331), .B2(new_n332), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n339), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n283), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  AOI211_X1 g159(.A(new_n351), .B(new_n340), .C1(new_n346), .C2(new_n348), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n357), .B(new_n282), .C1(new_n361), .C2(new_n335), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT82), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT6), .B(new_n283), .C1(new_n350), .C2(new_n358), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n359), .A2(new_n366), .A3(new_n360), .A4(new_n362), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G197gat), .B(G204gat), .ZN(new_n372));
  INV_X1    g171(.A(G211gat), .ZN(new_n373));
  INV_X1    g172(.A(G218gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n372), .B1(KEYINPUT22), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G211gat), .B(G218gat), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G226gat), .ZN(new_n380));
  INV_X1    g179(.A(G233gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(G183gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G183gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n387), .A3(KEYINPUT27), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n384), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(KEYINPUT66), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT66), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT65), .B(G183gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT28), .ZN(new_n395));
  INV_X1    g194(.A(G190gat), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n391), .A2(new_n394), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT26), .ZN(new_n398));
  INV_X1    g197(.A(G169gat), .ZN(new_n399));
  INV_X1    g198(.A(G176gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT27), .B(G183gat), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n395), .B1(new_n407), .B2(new_n396), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT23), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT64), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n399), .A2(new_n400), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT23), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n411), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n412), .B(new_n402), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT24), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n405), .B(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(G190gat), .B1(new_n385), .B2(new_n387), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT25), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n405), .B(KEYINPUT24), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n384), .A2(new_n396), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT25), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n417), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT64), .B1(new_n411), .B2(KEYINPUT23), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n426), .A2(new_n412), .A3(new_n429), .A4(new_n402), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n423), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT76), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n410), .A2(new_n430), .A3(new_n423), .A4(KEYINPUT76), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n383), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n382), .A2(KEYINPUT29), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n379), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n410), .A2(new_n423), .A3(new_n430), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n382), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n378), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n371), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT30), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n442), .A3(new_n371), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n446), .A2(KEYINPUT77), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n443), .A2(KEYINPUT30), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n446), .B2(KEYINPUT77), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n368), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT29), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n378), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n324), .B1(new_n452), .B2(new_n337), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n378), .B1(new_n338), .B2(new_n451), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G78gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT31), .B(G50gat), .Z(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G228gat), .A2(G233gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G22gat), .ZN(new_n461));
  INV_X1    g260(.A(G106gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n459), .B(new_n463), .Z(new_n464));
  OAI21_X1  g263(.A(new_n440), .B1(new_n343), .B2(new_n341), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OR3_X1    g266(.A1(new_n440), .A2(new_n341), .A3(new_n343), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n440), .B(KEYINPUT72), .C1(new_n343), .C2(new_n341), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(G227gat), .A2(G233gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G43gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G99gat), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT74), .B(G71gat), .Z(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT33), .B1(new_n470), .B2(new_n471), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n470), .B2(new_n471), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT73), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n475), .A2(new_n479), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n479), .A2(KEYINPUT33), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI22_X1  g286(.A1(new_n470), .A2(new_n471), .B1(KEYINPUT75), .B2(KEYINPUT34), .ZN(new_n488));
  NAND2_X1  g287(.A1(KEYINPUT75), .A2(KEYINPUT34), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n485), .B2(new_n487), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n464), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT35), .B1(new_n450), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(KEYINPUT86), .A2(KEYINPUT35), .ZN(new_n495));
  INV_X1    g294(.A(new_n448), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n444), .A3(new_n445), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n363), .B2(new_n365), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n459), .B(new_n463), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n488), .B(new_n489), .Z(new_n502));
  OAI21_X1  g301(.A(new_n479), .B1(new_n483), .B2(KEYINPUT73), .ZN(new_n503));
  AOI211_X1 g302(.A(new_n474), .B(new_n482), .C1(new_n470), .C2(new_n471), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n503), .A2(new_n480), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n487), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(KEYINPUT86), .A2(KEYINPUT35), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n363), .A2(new_n365), .ZN(new_n511));
  INV_X1    g310(.A(new_n497), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n500), .A2(new_n509), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n507), .A2(KEYINPUT36), .A3(new_n508), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT36), .B1(new_n507), .B2(new_n508), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n450), .A2(new_n501), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n339), .B1(new_n355), .B2(new_n356), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n351), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n333), .A2(new_n334), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT39), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT39), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n525), .A3(new_n351), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n526), .A2(KEYINPUT83), .A3(new_n282), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT83), .B1(new_n526), .B2(new_n282), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT40), .B(new_n524), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n531), .A2(new_n359), .A3(new_n497), .A4(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n438), .A2(new_n442), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT37), .B1(new_n438), .B2(new_n442), .ZN(new_n538));
  INV_X1    g337(.A(new_n371), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT38), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n538), .A2(new_n539), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n536), .B2(new_n535), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(KEYINPUT84), .A3(KEYINPUT38), .ZN(new_n545));
  INV_X1    g344(.A(new_n443), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n435), .A2(new_n379), .A3(new_n437), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n378), .B1(new_n439), .B2(new_n441), .ZN(new_n548));
  OR3_X1    g347(.A1(new_n547), .A2(new_n548), .A3(new_n536), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n543), .A2(new_n541), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n542), .A2(new_n545), .A3(new_n546), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n533), .B(new_n464), .C1(new_n511), .C2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n519), .A2(new_n520), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n278), .B1(new_n516), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT102), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(G71gat), .A2(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n456), .ZN(new_n564));
  NAND3_X1  g363(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT93), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n571));
  INV_X1    g370(.A(G57gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(G64gat), .ZN(new_n573));
  INV_X1    g372(.A(G64gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(G57gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(G57gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n572), .A2(G64gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT94), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n576), .A2(new_n579), .A3(new_n580), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n570), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n577), .B(KEYINPUT95), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n581), .A2(new_n582), .B1(new_n564), .B2(new_n560), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT96), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n570), .A2(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n559), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(G183gat), .B1(new_n594), .B2(new_n241), .ZN(new_n595));
  AOI221_X4 g394(.A(KEYINPUT96), .B1(new_n587), .B2(new_n586), .C1(new_n570), .C2(new_n584), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n592), .B1(new_n585), .B2(new_n588), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT21), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n384), .A3(new_n242), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n591), .A2(KEYINPUT21), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n595), .B2(new_n599), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n558), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n595), .A2(new_n599), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n607), .A2(new_n602), .A3(G231gat), .A4(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G211gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n605), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n605), .B2(new_n608), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n557), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n605), .A2(new_n608), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n610), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n605), .A2(new_n608), .A3(new_n611), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n556), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n622));
  AND2_X1   g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(G99gat), .A2(G106gat), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G99gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n462), .ZN(new_n627));
  NAND2_X1  g426(.A1(G99gat), .A2(G106gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(KEYINPUT98), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  AND2_X1   g430(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(KEYINPUT97), .A2(G92gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G85gat), .A2(G92gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT7), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT7), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(G85gat), .A3(G92gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n628), .A2(KEYINPUT8), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n634), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n630), .A2(KEYINPUT99), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n630), .A2(new_n641), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n636), .A2(new_n638), .B1(KEYINPUT8), .B2(new_n628), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n634), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n643), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n228), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n224), .ZN(new_n651));
  NAND3_X1  g450(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT100), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n657));
  NAND2_X1  g456(.A1(G232gat), .A2(G233gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n657), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n660), .B(new_n649), .C1(new_n654), .C2(new_n655), .ZN(new_n661));
  XNOR2_X1  g460(.A(G134gat), .B(G162gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT101), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n659), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n659), .B2(new_n661), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n621), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n659), .A2(new_n661), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n663), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n620), .A3(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n555), .B1(new_n619), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(new_n614), .A3(new_n618), .A4(KEYINPUT102), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G120gat), .B(G148gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(G176gat), .B(G204gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n585), .A2(new_n588), .A3(new_n643), .A4(new_n647), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n650), .B2(new_n591), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(G230gat), .A3(G233gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(G230gat), .A2(G233gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT103), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT10), .B(new_n650), .C1(new_n596), .C2(new_n597), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT10), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n688), .B(new_n680), .C1(new_n650), .C2(new_n591), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n679), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n687), .A2(new_n689), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n684), .ZN(new_n693));
  INV_X1    g492(.A(new_n679), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n682), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n676), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n554), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n368), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n232), .ZN(G1324gat));
  NAND3_X1  g500(.A1(new_n554), .A2(new_n698), .A3(new_n497), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT16), .B(G8gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT105), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n702), .B(KEYINPUT104), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n707), .B2(G8gat), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n705), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(G1325gat));
  INV_X1    g509(.A(G15gat), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n699), .A2(new_n711), .A3(new_n519), .ZN(new_n712));
  INV_X1    g511(.A(new_n699), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n491), .A2(new_n492), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n711), .B2(new_n716), .ZN(G1326gat));
  NOR2_X1   g516(.A1(new_n699), .A2(new_n464), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  AOI21_X1  g519(.A(new_n674), .B1(new_n516), .B2(new_n553), .ZN(new_n721));
  INV_X1    g520(.A(new_n619), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n696), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n277), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n368), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n210), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n516), .A2(new_n553), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n672), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n721), .A2(KEYINPUT44), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n275), .A2(KEYINPUT106), .A3(new_n276), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT106), .B1(new_n275), .B2(new_n276), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n731), .A2(new_n723), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n368), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n727), .A2(new_n738), .ZN(G1328gat));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n211), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT46), .B1(new_n740), .B2(new_n512), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n737), .B2(new_n512), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n740), .A2(KEYINPUT46), .A3(new_n512), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n740), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n512), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n741), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(G1329gat));
  OAI21_X1  g546(.A(G43gat), .B1(new_n737), .B2(new_n519), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n724), .A2(new_n219), .A3(new_n715), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1330gat));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT48), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n721), .A2(new_n277), .A3(new_n723), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n217), .B1(new_n756), .B2(new_n464), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n501), .A2(G50gat), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n755), .B(new_n757), .C1(new_n737), .C2(new_n758), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n754), .A2(KEYINPUT48), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n736), .A2(new_n697), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n728), .A2(new_n676), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n728), .A2(KEYINPUT109), .A3(new_n676), .A4(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n368), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n572), .ZN(G1332gat));
  NOR2_X1   g568(.A1(new_n767), .A2(new_n512), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  AND2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n770), .B2(new_n771), .ZN(G1333gat));
  OAI21_X1  g573(.A(G71gat), .B1(new_n767), .B2(new_n519), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n765), .A2(new_n563), .A3(new_n715), .A4(new_n766), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n767), .A2(new_n464), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n456), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n722), .A2(new_n736), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n731), .A2(new_n696), .A3(new_n732), .A4(new_n783), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n784), .A2(new_n631), .A3(new_n368), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n728), .A2(new_n672), .A3(new_n788), .A4(new_n783), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n790), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n721), .A2(new_n792), .A3(new_n788), .A4(new_n783), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n791), .A2(new_n725), .A3(new_n696), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n785), .B1(new_n631), .B2(new_n794), .ZN(G1336gat));
  NOR2_X1   g594(.A1(new_n632), .A2(new_n633), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n784), .B2(new_n512), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n791), .A2(new_n793), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n512), .A2(G92gat), .A3(new_n697), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n800), .B(KEYINPUT111), .Z(new_n802));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n721), .B(new_n730), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n804), .A2(new_n696), .A3(new_n497), .A4(new_n783), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n805), .B2(new_n796), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n801), .B1(new_n806), .B2(new_n798), .ZN(G1337gat));
  OAI21_X1  g606(.A(G99gat), .B1(new_n784), .B2(new_n519), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n714), .A2(G99gat), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n791), .A2(new_n696), .A3(new_n793), .A4(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n808), .B2(new_n811), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(G1338gat));
  NAND4_X1  g613(.A1(new_n791), .A2(new_n696), .A3(new_n501), .A4(new_n793), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n462), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n464), .A2(new_n462), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n804), .A2(new_n696), .A3(new_n783), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n818), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1339gat));
  NAND4_X1  g622(.A1(new_n673), .A2(new_n675), .A3(new_n697), .A4(new_n735), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n248), .B1(new_n246), .B2(new_n247), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n263), .A2(new_n247), .A3(new_n265), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT115), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n271), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n276), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n829), .B1(new_n668), .B2(new_n671), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n687), .A2(new_n689), .A3(new_n686), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n693), .A2(KEYINPUT54), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n694), .B1(new_n690), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(KEYINPUT55), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n695), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT113), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n834), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n835), .A2(new_n841), .A3(new_n695), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT114), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n837), .A2(new_n845), .A3(new_n840), .A4(new_n842), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n276), .A2(new_n828), .A3(new_n696), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n846), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n735), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(new_n674), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n824), .B1(new_n852), .B2(new_n722), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n509), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n368), .A2(new_n497), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT116), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n294), .A3(new_n736), .ZN(new_n858));
  OAI21_X1  g657(.A(G113gat), .B1(new_n856), .B2(new_n278), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1340gat));
  OR2_X1    g659(.A1(new_n301), .A2(new_n302), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n857), .A2(new_n861), .A3(new_n696), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n696), .A3(new_n855), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n863), .A2(new_n864), .A3(G120gat), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n863), .B2(G120gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(G1341gat));
  NOR2_X1   g666(.A1(new_n856), .A2(new_n619), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n286), .A2(new_n287), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n868), .B(new_n869), .ZN(G1342gat));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n672), .A3(new_n855), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT56), .B1(new_n871), .B2(G134gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(G134gat), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n871), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR4_X1   g675(.A1(new_n871), .A2(KEYINPUT118), .A3(KEYINPUT56), .A4(G134gat), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n872), .B(new_n873), .C1(new_n876), .C2(new_n877), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n853), .A2(new_n501), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n836), .ZN(new_n882));
  XOR2_X1   g681(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n883));
  NAND2_X1  g682(.A1(new_n838), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n277), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n849), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n885), .B2(new_n849), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n674), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n722), .B1(new_n888), .B2(new_n847), .ZN(new_n889));
  AND4_X1   g688(.A1(new_n673), .A2(new_n675), .A3(new_n697), .A4(new_n735), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT57), .B(new_n501), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n885), .A2(new_n849), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n849), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n672), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n619), .B1(new_n898), .B2(new_n848), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n824), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n900), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n501), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n893), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n519), .A2(new_n855), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT119), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n277), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n310), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n853), .A2(new_n501), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n903), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(G141gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT58), .B1(new_n909), .B2(new_n277), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n908), .A2(G141gat), .A3(new_n278), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n902), .A2(new_n736), .A3(new_n904), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n310), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n911), .B1(new_n912), .B2(new_n915), .ZN(G1344gat));
  OAI21_X1  g715(.A(KEYINPUT59), .B1(new_n908), .B2(new_n697), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n308), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n904), .A2(new_n696), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(KEYINPUT59), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n902), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n879), .A2(KEYINPUT57), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n676), .A2(new_n697), .A3(new_n278), .ZN(new_n923));
  INV_X1    g722(.A(new_n843), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n830), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n722), .B1(new_n888), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n880), .B(new_n501), .C1(new_n923), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT59), .B(G148gat), .C1(new_n928), .C2(new_n919), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n921), .A3(new_n929), .ZN(G1345gat));
  INV_X1    g729(.A(new_n908), .ZN(new_n931));
  AOI21_X1  g730(.A(G155gat), .B1(new_n931), .B2(new_n722), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n902), .A2(new_n904), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n619), .A2(new_n313), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G1346gat));
  AOI21_X1  g734(.A(G162gat), .B1(new_n931), .B2(new_n672), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n674), .A2(new_n314), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n933), .B2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n725), .A2(new_n512), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n854), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n399), .A3(new_n736), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(new_n277), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n399), .ZN(G1348gat));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n696), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g744(.A1(new_n940), .A2(new_n722), .A3(new_n407), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n854), .A2(new_n722), .A3(new_n939), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n393), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n854), .A2(new_n672), .A3(new_n939), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G190gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(KEYINPUT61), .A3(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(KEYINPUT123), .A3(new_n960), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n959), .B(new_n961), .C1(G190gat), .C2(new_n954), .ZN(G1351gat));
  XNOR2_X1  g761(.A(KEYINPUT124), .B(G197gat), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n519), .A2(new_n939), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n922), .A2(new_n927), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n965), .B2(new_n278), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n907), .A2(new_n964), .ZN(new_n967));
  INV_X1    g766(.A(new_n963), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n736), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1352gat));
  INV_X1    g769(.A(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n971), .A3(new_n696), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G204gat), .B1(new_n965), .B2(new_n697), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT62), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(G1353gat));
  NAND4_X1  g779(.A1(new_n922), .A2(new_n927), .A3(new_n722), .A4(new_n964), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G211gat), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT63), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n983), .A2(KEYINPUT63), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(KEYINPUT63), .ZN(new_n986));
  NAND4_X1  g785(.A1(new_n981), .A2(G211gat), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n967), .A2(new_n373), .A3(new_n722), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(G1354gat));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n965), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n672), .B1(new_n965), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g791(.A(G218gat), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n967), .A2(new_n374), .A3(new_n672), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1355gat));
endmodule


