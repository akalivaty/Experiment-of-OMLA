//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n435, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(new_n435));
  INV_X1    g010(.A(new_n435), .ZN(G219));
  XOR2_X1   g011(.A(KEYINPUT0), .B(G82), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n435), .A2(new_n437), .A3(G44), .A4(G96), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  OR2_X1    g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n454), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n470), .B1(new_n464), .B2(new_n465), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT66), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n479));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n463), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n482), .B1(new_n483), .B2(G136), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n479), .A2(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n464), .B2(new_n465), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n465), .C2(new_n464), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  OR2_X1    g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT67), .A3(G62), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT67), .B1(new_n501), .B2(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(G651), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n499), .A2(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(G88), .B1(new_n513), .B2(G50), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n508), .A2(new_n514), .ZN(G166));
  XOR2_X1   g090(.A(KEYINPUT69), .B(KEYINPUT7), .Z(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(G51), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(G89), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n518), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n510), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(G543), .B1(new_n527), .B2(new_n528), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n526), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n525), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n531), .A2(new_n539), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n513), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n529), .A2(new_n530), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G651), .B1(new_n511), .B2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(G299));
  INV_X1    g130(.A(G171), .ZN(G301));
  NAND2_X1  g131(.A1(new_n508), .A2(new_n514), .ZN(G303));
  NAND2_X1  g132(.A1(new_n511), .A2(G87), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n513), .A2(G49), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G288));
  AOI22_X1  g137(.A1(new_n511), .A2(G86), .B1(new_n513), .B2(G48), .ZN(new_n563));
  OAI21_X1  g138(.A(G61), .B1(new_n529), .B2(new_n530), .ZN(new_n564));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n525), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(new_n567), .A3(KEYINPUT70), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  INV_X1    g145(.A(G48), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n531), .A2(new_n570), .B1(new_n533), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n569), .B1(new_n572), .B2(new_n566), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G305));
  NAND2_X1  g150(.A1(new_n501), .A2(G60), .ZN(new_n576));
  NAND2_X1  g151(.A1(G72), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n525), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(KEYINPUT71), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(KEYINPUT71), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n511), .A2(G85), .B1(new_n513), .B2(G47), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT72), .Z(new_n584));
  OAI21_X1  g159(.A(G66), .B1(new_n529), .B2(new_n530), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n525), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(G54), .B(G543), .C1(new_n527), .C2(new_n528), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT73), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT73), .ZN(new_n591));
  INV_X1    g166(.A(new_n586), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n501), .B2(G66), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n588), .C1(new_n593), .C2(new_n525), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n511), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n531), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n595), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n596), .B1(new_n595), .B2(new_n601), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n584), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n584), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g191(.A(KEYINPUT3), .B(G2104), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n473), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  AOI22_X1  g196(.A1(G123), .A2(new_n482), .B1(new_n483), .B2(G135), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(KEYINPUT76), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(KEYINPUT76), .ZN(new_n625));
  OR3_X1    g200(.A1(new_n463), .A2(KEYINPUT75), .A3(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT75), .B1(new_n463), .B2(G111), .ZN(new_n627));
  NAND4_X1  g202(.A1(new_n624), .A2(new_n625), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT77), .B(G2096), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n621), .A2(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT78), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2096), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1991), .B(G1996), .Z(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(KEYINPUT79), .ZN(new_n666));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(KEYINPUT79), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n663), .A2(new_n664), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(new_n665), .ZN(new_n673));
  MUX2_X1   g248(.A(new_n673), .B(new_n672), .S(new_n668), .Z(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n675), .B1(new_n671), .B2(new_n674), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n662), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n678), .ZN(new_n680));
  INV_X1    g255(.A(new_n662), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(new_n676), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n682), .A3(new_n684), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n690));
  NOR2_X1   g265(.A1(G16), .A2(G24), .ZN(new_n691));
  XNOR2_X1  g266(.A(G290), .B(KEYINPUT83), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT84), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  INV_X1    g273(.A(G107), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G2105), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n617), .A2(G2105), .ZN(new_n701));
  INV_X1    g276(.A(G119), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT81), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n482), .A2(new_n704), .A3(G119), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n700), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n617), .A2(G131), .A3(new_n463), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT80), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT82), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n706), .B2(new_n708), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n697), .B1(new_n712), .B2(new_n696), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XOR2_X1   g289(.A(new_n713), .B(new_n714), .Z(new_n715));
  NOR2_X1   g290(.A1(new_n695), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT86), .Z(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n721), .ZN(new_n724));
  NOR2_X1   g299(.A1(G6), .A2(G16), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n574), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT32), .B(G1981), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT85), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n717), .A2(G23), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n561), .B2(new_n717), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT33), .B(G1976), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n716), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n722), .A2(new_n724), .A3(new_n734), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(KEYINPUT34), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n690), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(new_n690), .A3(new_n738), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n696), .A2(G32), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  INV_X1    g319(.A(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n701), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n483), .A2(G141), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n473), .A2(G105), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n742), .B1(new_n750), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n696), .B1(KEYINPUT24), .B2(G34), .ZN(new_n755));
  OAI22_X1  g330(.A1(G160), .A2(new_n696), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  NOR2_X1   g332(.A1(G171), .A2(new_n717), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G5), .B2(new_n717), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n753), .B1(G2084), .B2(new_n756), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n696), .A2(G35), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT94), .Z(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n696), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n760), .B1(new_n764), .B2(G2090), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n751), .A2(new_n752), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT31), .B(G11), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT93), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n629), .A2(new_n696), .ZN(new_n769));
  INV_X1    g344(.A(G28), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(KEYINPUT30), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n768), .B(new_n769), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n756), .A2(G2084), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n759), .A2(new_n757), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n766), .A2(new_n773), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n717), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n717), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1966), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n696), .A2(G27), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n696), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2078), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n776), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n717), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n542), .B2(new_n717), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT88), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT87), .B(G1341), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n765), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n717), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT23), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n608), .B2(new_n717), .ZN(new_n792));
  INV_X1    g367(.A(G1956), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n764), .B2(G2090), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n696), .A2(G33), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT25), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G139), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n617), .A2(new_n463), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n617), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n463), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n796), .B1(new_n805), .B2(new_n696), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT92), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2072), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n789), .A2(new_n795), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n717), .A2(G4), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n604), .B2(new_n717), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n696), .A2(G26), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT28), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n483), .A2(G140), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n482), .A2(G128), .ZN(new_n817));
  OR2_X1    g392(.A1(G104), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT89), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT89), .A4(new_n819), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n824), .A2(KEYINPUT90), .A3(G29), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT90), .B1(new_n824), .B2(G29), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n815), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT91), .B(G2067), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n813), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT95), .B1(new_n809), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n795), .A2(new_n808), .ZN(new_n832));
  OR4_X1    g407(.A1(KEYINPUT95), .A2(new_n789), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n740), .A2(new_n741), .B1(new_n831), .B2(new_n833), .ZN(G311));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n833), .ZN(new_n835));
  INV_X1    g410(.A(new_n741), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n739), .B2(new_n836), .ZN(G150));
  AOI22_X1  g412(.A1(new_n501), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n525), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n531), .A2(new_n840), .B1(new_n533), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n844), .B(new_n845), .C1(new_n538), .C2(new_n541), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(KEYINPUT96), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n839), .B2(new_n842), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n542), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n604), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n844), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(G145));
  XNOR2_X1  g434(.A(new_n629), .B(G160), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G162), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n710), .A2(new_n711), .ZN(new_n863));
  INV_X1    g438(.A(new_n619), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n866));
  INV_X1    g441(.A(G130), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n701), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n482), .A2(KEYINPUT97), .A3(G130), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  INV_X1    g446(.A(G118), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(G2105), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n483), .B2(G142), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n865), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n870), .A2(new_n865), .A3(new_n874), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n864), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n879), .A2(new_n619), .A3(new_n875), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n863), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n619), .B1(new_n879), .B2(new_n875), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n876), .A2(new_n864), .A3(new_n877), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n712), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(G164), .B1(new_n822), .B2(new_n823), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n822), .A2(G164), .A3(new_n823), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n750), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n750), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  OAI22_X1  g466(.A1(new_n890), .A2(new_n891), .B1(new_n804), .B2(new_n802), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n805), .A3(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n885), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n894), .ZN(new_n898));
  INV_X1    g473(.A(new_n885), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n899), .A3(new_n896), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n862), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n895), .A2(new_n862), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n885), .B1(new_n894), .B2(new_n892), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT100), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n896), .B2(new_n895), .ZN(new_n909));
  INV_X1    g484(.A(new_n902), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n861), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  INV_X1    g487(.A(new_n907), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n908), .A2(new_n914), .A3(KEYINPUT40), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n908), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(G395));
  XNOR2_X1  g492(.A(new_n613), .B(KEYINPUT101), .ZN(new_n918));
  INV_X1    g493(.A(new_n850), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n613), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n850), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n595), .A2(new_n601), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n925), .A2(G299), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(G299), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT41), .B1(new_n926), .B2(new_n927), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(KEYINPUT102), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n928), .A2(new_n935), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n920), .A2(new_n923), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(G305), .A2(G290), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G305), .A2(G290), .ZN(new_n941));
  NAND2_X1  g516(.A1(G166), .A2(G288), .ZN(new_n942));
  NAND2_X1  g517(.A1(G303), .A2(new_n561), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n940), .A2(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n943), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n945), .A2(new_n946), .A3(new_n939), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT42), .Z(new_n949));
  AND3_X1   g524(.A1(new_n930), .A2(new_n938), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n930), .B2(new_n938), .ZN(new_n951));
  OAI21_X1  g526(.A(G868), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g528(.A(new_n952), .B1(G868), .B2(new_n843), .ZN(G331));
  NAND2_X1  g529(.A1(G171), .A2(KEYINPUT103), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n526), .B2(new_n535), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(G286), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(G286), .A2(new_n958), .A3(new_n956), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n961), .ZN(new_n963));
  INV_X1    g538(.A(new_n955), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n963), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n850), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(new_n961), .A3(new_n955), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n964), .B1(new_n963), .B2(new_n959), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n919), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n928), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n934), .A2(new_n966), .A3(new_n936), .A4(new_n969), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n948), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n904), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n944), .B2(new_n947), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n940), .A2(new_n942), .A3(new_n943), .A4(new_n941), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n946), .B1(new_n945), .B2(new_n939), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT105), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n972), .B2(new_n971), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n980), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n970), .B1(new_n932), .B2(new_n933), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n929), .B1(new_n966), .B2(new_n969), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n904), .A4(new_n973), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n974), .B2(new_n981), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n986), .A2(KEYINPUT43), .A3(new_n904), .A4(new_n973), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  MUX2_X1   g567(.A(new_n989), .B(new_n992), .S(KEYINPUT44), .Z(G397));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n549), .A2(new_n994), .A3(new_n554), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n549), .B2(new_n554), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n998));
  INV_X1    g573(.A(G125), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n480), .B2(new_n481), .ZN(new_n1000));
  INV_X1    g575(.A(new_n467), .ZN(new_n1001));
  OAI21_X1  g576(.A(G2105), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n617), .A2(new_n470), .B1(G101), .B2(new_n473), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1002), .A2(KEYINPUT106), .A3(G40), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n468), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  INV_X1    g585(.A(new_n497), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n496), .B1(new_n617), .B2(new_n493), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1009), .B(new_n1010), .C1(new_n1013), .C2(new_n491), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n998), .A2(new_n1008), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n793), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(G164), .B2(G1384), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT45), .B(new_n1010), .C1(new_n1013), .C2(new_n491), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1008), .A3(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT56), .B(G2072), .Z(new_n1021));
  OAI211_X1 g596(.A(new_n997), .B(new_n1016), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1015), .A2(new_n812), .ZN(new_n1023));
  INV_X1    g598(.A(G2067), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n495), .A2(new_n497), .ZN(new_n1025));
  INV_X1    g600(.A(new_n491), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1384), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1008), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(new_n604), .A3(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n995), .A2(new_n996), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1010), .B1(new_n1013), .B2(new_n491), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1032), .A2(KEYINPUT50), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1956), .B1(new_n1033), .B2(new_n1014), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1022), .A3(KEYINPUT61), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1036), .A2(new_n1022), .A3(KEYINPUT116), .A4(KEYINPUT61), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1008), .A2(new_n1027), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT58), .B(G1341), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n1044), .A2(new_n1045), .B1(new_n1020), .B2(G1996), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n542), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(KEYINPUT59), .A3(new_n542), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT61), .B1(new_n1036), .B2(new_n1022), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1042), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT60), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n602), .A2(new_n603), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT60), .A3(new_n1023), .A4(new_n1028), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT117), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1023), .A2(KEYINPUT60), .A3(new_n1028), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1059), .A2(KEYINPUT118), .A3(new_n604), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT118), .B1(new_n1059), .B2(new_n604), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1055), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1037), .B1(new_n1054), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1015), .A2(new_n757), .ZN(new_n1066));
  INV_X1    g641(.A(G2078), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1018), .A2(new_n1019), .A3(new_n1008), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT53), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1065), .B(new_n1066), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1068), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT121), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1068), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1073), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT119), .A3(new_n1067), .A4(new_n1008), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(KEYINPUT53), .A3(new_n1070), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1065), .B1(new_n1083), .B2(new_n1066), .ZN(new_n1084));
  OAI21_X1  g659(.A(G301), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1003), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n475), .A2(KEYINPUT122), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(G40), .A4(new_n1002), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT123), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1002), .A2(G40), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1074), .A2(G2078), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1090), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1095), .A2(new_n1081), .B1(new_n757), .B2(new_n1015), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1077), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1068), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT124), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1079), .A2(new_n1101), .A3(new_n1096), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(G171), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1085), .A2(new_n1103), .A3(KEYINPUT54), .ZN(new_n1104));
  OAI21_X1  g679(.A(G171), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1099), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT54), .B1(new_n1106), .B2(G301), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G303), .A2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT109), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G8), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1020), .A2(new_n721), .ZN(new_n1118));
  INV_X1    g693(.A(G2090), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n998), .A2(new_n1014), .A3(new_n1008), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1112), .A2(KEYINPUT109), .A3(new_n1113), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1116), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT49), .ZN(new_n1124));
  INV_X1    g699(.A(G1981), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n563), .B2(new_n567), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n572), .A2(new_n566), .A3(G1981), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n563), .A2(new_n567), .A3(new_n1125), .ZN(new_n1129));
  OAI21_X1  g704(.A(G1981), .B1(new_n572), .B2(new_n566), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(KEYINPUT49), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1128), .A2(new_n1043), .A3(G8), .A4(new_n1131), .ZN(new_n1132));
  AOI221_X4 g707(.A(new_n1117), .B1(new_n561), .B2(G1976), .C1(new_n1008), .C2(new_n1027), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n561), .A2(G1976), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(G8), .A3(new_n1043), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT110), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1133), .A2(KEYINPUT110), .A3(new_n1137), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G8), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT112), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT112), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1121), .A2(new_n1148), .A3(new_n1114), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1123), .B(new_n1143), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1966), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1020), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(G2084), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n998), .A2(new_n1014), .A3(new_n1008), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(G168), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(G8), .ZN(new_n1156));
  AOI21_X1  g731(.A(G168), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT51), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(new_n1159), .A3(G8), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1150), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1064), .A2(new_n1109), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1132), .A2(new_n1136), .A3(new_n561), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1129), .B(KEYINPUT111), .ZN(new_n1164));
  OAI211_X1 g739(.A(G8), .B(new_n1043), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1143), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1123), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1158), .A2(new_n1160), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1158), .B2(new_n1160), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1169), .A2(new_n1170), .A3(new_n1150), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1105), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1167), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1148), .B1(new_n1121), .B2(new_n1114), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n998), .A2(new_n1008), .A3(new_n1014), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1175), .A2(new_n1119), .B1(new_n1020), .B2(new_n721), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1146), .B(KEYINPUT112), .C1(new_n1176), .C2(new_n1117), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1175), .A2(new_n1153), .B1(new_n1020), .B2(new_n1151), .ZN(new_n1179));
  NOR2_X1   g754(.A1(G286), .A2(new_n1117), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT113), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT113), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1180), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1178), .A2(new_n1123), .A3(new_n1186), .A4(new_n1143), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT114), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT114), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1187), .A2(new_n1191), .A3(new_n1188), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1114), .B1(new_n1121), .B2(KEYINPUT115), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1193), .B1(KEYINPUT115), .B2(new_n1121), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1188), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1194), .A2(new_n1195), .A3(new_n1123), .A4(new_n1143), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1190), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1162), .A2(new_n1173), .A3(new_n1197), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1018), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n824), .B(new_n1024), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n1201), .A2(KEYINPUT108), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(KEYINPUT108), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n750), .B(G1996), .Z(new_n1204));
  NAND3_X1  g779(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n712), .B(new_n714), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(G290), .ZN(new_n1208));
  INV_X1    g783(.A(G1986), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT107), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1211), .B1(new_n1209), .B2(new_n1208), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1200), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1198), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1200), .B1(new_n1215), .B2(new_n750), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1199), .A2(new_n1018), .A3(G1996), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT46), .Z(new_n1218));
  NAND2_X1  g793(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1219), .B(KEYINPUT47), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n712), .A2(new_n714), .ZN(new_n1221));
  XOR2_X1   g796(.A(new_n1221), .B(KEYINPUT125), .Z(new_n1222));
  OAI22_X1  g797(.A1(new_n1222), .A2(new_n1205), .B1(G2067), .B2(new_n824), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1223), .A2(new_n1200), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1220), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1207), .A2(new_n1200), .ZN(new_n1226));
  XOR2_X1   g801(.A(new_n1226), .B(KEYINPUT126), .Z(new_n1227));
  NOR3_X1   g802(.A1(new_n1211), .A2(new_n1199), .A3(new_n1018), .ZN(new_n1228));
  XOR2_X1   g803(.A(new_n1228), .B(KEYINPUT48), .Z(new_n1229));
  AOI21_X1  g804(.A(new_n1225), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1214), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n1233));
  NOR2_X1   g807(.A1(G227), .A2(new_n461), .ZN(new_n1234));
  OAI21_X1  g808(.A(new_n1234), .B1(new_n647), .B2(new_n646), .ZN(new_n1235));
  INV_X1    g809(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1233), .B1(new_n688), .B2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g811(.A(KEYINPUT127), .B(new_n1235), .C1(new_n686), .C2(new_n687), .ZN(new_n1238));
  NOR2_X1   g812(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g813(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g814(.A1(new_n908), .A2(new_n914), .ZN(new_n1241));
  AND3_X1   g815(.A1(new_n1240), .A2(new_n1241), .A3(new_n989), .ZN(G308));
  NAND3_X1  g816(.A1(new_n1240), .A2(new_n1241), .A3(new_n989), .ZN(G225));
endmodule


