

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U547 ( .A(n517), .B(n516), .ZN(n529) );
  NOR2_X1 U548 ( .A1(n741), .A2(n723), .ZN(n515) );
  NOR2_X2 U549 ( .A1(G2105), .A2(n521), .ZN(n892) );
  XNOR2_X1 U550 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n757) );
  XNOR2_X1 U551 ( .A(n758), .B(n757), .ZN(G329) );
  XNOR2_X1 U552 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n517) );
  NOR2_X1 U553 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  NAND2_X1 U554 ( .A1(n529), .A2(G137), .ZN(n519) );
  AND2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U556 ( .A1(n888), .A2(G113), .ZN(n518) );
  NAND2_X1 U557 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U558 ( .A(n520), .B(KEYINPUT68), .ZN(n527) );
  INV_X1 U559 ( .A(G2104), .ZN(n521) );
  AND2_X1 U560 ( .A1(n521), .A2(G2105), .ZN(n889) );
  NAND2_X1 U561 ( .A1(n889), .A2(G125), .ZN(n525) );
  XNOR2_X1 U562 ( .A(KEYINPUT23), .B(KEYINPUT66), .ZN(n523) );
  NAND2_X1 U563 ( .A1(n892), .A2(G101), .ZN(n522) );
  XOR2_X1 U564 ( .A(n523), .B(n522), .Z(n524) );
  NAND2_X1 U565 ( .A1(n525), .A2(n524), .ZN(n526) );
  OR2_X1 U566 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X2 U567 ( .A(n528), .B(KEYINPUT65), .ZN(G160) );
  NAND2_X1 U568 ( .A1(G138), .A2(n529), .ZN(n531) );
  NAND2_X1 U569 ( .A1(G126), .A2(n889), .ZN(n530) );
  NAND2_X1 U570 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U571 ( .A1(G114), .A2(n888), .ZN(n533) );
  NAND2_X1 U572 ( .A1(G102), .A2(n892), .ZN(n532) );
  NAND2_X1 U573 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U574 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U575 ( .A(KEYINPUT93), .B(n536), .Z(G164) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n587) );
  INV_X1 U577 ( .A(G651), .ZN(n541) );
  NOR2_X1 U578 ( .A1(n587), .A2(n541), .ZN(n801) );
  NAND2_X1 U579 ( .A1(G72), .A2(n801), .ZN(n538) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n802) );
  NAND2_X1 U581 ( .A1(G85), .A2(n802), .ZN(n537) );
  NAND2_X1 U582 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U583 ( .A(KEYINPUT69), .B(n539), .ZN(n546) );
  NOR2_X1 U584 ( .A1(G651), .A2(n587), .ZN(n540) );
  XNOR2_X1 U585 ( .A(KEYINPUT64), .B(n540), .ZN(n798) );
  NAND2_X1 U586 ( .A1(n798), .A2(G47), .ZN(n544) );
  NOR2_X1 U587 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n542), .Z(n797) );
  NAND2_X1 U589 ( .A1(G60), .A2(n797), .ZN(n543) );
  AND2_X1 U590 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U591 ( .A1(n546), .A2(n545), .ZN(G290) );
  NAND2_X1 U592 ( .A1(n802), .A2(G89), .ZN(n547) );
  XNOR2_X1 U593 ( .A(n547), .B(KEYINPUT4), .ZN(n549) );
  NAND2_X1 U594 ( .A1(G76), .A2(n801), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U596 ( .A(KEYINPUT5), .B(n550), .ZN(n558) );
  NAND2_X1 U597 ( .A1(G63), .A2(n797), .ZN(n553) );
  NAND2_X1 U598 ( .A1(G51), .A2(n798), .ZN(n551) );
  XOR2_X1 U599 ( .A(KEYINPUT79), .B(n551), .Z(n552) );
  NAND2_X1 U600 ( .A1(n553), .A2(n552), .ZN(n556) );
  XNOR2_X1 U601 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n554) );
  XNOR2_X1 U602 ( .A(n554), .B(KEYINPUT6), .ZN(n555) );
  XNOR2_X1 U603 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U604 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U605 ( .A(KEYINPUT7), .B(n559), .ZN(G168) );
  XNOR2_X1 U606 ( .A(KEYINPUT71), .B(KEYINPUT9), .ZN(n563) );
  NAND2_X1 U607 ( .A1(G77), .A2(n801), .ZN(n561) );
  NAND2_X1 U608 ( .A1(G90), .A2(n802), .ZN(n560) );
  NAND2_X1 U609 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U610 ( .A(n563), .B(n562), .ZN(n568) );
  NAND2_X1 U611 ( .A1(G52), .A2(n798), .ZN(n564) );
  XNOR2_X1 U612 ( .A(n564), .B(KEYINPUT70), .ZN(n566) );
  NAND2_X1 U613 ( .A1(G64), .A2(n797), .ZN(n565) );
  NAND2_X1 U614 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U615 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U616 ( .A(KEYINPUT72), .B(n569), .ZN(G171) );
  NAND2_X1 U617 ( .A1(G75), .A2(n801), .ZN(n571) );
  NAND2_X1 U618 ( .A1(G88), .A2(n802), .ZN(n570) );
  NAND2_X1 U619 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U620 ( .A1(G62), .A2(n797), .ZN(n573) );
  NAND2_X1 U621 ( .A1(G50), .A2(n798), .ZN(n572) );
  NAND2_X1 U622 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U623 ( .A1(n575), .A2(n574), .ZN(G166) );
  INV_X1 U624 ( .A(G166), .ZN(G303) );
  NAND2_X1 U625 ( .A1(G65), .A2(n797), .ZN(n576) );
  XNOR2_X1 U626 ( .A(n576), .B(KEYINPUT74), .ZN(n583) );
  NAND2_X1 U627 ( .A1(G78), .A2(n801), .ZN(n578) );
  NAND2_X1 U628 ( .A1(G91), .A2(n802), .ZN(n577) );
  NAND2_X1 U629 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U630 ( .A1(G53), .A2(n798), .ZN(n579) );
  XNOR2_X1 U631 ( .A(KEYINPUT75), .B(n579), .ZN(n580) );
  NOR2_X1 U632 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U633 ( .A1(n583), .A2(n582), .ZN(G299) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G651), .A2(G74), .ZN(n585) );
  NAND2_X1 U636 ( .A1(G49), .A2(n798), .ZN(n584) );
  NAND2_X1 U637 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U638 ( .A1(n797), .A2(n586), .ZN(n589) );
  NAND2_X1 U639 ( .A1(n587), .A2(G87), .ZN(n588) );
  NAND2_X1 U640 ( .A1(n589), .A2(n588), .ZN(G288) );
  NAND2_X1 U641 ( .A1(n801), .A2(G73), .ZN(n590) );
  XNOR2_X1 U642 ( .A(n590), .B(KEYINPUT2), .ZN(n592) );
  NAND2_X1 U643 ( .A1(G61), .A2(n797), .ZN(n591) );
  NAND2_X1 U644 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U645 ( .A1(G86), .A2(n802), .ZN(n593) );
  XNOR2_X1 U646 ( .A(KEYINPUT87), .B(n593), .ZN(n594) );
  NOR2_X1 U647 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U648 ( .A(KEYINPUT88), .B(n596), .ZN(n598) );
  NAND2_X1 U649 ( .A1(n798), .A2(G48), .ZN(n597) );
  NAND2_X1 U650 ( .A1(n598), .A2(n597), .ZN(G305) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n641) );
  INV_X1 U652 ( .A(KEYINPUT94), .ZN(n600) );
  NAND2_X1 U653 ( .A1(G40), .A2(G160), .ZN(n599) );
  XNOR2_X1 U654 ( .A(n600), .B(n599), .ZN(n640) );
  INV_X1 U655 ( .A(n640), .ZN(n601) );
  NOR2_X1 U656 ( .A1(n641), .A2(n601), .ZN(n602) );
  XNOR2_X1 U657 ( .A(n602), .B(KEYINPUT95), .ZN(n749) );
  NAND2_X1 U658 ( .A1(G116), .A2(n888), .ZN(n604) );
  NAND2_X1 U659 ( .A1(G128), .A2(n889), .ZN(n603) );
  NAND2_X1 U660 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U661 ( .A(KEYINPUT35), .B(n605), .ZN(n611) );
  NAND2_X1 U662 ( .A1(n529), .A2(G140), .ZN(n606) );
  XNOR2_X1 U663 ( .A(n606), .B(KEYINPUT96), .ZN(n608) );
  NAND2_X1 U664 ( .A1(G104), .A2(n892), .ZN(n607) );
  NAND2_X1 U665 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U666 ( .A(KEYINPUT34), .B(n609), .Z(n610) );
  NAND2_X1 U667 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U668 ( .A(KEYINPUT36), .B(n612), .Z(n885) );
  XNOR2_X1 U669 ( .A(G2067), .B(KEYINPUT37), .ZN(n613) );
  AND2_X1 U670 ( .A1(n885), .A2(n613), .ZN(n985) );
  NOR2_X1 U671 ( .A1(n885), .A2(n613), .ZN(n986) );
  NAND2_X1 U672 ( .A1(G105), .A2(n892), .ZN(n614) );
  XNOR2_X1 U673 ( .A(n614), .B(KEYINPUT38), .ZN(n621) );
  NAND2_X1 U674 ( .A1(G141), .A2(n529), .ZN(n616) );
  NAND2_X1 U675 ( .A1(G129), .A2(n889), .ZN(n615) );
  NAND2_X1 U676 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U677 ( .A1(n888), .A2(G117), .ZN(n617) );
  XOR2_X1 U678 ( .A(KEYINPUT98), .B(n617), .Z(n618) );
  NOR2_X1 U679 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U680 ( .A1(n621), .A2(n620), .ZN(n883) );
  NOR2_X1 U681 ( .A1(G1996), .A2(n883), .ZN(n977) );
  NAND2_X1 U682 ( .A1(G131), .A2(n529), .ZN(n623) );
  NAND2_X1 U683 ( .A1(G119), .A2(n889), .ZN(n622) );
  NAND2_X1 U684 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U685 ( .A1(G107), .A2(n888), .ZN(n625) );
  NAND2_X1 U686 ( .A1(G95), .A2(n892), .ZN(n624) );
  NAND2_X1 U687 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U688 ( .A1(n627), .A2(n626), .ZN(n898) );
  NAND2_X1 U689 ( .A1(G1991), .A2(n898), .ZN(n628) );
  XNOR2_X1 U690 ( .A(n628), .B(KEYINPUT97), .ZN(n630) );
  AND2_X1 U691 ( .A1(G1996), .A2(n883), .ZN(n629) );
  NOR2_X1 U692 ( .A1(n630), .A2(n629), .ZN(n982) );
  INV_X1 U693 ( .A(n982), .ZN(n633) );
  NOR2_X1 U694 ( .A1(G1986), .A2(G290), .ZN(n631) );
  NOR2_X1 U695 ( .A1(G1991), .A2(n898), .ZN(n973) );
  NOR2_X1 U696 ( .A1(n631), .A2(n973), .ZN(n632) );
  NOR2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U698 ( .A1(n977), .A2(n634), .ZN(n635) );
  XOR2_X1 U699 ( .A(KEYINPUT39), .B(n635), .Z(n636) );
  NOR2_X1 U700 ( .A1(n986), .A2(n636), .ZN(n637) );
  NOR2_X1 U701 ( .A1(n985), .A2(n637), .ZN(n638) );
  NOR2_X1 U702 ( .A1(n749), .A2(n638), .ZN(n639) );
  XNOR2_X1 U703 ( .A(n639), .B(KEYINPUT106), .ZN(n756) );
  NAND2_X2 U704 ( .A1(n641), .A2(n640), .ZN(n684) );
  NAND2_X1 U705 ( .A1(G8), .A2(n684), .ZN(n741) );
  NOR2_X1 U706 ( .A1(G1966), .A2(n741), .ZN(n712) );
  NOR2_X1 U707 ( .A1(G2084), .A2(n684), .ZN(n711) );
  NOR2_X1 U708 ( .A1(n712), .A2(n711), .ZN(n643) );
  INV_X1 U709 ( .A(KEYINPUT103), .ZN(n642) );
  XNOR2_X1 U710 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U711 ( .A1(G8), .A2(n644), .ZN(n645) );
  XNOR2_X1 U712 ( .A(n645), .B(KEYINPUT30), .ZN(n646) );
  NOR2_X1 U713 ( .A1(G168), .A2(n646), .ZN(n650) );
  XNOR2_X1 U714 ( .A(G1961), .B(KEYINPUT101), .ZN(n916) );
  NAND2_X1 U715 ( .A1(n684), .A2(n916), .ZN(n648) );
  INV_X1 U716 ( .A(n684), .ZN(n668) );
  XNOR2_X1 U717 ( .A(KEYINPUT25), .B(G2078), .ZN(n949) );
  NAND2_X1 U718 ( .A1(n668), .A2(n949), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n700) );
  NOR2_X1 U720 ( .A1(n700), .A2(G171), .ZN(n649) );
  NOR2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U722 ( .A(n651), .B(KEYINPUT31), .Z(n709) );
  INV_X1 U723 ( .A(G8), .ZN(n656) );
  NOR2_X1 U724 ( .A1(G1971), .A2(n741), .ZN(n653) );
  NOR2_X1 U725 ( .A1(G2090), .A2(n684), .ZN(n652) );
  NOR2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n654), .A2(G303), .ZN(n655) );
  OR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n704) );
  AND2_X1 U729 ( .A1(n709), .A2(n704), .ZN(n703) );
  NAND2_X1 U730 ( .A1(n668), .A2(G2072), .ZN(n657) );
  XOR2_X1 U731 ( .A(KEYINPUT27), .B(n657), .Z(n659) );
  NAND2_X1 U732 ( .A1(G1956), .A2(n684), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n693) );
  NAND2_X1 U734 ( .A1(G299), .A2(n693), .ZN(n660) );
  XOR2_X1 U735 ( .A(KEYINPUT28), .B(n660), .Z(n698) );
  NAND2_X1 U736 ( .A1(G66), .A2(n797), .ZN(n662) );
  NAND2_X1 U737 ( .A1(G54), .A2(n798), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U739 ( .A1(G79), .A2(n801), .ZN(n664) );
  NAND2_X1 U740 ( .A1(G92), .A2(n802), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n667), .B(KEYINPUT15), .ZN(n779) );
  NAND2_X1 U744 ( .A1(G1348), .A2(n684), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n668), .A2(G2067), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n670), .A2(n669), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n779), .A2(n690), .ZN(n689) );
  NAND2_X1 U748 ( .A1(n802), .A2(G81), .ZN(n671) );
  XNOR2_X1 U749 ( .A(n671), .B(KEYINPUT12), .ZN(n673) );
  NAND2_X1 U750 ( .A1(G68), .A2(n801), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U752 ( .A(n674), .B(KEYINPUT13), .ZN(n676) );
  NAND2_X1 U753 ( .A1(G43), .A2(n798), .ZN(n675) );
  NAND2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n680) );
  NAND2_X1 U755 ( .A1(G56), .A2(n797), .ZN(n677) );
  XNOR2_X1 U756 ( .A(n677), .B(KEYINPUT14), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n678), .B(KEYINPUT77), .ZN(n679) );
  NOR2_X1 U758 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U759 ( .A(KEYINPUT78), .B(n681), .Z(n1010) );
  INV_X1 U760 ( .A(G1996), .ZN(n682) );
  NOR2_X1 U761 ( .A1(n684), .A2(n682), .ZN(n683) );
  XOR2_X1 U762 ( .A(n683), .B(KEYINPUT26), .Z(n686) );
  NAND2_X1 U763 ( .A1(n684), .A2(G1341), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U765 ( .A1(n1010), .A2(n687), .ZN(n688) );
  NOR2_X1 U766 ( .A1(n689), .A2(n688), .ZN(n692) );
  AND2_X1 U767 ( .A1(n779), .A2(n690), .ZN(n691) );
  NOR2_X1 U768 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U769 ( .A1(G299), .A2(n693), .ZN(n694) );
  NOR2_X1 U770 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U771 ( .A(n696), .B(KEYINPUT102), .ZN(n697) );
  NOR2_X1 U772 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n699), .B(KEYINPUT29), .ZN(n702) );
  NAND2_X1 U774 ( .A1(n700), .A2(G171), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n710) );
  NAND2_X1 U776 ( .A1(n703), .A2(n710), .ZN(n707) );
  INV_X1 U777 ( .A(n704), .ZN(n705) );
  OR2_X1 U778 ( .A1(n705), .A2(G286), .ZN(n706) );
  NAND2_X1 U779 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U780 ( .A(n708), .B(KEYINPUT32), .ZN(n717) );
  AND2_X1 U781 ( .A1(n710), .A2(n709), .ZN(n715) );
  AND2_X1 U782 ( .A1(G8), .A2(n711), .ZN(n713) );
  OR2_X1 U783 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U784 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n737) );
  NOR2_X1 U786 ( .A1(G1976), .A2(G288), .ZN(n997) );
  INV_X1 U787 ( .A(n997), .ZN(n720) );
  NOR2_X1 U788 ( .A1(G1971), .A2(G303), .ZN(n718) );
  XOR2_X1 U789 ( .A(n718), .B(KEYINPUT104), .Z(n719) );
  AND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n721) );
  AND2_X1 U791 ( .A1(n737), .A2(n721), .ZN(n722) );
  XNOR2_X1 U792 ( .A(n722), .B(KEYINPUT105), .ZN(n728) );
  NAND2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n1006) );
  INV_X1 U794 ( .A(n1006), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n997), .A2(KEYINPUT33), .ZN(n724) );
  NOR2_X1 U796 ( .A1(n724), .A2(n741), .ZN(n730) );
  INV_X1 U797 ( .A(n730), .ZN(n725) );
  AND2_X1 U798 ( .A1(n515), .A2(n725), .ZN(n726) );
  XOR2_X1 U799 ( .A(G1981), .B(G305), .Z(n993) );
  AND2_X1 U800 ( .A1(n726), .A2(n993), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n734) );
  INV_X1 U802 ( .A(n993), .ZN(n732) );
  INV_X1 U803 ( .A(KEYINPUT33), .ZN(n729) );
  OR2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n731) );
  OR2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n734), .A2(n733), .ZN(n746) );
  NOR2_X1 U807 ( .A1(G2090), .A2(G303), .ZN(n735) );
  NAND2_X1 U808 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  AND2_X1 U810 ( .A1(n738), .A2(n741), .ZN(n744) );
  NOR2_X1 U811 ( .A1(G1981), .A2(G305), .ZN(n739) );
  XOR2_X1 U812 ( .A(n739), .B(KEYINPUT24), .Z(n740) );
  NOR2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U814 ( .A(n742), .B(KEYINPUT100), .ZN(n743) );
  OR2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U816 ( .A1(n746), .A2(n745), .ZN(n754) );
  NOR2_X1 U817 ( .A1(n986), .A2(n633), .ZN(n747) );
  NOR2_X1 U818 ( .A1(n749), .A2(n747), .ZN(n748) );
  XNOR2_X1 U819 ( .A(n748), .B(KEYINPUT99), .ZN(n752) );
  INV_X1 U820 ( .A(n749), .ZN(n750) );
  XNOR2_X1 U821 ( .A(G1986), .B(G290), .ZN(n999) );
  NAND2_X1 U822 ( .A1(n750), .A2(n999), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U824 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U825 ( .A1(n756), .A2(n755), .ZN(n758) );
  INV_X1 U826 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U827 ( .A(G2451), .B(G2446), .ZN(n768) );
  XOR2_X1 U828 ( .A(G2430), .B(KEYINPUT109), .Z(n760) );
  XNOR2_X1 U829 ( .A(G2454), .B(G2435), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n760), .B(n759), .ZN(n764) );
  XOR2_X1 U831 ( .A(G2438), .B(KEYINPUT108), .Z(n762) );
  XNOR2_X1 U832 ( .A(G1341), .B(G1348), .ZN(n761) );
  XNOR2_X1 U833 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U834 ( .A(n764), .B(n763), .Z(n766) );
  XNOR2_X1 U835 ( .A(G2443), .B(G2427), .ZN(n765) );
  XNOR2_X1 U836 ( .A(n766), .B(n765), .ZN(n767) );
  XNOR2_X1 U837 ( .A(n768), .B(n767), .ZN(n769) );
  AND2_X1 U838 ( .A1(n769), .A2(G14), .ZN(G401) );
  INV_X1 U839 ( .A(G860), .ZN(n778) );
  OR2_X1 U840 ( .A1(n778), .A2(n1010), .ZN(G153) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  INV_X1 U843 ( .A(G120), .ZN(G236) );
  INV_X1 U844 ( .A(G69), .ZN(G235) );
  INV_X1 U845 ( .A(G108), .ZN(G238) );
  NAND2_X1 U846 ( .A1(G94), .A2(G452), .ZN(n770) );
  XNOR2_X1 U847 ( .A(n770), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U849 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U850 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n773) );
  INV_X1 U851 ( .A(G223), .ZN(n837) );
  NAND2_X1 U852 ( .A1(G567), .A2(n837), .ZN(n772) );
  XNOR2_X1 U853 ( .A(n773), .B(n772), .ZN(G234) );
  NAND2_X1 U854 ( .A1(G301), .A2(G868), .ZN(n775) );
  INV_X1 U855 ( .A(G868), .ZN(n818) );
  NAND2_X1 U856 ( .A1(n779), .A2(n818), .ZN(n774) );
  NAND2_X1 U857 ( .A1(n775), .A2(n774), .ZN(G284) );
  NOR2_X1 U858 ( .A1(G286), .A2(n818), .ZN(n777) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n776) );
  NOR2_X1 U860 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U861 ( .A1(n778), .A2(G559), .ZN(n780) );
  INV_X1 U862 ( .A(n779), .ZN(n996) );
  NAND2_X1 U863 ( .A1(n780), .A2(n996), .ZN(n781) );
  XNOR2_X1 U864 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U865 ( .A1(n996), .A2(G868), .ZN(n782) );
  NOR2_X1 U866 ( .A1(G559), .A2(n782), .ZN(n783) );
  XNOR2_X1 U867 ( .A(n783), .B(KEYINPUT82), .ZN(n785) );
  NOR2_X1 U868 ( .A1(n1010), .A2(G868), .ZN(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(G282) );
  XNOR2_X1 U870 ( .A(G2100), .B(KEYINPUT85), .ZN(n796) );
  XOR2_X1 U871 ( .A(KEYINPUT18), .B(KEYINPUT84), .Z(n787) );
  NAND2_X1 U872 ( .A1(G123), .A2(n889), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U874 ( .A(n788), .B(KEYINPUT83), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n888), .A2(G111), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U877 ( .A1(G135), .A2(n529), .ZN(n792) );
  NAND2_X1 U878 ( .A1(G99), .A2(n892), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n972) );
  XNOR2_X1 U881 ( .A(n972), .B(G2096), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(G156) );
  NAND2_X1 U883 ( .A1(G67), .A2(n797), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n806) );
  NAND2_X1 U886 ( .A1(G80), .A2(n801), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U889 ( .A1(n806), .A2(n805), .ZN(n817) );
  NAND2_X1 U890 ( .A1(G559), .A2(n996), .ZN(n807) );
  XNOR2_X1 U891 ( .A(n807), .B(n1010), .ZN(n815) );
  XNOR2_X1 U892 ( .A(KEYINPUT86), .B(n815), .ZN(n808) );
  NOR2_X1 U893 ( .A1(G860), .A2(n808), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n817), .B(n809), .ZN(G145) );
  XNOR2_X1 U895 ( .A(KEYINPUT19), .B(G288), .ZN(n814) );
  XNOR2_X1 U896 ( .A(G166), .B(n817), .ZN(n812) );
  XNOR2_X1 U897 ( .A(G305), .B(G299), .ZN(n810) );
  XNOR2_X1 U898 ( .A(n810), .B(G290), .ZN(n811) );
  XNOR2_X1 U899 ( .A(n812), .B(n811), .ZN(n813) );
  XNOR2_X1 U900 ( .A(n814), .B(n813), .ZN(n844) );
  XNOR2_X1 U901 ( .A(n815), .B(n844), .ZN(n816) );
  NAND2_X1 U902 ( .A1(n816), .A2(G868), .ZN(n820) );
  NAND2_X1 U903 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U904 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U905 ( .A(KEYINPUT89), .B(n821), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U910 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G235), .A2(G236), .ZN(n826) );
  XOR2_X1 U913 ( .A(KEYINPUT90), .B(n826), .Z(n827) );
  NOR2_X1 U914 ( .A1(G238), .A2(n827), .ZN(n828) );
  NAND2_X1 U915 ( .A1(G57), .A2(n828), .ZN(n913) );
  NAND2_X1 U916 ( .A1(n913), .A2(G567), .ZN(n833) );
  NOR2_X1 U917 ( .A1(G220), .A2(G219), .ZN(n829) );
  XOR2_X1 U918 ( .A(KEYINPUT22), .B(n829), .Z(n830) );
  NOR2_X1 U919 ( .A1(G218), .A2(n830), .ZN(n831) );
  NAND2_X1 U920 ( .A1(G96), .A2(n831), .ZN(n914) );
  NAND2_X1 U921 ( .A1(n914), .A2(G2106), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n833), .A2(n832), .ZN(n915) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n834) );
  XOR2_X1 U924 ( .A(KEYINPUT91), .B(n834), .Z(n835) );
  NOR2_X1 U925 ( .A1(n915), .A2(n835), .ZN(n836) );
  XNOR2_X1 U926 ( .A(KEYINPUT92), .B(n836), .ZN(n840) );
  NAND2_X1 U927 ( .A1(G36), .A2(n840), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U930 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U933 ( .A(KEYINPUT110), .B(n841), .ZN(G188) );
  XOR2_X1 U934 ( .A(KEYINPUT114), .B(n996), .Z(n843) );
  XNOR2_X1 U935 ( .A(G301), .B(n1010), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(n846) );
  XNOR2_X1 U937 ( .A(G286), .B(n844), .ZN(n845) );
  XNOR2_X1 U938 ( .A(n846), .B(n845), .ZN(n847) );
  NOR2_X1 U939 ( .A1(G37), .A2(n847), .ZN(n848) );
  XOR2_X1 U940 ( .A(KEYINPUT115), .B(n848), .Z(G397) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2084), .Z(n850) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2072), .ZN(n849) );
  XNOR2_X1 U943 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U944 ( .A(n851), .B(G2096), .Z(n853) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2090), .ZN(n852) );
  XNOR2_X1 U946 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U947 ( .A(G2100), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U948 ( .A(KEYINPUT111), .B(G2678), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U950 ( .A(n857), .B(n856), .Z(G227) );
  XNOR2_X1 U951 ( .A(G1991), .B(KEYINPUT41), .ZN(n867) );
  XOR2_X1 U952 ( .A(G1986), .B(G1971), .Z(n859) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1956), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U955 ( .A(G1961), .B(G1966), .Z(n861) );
  XNOR2_X1 U956 ( .A(G1981), .B(G1976), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U958 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U959 ( .A(KEYINPUT112), .B(G2474), .ZN(n864) );
  XNOR2_X1 U960 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U961 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G124), .A2(n889), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n888), .A2(G112), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U966 ( .A1(G136), .A2(n529), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G100), .A2(n892), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U969 ( .A1(n874), .A2(n873), .ZN(G162) );
  XNOR2_X1 U970 ( .A(n972), .B(G162), .ZN(n882) );
  NAND2_X1 U971 ( .A1(G139), .A2(n529), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G103), .A2(n892), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U974 ( .A1(G115), .A2(n888), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G127), .A2(n889), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n968) );
  XNOR2_X1 U979 ( .A(n882), .B(n968), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n884), .B(n883), .ZN(n887) );
  XOR2_X1 U981 ( .A(G160), .B(n885), .Z(n886) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n904) );
  NAND2_X1 U983 ( .A1(G118), .A2(n888), .ZN(n891) );
  NAND2_X1 U984 ( .A1(G130), .A2(n889), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n897) );
  NAND2_X1 U986 ( .A1(G142), .A2(n529), .ZN(n894) );
  NAND2_X1 U987 ( .A1(G106), .A2(n892), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U989 ( .A(n895), .B(KEYINPUT45), .Z(n896) );
  NOR2_X1 U990 ( .A1(n897), .A2(n896), .ZN(n899) );
  XNOR2_X1 U991 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U992 ( .A(n900), .B(KEYINPUT48), .Z(n902) );
  XNOR2_X1 U993 ( .A(G164), .B(KEYINPUT46), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U995 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U996 ( .A1(G37), .A2(n905), .ZN(n906) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(n906), .Z(G395) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U999 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1000 ( .A1(G397), .A2(n908), .ZN(n912) );
  NOR2_X1 U1001 ( .A1(n915), .A2(G401), .ZN(n909) );
  XOR2_X1 U1002 ( .A(KEYINPUT116), .B(n909), .Z(n910) );
  NOR2_X1 U1003 ( .A1(G395), .A2(n910), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(n912), .A2(n911), .ZN(G225) );
  XNOR2_X1 U1005 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(G325) );
  INV_X1 U1009 ( .A(G325), .ZN(G261) );
  INV_X1 U1010 ( .A(n915), .ZN(G319) );
  INV_X1 U1011 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1012 ( .A(G5), .B(n916), .ZN(n937) );
  XOR2_X1 U1013 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n923) );
  XNOR2_X1 U1014 ( .A(G1971), .B(G22), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(G24), .B(G1986), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1017 ( .A(G1976), .B(KEYINPUT126), .Z(n919) );
  XNOR2_X1 U1018 ( .A(G23), .B(n919), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n935) );
  XNOR2_X1 U1021 ( .A(G1348), .B(KEYINPUT59), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(G4), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(G1981), .B(G6), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G1341), .B(G19), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(KEYINPUT124), .B(G1956), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(G20), .B(n929), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT125), .B(n932), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT60), .B(n933), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(G21), .B(G1966), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n940), .B(KEYINPUT61), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(G16), .B(KEYINPUT123), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(G11), .A2(n943), .ZN(n967) );
  XOR2_X1 U1040 ( .A(G34), .B(KEYINPUT121), .Z(n945) );
  XNOR2_X1 U1041 ( .A(G2084), .B(KEYINPUT54), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n945), .B(n944), .ZN(n963) );
  XNOR2_X1 U1043 ( .A(G1996), .B(G32), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n954) );
  XOR2_X1 U1046 ( .A(G2067), .B(G26), .Z(n948) );
  NAND2_X1 U1047 ( .A1(n948), .A2(G28), .ZN(n952) );
  XOR2_X1 U1048 ( .A(G27), .B(n949), .Z(n950) );
  XNOR2_X1 U1049 ( .A(KEYINPUT118), .B(n950), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G25), .B(G1991), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1054 ( .A(n957), .B(KEYINPUT119), .Z(n958) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G35), .B(G2090), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1058 ( .A(KEYINPUT120), .B(n961), .Z(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n964), .ZN(n965) );
  XOR2_X1 U1061 ( .A(KEYINPUT55), .B(n965), .Z(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n992) );
  XOR2_X1 U1063 ( .A(G2072), .B(n968), .Z(n970) );
  XOR2_X1 U1064 ( .A(G164), .B(G2078), .Z(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(KEYINPUT50), .B(n971), .ZN(n975) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n980) );
  XOR2_X1 U1069 ( .A(G2090), .B(G162), .Z(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n978), .B(KEYINPUT51), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G160), .B(G2084), .Z(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n988) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(KEYINPUT52), .B(n989), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n990), .A2(G29), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n1018) );
  XOR2_X1 U1081 ( .A(KEYINPUT56), .B(G16), .Z(n1016) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G168), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(KEYINPUT57), .ZN(n1005) );
  XNOR2_X1 U1085 ( .A(n996), .B(G1348), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(KEYINPUT122), .B(n997), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G301), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1014) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G166), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G299), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1096 ( .A(n1010), .B(G1341), .Z(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1099 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1100 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(n1019), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1102 ( .A(G311), .ZN(G150) );
endmodule

