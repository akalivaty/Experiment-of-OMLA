//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n474), .A2(G137), .A3(new_n475), .A4(new_n464), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND3_X1   g055(.A1(new_n474), .A2(G2105), .A3(new_n464), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n475), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n474), .A2(new_n475), .A3(new_n464), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n486), .A2(KEYINPUT69), .A3(G136), .ZN(new_n487));
  AOI21_X1  g062(.A(KEYINPUT69), .B1(new_n486), .B2(G136), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n482), .B1(new_n483), .B2(new_n484), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  AND2_X1   g067(.A1(new_n475), .A2(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n474), .A2(new_n464), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n467), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n475), .C1(new_n496), .C2(KEYINPUT73), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n496), .A2(KEYINPUT73), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n474), .A2(new_n464), .A3(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(KEYINPUT72), .A3(new_n504), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n500), .B1(new_n507), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT74), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT74), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n516), .A2(G50), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n513), .A2(new_n514), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n521), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT75), .B(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n516), .A2(G51), .ZN(new_n531));
  INV_X1    g106(.A(new_n521), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n532), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n526), .A2(G89), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND2_X1  g116(.A1(new_n526), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n516), .A2(G52), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n521), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(new_n517), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n521), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n516), .A2(G43), .B1(new_n517), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n526), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n521), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n526), .A2(G91), .B1(G651), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(G53), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n566));
  XOR2_X1   g141(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n567));
  OR2_X1    g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n566), .B1(KEYINPUT76), .B2(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(KEYINPUT77), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT77), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n526), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n516), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n521), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n526), .A2(G86), .B1(new_n517), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n516), .A2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(G85), .A2(new_n526), .B1(new_n516), .B2(G47), .ZN(new_n584));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n521), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n587), .A2(KEYINPUT78), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n517), .B1(new_n587), .B2(KEYINPUT78), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G171), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n526), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n515), .A2(KEYINPUT79), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n515), .B2(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT80), .Z(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n521), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n595), .A2(new_n597), .B1(G651), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n594), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n591), .B1(new_n608), .B2(G868), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT82), .ZN(G284));
  XOR2_X1   g185(.A(new_n609), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(new_n565), .ZN(new_n613));
  INV_X1    g188(.A(new_n572), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n570), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n612), .B1(new_n615), .B2(G868), .ZN(G280));
  XOR2_X1   g191(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n607), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND3_X1  g194(.A1(new_n607), .A2(KEYINPUT85), .A3(new_n618), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(KEYINPUT85), .B1(new_n607), .B2(new_n618), .ZN(new_n622));
  OAI21_X1  g197(.A(G868), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n556), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT86), .Z(G323));
  XNOR2_X1  g200(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n626));
  XNOR2_X1  g201(.A(G323), .B(new_n626), .ZN(G282));
  NAND2_X1  g202(.A1(new_n495), .A2(new_n477), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n486), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n475), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT88), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(G14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT89), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n669), .A2(new_n671), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n674), .A3(new_n672), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n676), .B(new_n679), .C1(new_n674), .C2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(G229));
  NAND2_X1  g263(.A1(G115), .A2(G2104), .ZN(new_n689));
  INV_X1    g264(.A(G127), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n467), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G2105), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT25), .Z(new_n694));
  INV_X1    g269(.A(G139), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n692), .B(new_n694), .C1(new_n485), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT99), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n698), .B2(G33), .ZN(new_n700));
  INV_X1    g275(.A(G2072), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT100), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n698), .A2(G27), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G164), .B2(new_n698), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G2078), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(G2078), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT30), .B(G28), .ZN(new_n710));
  OR2_X1    g285(.A1(KEYINPUT31), .A2(G11), .ZN(new_n711));
  NAND2_X1  g286(.A1(KEYINPUT31), .A2(G11), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n710), .A2(new_n698), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n714), .A2(G34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(G34), .ZN(new_n716));
  AOI21_X1  g291(.A(G29), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n479), .B2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G2084), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n713), .B1(new_n636), .B2(new_n698), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(new_n718), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G5), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G171), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1966), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n722), .A2(G21), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G286), .B2(G16), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n721), .B1(G1961), .B2(new_n724), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n727), .A2(new_n725), .B1(new_n724), .B2(G1961), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n698), .A2(G32), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n486), .A2(G141), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n481), .A2(G129), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AOI22_X1  g311(.A1(G105), .A2(new_n477), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n731), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n730), .B1(new_n739), .B2(new_n698), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n729), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n728), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n703), .A2(new_n709), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n698), .A2(G35), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT101), .Z(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n698), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT29), .B(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n722), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n615), .B2(new_n722), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n722), .A2(G4), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n607), .B2(new_n722), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT96), .B(G1348), .Z(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n722), .A2(G19), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n556), .B2(new_n722), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1341), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n486), .A2(G140), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n481), .A2(G128), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n475), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G29), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n698), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT97), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n761), .A2(new_n762), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n761), .A2(new_n780), .A3(new_n762), .A4(new_n777), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n746), .A2(new_n757), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(KEYINPUT103), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n745), .A2(new_n751), .A3(new_n756), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT103), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n784), .A2(new_n785), .A3(new_n779), .A4(new_n781), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT104), .ZN(new_n788));
  NOR2_X1   g363(.A1(G16), .A2(G23), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G288), .B2(new_n722), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT95), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT33), .B(G1976), .Z(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n722), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n722), .ZN(new_n798));
  INV_X1    g373(.A(G1971), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n795), .A2(new_n796), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n698), .A2(G25), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n486), .A2(G131), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT92), .Z(new_n808));
  OR2_X1    g383(.A1(new_n475), .A2(G107), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n481), .A2(G119), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n806), .B1(new_n814), .B2(new_n698), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT93), .Z(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  OR2_X1    g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n819));
  MUX2_X1   g394(.A(G24), .B(G290), .S(G16), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1986), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n816), .B2(new_n817), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n805), .A2(new_n818), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT36), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n787), .A2(new_n788), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n788), .B1(new_n787), .B2(new_n824), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n787), .A2(new_n824), .ZN(G150));
  NAND2_X1  g403(.A1(new_n607), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n521), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n516), .A2(G55), .B1(new_n517), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n526), .A2(G93), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(new_n555), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n555), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n830), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n836), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(new_n813), .B(new_n629), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n486), .A2(G142), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n481), .A2(G130), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n851));
  INV_X1    g426(.A(G118), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n850), .A2(new_n851), .B1(new_n852), .B2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n851), .B2(new_n850), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n847), .B(new_n855), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n499), .A2(new_n495), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n502), .A3(new_n504), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n770), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n738), .ZN(new_n862));
  INV_X1    g437(.A(new_n697), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n696), .B2(new_n862), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n856), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n856), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n636), .B(new_n479), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n491), .B(new_n869), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT106), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n866), .A2(new_n867), .A3(new_n873), .A4(new_n870), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n868), .B2(new_n871), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g453(.A1(new_n615), .A2(new_n594), .A3(new_n602), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n603), .A2(G299), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT107), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n839), .ZN(new_n884));
  INV_X1    g459(.A(new_n622), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n620), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n621), .A2(new_n622), .A3(new_n839), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n839), .B1(new_n621), .B2(new_n622), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n620), .A3(new_n884), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n879), .A2(new_n880), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n881), .A2(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n888), .A2(KEYINPUT108), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n898), .B(new_n883), .C1(new_n886), .C2(new_n887), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n901));
  INV_X1    g476(.A(G288), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G166), .B(G305), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n903), .B(new_n904), .Z(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n906), .A3(new_n899), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n901), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n905), .B1(new_n901), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g484(.A(G868), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G868), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n836), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(G295));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n912), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n837), .A2(G301), .A3(new_n838), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G301), .B1(new_n837), .B2(new_n838), .ZN(new_n920));
  OAI21_X1  g495(.A(G286), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n920), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(G168), .A3(new_n918), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n881), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n893), .A2(new_n894), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n923), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n917), .B1(new_n928), .B2(new_n905), .ZN(new_n929));
  INV_X1    g504(.A(new_n927), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n924), .B1(new_n930), .B2(new_n895), .ZN(new_n931));
  INV_X1    g506(.A(new_n905), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n916), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n882), .B2(new_n927), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n926), .A2(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n894), .A2(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n931), .B2(new_n932), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT43), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n915), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n929), .B2(new_n933), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n940), .A3(new_n916), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n942), .A2(new_n945), .A3(KEYINPUT110), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n934), .A2(new_n941), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT44), .ZN(new_n949));
  INV_X1    g524(.A(new_n944), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n928), .A2(new_n905), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n916), .B1(new_n940), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n915), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n947), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n946), .A2(new_n954), .ZN(G397));
  XNOR2_X1  g530(.A(new_n770), .B(G2067), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT111), .ZN(new_n957));
  INV_X1    g532(.A(G1996), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n738), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n813), .B(new_n817), .Z(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n500), .B2(new_n505), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n470), .A2(G40), .A3(new_n476), .A4(new_n478), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n962), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT48), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n958), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT46), .Z(new_n975));
  NAND2_X1  g550(.A1(new_n957), .A2(new_n739), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(new_n968), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n814), .A2(new_n817), .ZN(new_n979));
  OAI22_X1  g554(.A1(new_n960), .A2(new_n979), .B1(G2067), .B2(new_n770), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n973), .B(new_n978), .C1(new_n968), .C2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT126), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n967), .B1(new_n964), .B2(KEYINPUT50), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n502), .A2(KEYINPUT72), .A3(new_n504), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT72), .B1(new_n502), .B2(new_n504), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n859), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n963), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1956), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n965), .C1(G164), .C2(G1384), .ZN(new_n993));
  INV_X1    g568(.A(new_n967), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT45), .B(new_n963), .C1(new_n500), .C2(new_n505), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n992), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT45), .B1(new_n986), .B2(new_n963), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n993), .B(new_n994), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT56), .B(G2072), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n991), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n613), .A2(KEYINPUT57), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n568), .A2(new_n569), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1005), .B1(new_n615), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1348), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n987), .B1(new_n986), .B2(new_n963), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n994), .B1(new_n964), .B2(KEYINPUT50), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OR3_X1    g587(.A1(new_n964), .A2(G2067), .A3(new_n967), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1008), .B1(new_n1015), .B2(new_n608), .ZN(new_n1016));
  AOI22_X1  g591(.A1(G299), .A2(KEYINPUT57), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n965), .B1(G164), .B2(G1384), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n996), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(new_n994), .A3(new_n993), .A4(new_n1000), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1020), .A3(new_n991), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n1021), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1008), .A2(KEYINPUT117), .A3(new_n1021), .A4(KEYINPUT61), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1012), .A2(KEYINPUT60), .A3(new_n1013), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1012), .A2(KEYINPUT118), .A3(KEYINPUT60), .A4(new_n1013), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n607), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT60), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1014), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1032), .B(new_n1034), .C1(new_n607), .C2(new_n1030), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT116), .B(G1996), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n964), .A2(new_n967), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT58), .B(G1341), .ZN(new_n1038));
  OAI22_X1  g613(.A1(new_n999), .A2(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n556), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT59), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1042), .A3(new_n556), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1008), .A2(new_n1021), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT61), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1035), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1022), .B1(new_n1027), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT119), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(new_n1022), .C1(new_n1027), .C2(new_n1048), .ZN(new_n1052));
  INV_X1    g627(.A(G2078), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1019), .A2(new_n1053), .A3(new_n994), .A4(new_n993), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n967), .B1(new_n964), .B2(new_n965), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n986), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1053), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT122), .A4(new_n1053), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT53), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1961), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1056), .A2(new_n1063), .A3(G301), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1055), .B(G2078), .C1(new_n967), .C2(KEYINPUT123), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(new_n995), .A3(new_n966), .A4(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1065), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT54), .B1(new_n1072), .B2(G301), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT125), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1056), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G171), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(KEYINPUT54), .A4(new_n1066), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1072), .A2(new_n1081), .A3(G301), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1056), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(G171), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT124), .B1(new_n1076), .B2(G171), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1082), .B(new_n1083), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G303), .A2(G8), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT55), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n989), .A2(G2090), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n799), .B2(new_n999), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT113), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1037), .A2(new_n1092), .ZN(new_n1095));
  INV_X1    g670(.A(G1976), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(G288), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT52), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  INV_X1    g674(.A(G1981), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n581), .A2(new_n1100), .A3(new_n582), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n581), .B2(new_n582), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(G305), .A2(G1981), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n581), .A2(new_n1100), .A3(new_n582), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(KEYINPUT49), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1106), .A3(new_n1095), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(G288), .B2(new_n1096), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1095), .B(new_n1108), .C1(new_n1096), .C2(G288), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1098), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n999), .A2(new_n799), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1112));
  INV_X1    g687(.A(G2090), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1092), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1089), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1110), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT113), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1118), .B(new_n1089), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1094), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1121), .A2(KEYINPUT51), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(KEYINPUT51), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n725), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1112), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(G2084), .ZN(new_n1128));
  OAI211_X1 g703(.A(G8), .B(new_n1124), .C1(new_n1128), .C2(G286), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(G8), .A3(G286), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1112), .A2(new_n719), .B1(new_n1125), .B2(new_n725), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1092), .B1(new_n1131), .B2(G168), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1129), .B(new_n1130), .C1(new_n1132), .C2(new_n1123), .ZN(new_n1133));
  AND4_X1   g708(.A1(new_n1080), .A2(new_n1087), .A3(new_n1120), .A4(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1050), .A2(new_n1052), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n1110), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1107), .A2(new_n1096), .A3(new_n902), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1105), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1095), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1133), .A2(KEYINPUT62), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1132), .A2(new_n1123), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1144), .A3(new_n1085), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1120), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1140), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1098), .A2(new_n1109), .A3(new_n1107), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT115), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1128), .A2(G8), .A3(G168), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT114), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT114), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1128), .A2(new_n1153), .A3(G8), .A4(G168), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1155), .A2(KEYINPUT63), .A3(new_n1136), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1155), .A2(new_n1094), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1150), .A2(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1147), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1135), .A2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(G290), .B(G1986), .Z(new_n1162));
  AOI21_X1  g737(.A(new_n969), .B1(new_n962), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n982), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  AOI211_X1 g740(.A(KEYINPUT126), .B(new_n1163), .C1(new_n1135), .C2(new_n1160), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n981), .B1(new_n1165), .B2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g742(.A1(new_n460), .A2(G227), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n654), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g744(.A(new_n1170), .B(KEYINPUT127), .Z(new_n1171));
  NOR2_X1   g745(.A1(new_n1171), .A2(G229), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n877), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n950), .A2(new_n952), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1173), .A2(new_n1174), .ZN(G308));
  INV_X1    g749(.A(G308), .ZN(G225));
endmodule


