//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT90), .B1(new_n208), .B2(G43gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n207), .A2(new_n213), .A3(new_n211), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT17), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT17), .A4(new_n216), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT91), .A2(G1gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT16), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(G1gat), .B1(new_n223), .B2(KEYINPUT91), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT92), .ZN(new_n228));
  OAI22_X1  g027(.A1(new_n226), .A2(new_n227), .B1(new_n228), .B2(G8gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(G8gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n229), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n222), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n229), .B(new_n230), .ZN(new_n235));
  INV_X1    g034(.A(new_n218), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n233), .A2(new_n234), .A3(new_n237), .A4(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n234), .B(KEYINPUT13), .Z(new_n243));
  INV_X1    g042(.A(new_n237), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n235), .A2(new_n236), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(G169gat), .B(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT12), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n240), .A2(new_n242), .A3(new_n246), .A4(new_n253), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT31), .B(G50gat), .Z(new_n259));
  NAND2_X1  g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT2), .ZN(new_n261));
  INV_X1    g060(.A(G141gat), .ZN(new_n262));
  INV_X1    g061(.A(G148gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT77), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G162gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n260), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n266), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT78), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(KEYINPUT78), .A3(new_n266), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n270), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  INV_X1    g083(.A(G218gat), .ZN(new_n285));
  OR2_X1    g084(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n283), .B(new_n284), .C1(new_n288), .C2(KEYINPUT22), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n287), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT75), .A2(G211gat), .ZN(new_n293));
  OAI21_X1  g092(.A(G218gat), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT22), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n296), .A2(KEYINPUT84), .A3(new_n283), .A4(new_n284), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n283), .B1(new_n288), .B2(KEYINPUT22), .ZN(new_n298));
  INV_X1    g097(.A(new_n284), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n291), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n282), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n289), .ZN(new_n306));
  INV_X1    g105(.A(new_n270), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n277), .A2(KEYINPUT78), .A3(new_n266), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT78), .B1(new_n277), .B2(new_n266), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n304), .B(new_n307), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n310), .B2(new_n302), .ZN(new_n311));
  INV_X1    g110(.A(G228gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  OAI22_X1  g112(.A1(new_n305), .A2(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n310), .A2(new_n302), .ZN(new_n315));
  INV_X1    g114(.A(new_n306), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n312), .A2(new_n313), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT3), .B1(new_n306), .B2(new_n302), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n317), .B(new_n318), .C1(new_n282), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G22gat), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n321), .B1(new_n314), .B2(new_n320), .ZN(new_n323));
  XNOR2_X1  g122(.A(G78gat), .B(G106gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n304), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n318), .B1(new_n329), .B2(new_n317), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n318), .B1(new_n319), .B2(new_n282), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(new_n311), .ZN(new_n332));
  OAI21_X1  g131(.A(G22gat), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n324), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n259), .B1(new_n326), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n325), .B1(new_n322), .B2(new_n323), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n334), .A3(new_n324), .ZN(new_n338));
  INV_X1    g137(.A(new_n259), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT39), .ZN(new_n342));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n282), .A2(new_n345), .A3(new_n304), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT79), .B1(new_n328), .B2(KEYINPUT3), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT69), .B(G127gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G134gat), .ZN(new_n349));
  INV_X1    g148(.A(G120gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G113gat), .ZN(new_n351));
  INV_X1    g150(.A(G113gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G120gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n355));
  INV_X1    g154(.A(G127gat), .ZN(new_n356));
  INV_X1    g155(.A(G134gat), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n354), .A2(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT70), .B(G113gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n351), .B1(new_n359), .B2(new_n350), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(G127gat), .A2(G134gat), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT1), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n349), .A2(new_n358), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n310), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n346), .A2(new_n347), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n282), .B2(new_n364), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n364), .B(new_n307), .C1(new_n308), .C2(new_n309), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(KEYINPUT4), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n282), .A2(KEYINPUT83), .A3(new_n368), .A4(new_n364), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n342), .B(new_n344), .C1(new_n367), .C2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT0), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT82), .ZN(new_n378));
  XOR2_X1   g177(.A(G57gat), .B(G85gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n374), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n347), .A2(new_n366), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n328), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n343), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n328), .A2(new_n365), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n371), .A3(new_n343), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT39), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(KEYINPUT85), .A3(KEYINPUT39), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n375), .B(new_n380), .C1(new_n385), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT40), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n386), .A2(new_n371), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n344), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT5), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n344), .B1(new_n382), .B2(new_n383), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n369), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT80), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT81), .B1(new_n371), .B2(KEYINPUT4), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n282), .A2(new_n406), .A3(new_n368), .A4(new_n364), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n402), .A2(new_n404), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n399), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n344), .A2(KEYINPUT5), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n367), .A2(new_n374), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n396), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n344), .B1(new_n367), .B2(new_n374), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n414), .A2(new_n390), .A3(new_n391), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n415), .A2(KEYINPUT40), .A3(new_n380), .A4(new_n375), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n395), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418));
  INV_X1    g217(.A(G169gat), .ZN(new_n419));
  INV_X1    g218(.A(G176gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT23), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT65), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT23), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(G169gat), .B2(G176gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT65), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n423), .B1(new_n421), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n428), .A2(KEYINPUT64), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(KEYINPUT64), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(G183gat), .A2(G190gat), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT25), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n428), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n421), .A2(new_n425), .A3(KEYINPUT25), .A4(new_n418), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT68), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n443), .A2(KEYINPUT26), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n418), .B1(new_n443), .B2(KEYINPUT26), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n433), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT27), .B(G183gat), .ZN(new_n447));
  INV_X1    g246(.A(G190gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n450));
  OR2_X1    g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n450), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G226gat), .A2(G233gat), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n442), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT66), .B1(new_n437), .B2(new_n441), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT25), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n426), .A2(new_n421), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n424), .A2(G169gat), .A3(G176gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n418), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n434), .B1(new_n430), .B2(new_n429), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464));
  INV_X1    g263(.A(new_n441), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n453), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n456), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n454), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(KEYINPUT29), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n455), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n316), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n456), .A2(new_n466), .A3(new_n467), .A4(new_n469), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n470), .B1(new_n442), .B2(new_n453), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n316), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n477), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT76), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n475), .B1(new_n471), .B2(new_n316), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT76), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n485), .A3(new_n480), .ZN(new_n486));
  AOI211_X1 g285(.A(new_n480), .B(new_n475), .C1(new_n316), .C2(new_n471), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n481), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n341), .B1(new_n417), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n381), .A2(new_n384), .A3(new_n410), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n400), .A2(new_n408), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n380), .B(new_n492), .C1(new_n493), .C2(new_n399), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n413), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n480), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n484), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n471), .B2(new_n306), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n473), .A2(new_n474), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n316), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT38), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n487), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(KEYINPUT6), .B(new_n396), .C1(new_n409), .C2(new_n412), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n496), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n506), .A2(KEYINPUT86), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n496), .A2(new_n504), .A3(new_n508), .A4(new_n505), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT37), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n499), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT38), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n491), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT87), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(KEYINPUT86), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n509), .A3(new_n512), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(KEYINPUT87), .A3(new_n491), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n505), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n490), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n516), .A2(new_n519), .B1(new_n523), .B2(new_n341), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n456), .A2(new_n364), .A3(new_n466), .A4(new_n467), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n468), .A2(new_n365), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n468), .A2(new_n526), .A3(new_n365), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(G227gat), .A3(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT32), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT33), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G15gat), .B(G43gat), .Z(new_n536));
  XNOR2_X1  g335(.A(G71gat), .B(G99gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n533), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n532), .B(KEYINPUT32), .C1(new_n534), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G227gat), .A2(G233gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n529), .A2(new_n543), .A3(new_n530), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT34), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT34), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n529), .A2(new_n549), .A3(new_n543), .A4(new_n530), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n550), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT72), .B1(new_n544), .B2(KEYINPUT34), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n547), .A2(KEYINPUT73), .A3(new_n548), .A4(new_n550), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n559), .A2(KEYINPUT74), .A3(new_n542), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT74), .B1(new_n559), .B2(new_n542), .ZN(new_n561));
  OAI211_X1 g360(.A(KEYINPUT36), .B(new_n553), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n542), .A2(new_n551), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n552), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n524), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n341), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n553), .B(new_n568), .C1(new_n560), .C2(new_n561), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT35), .B1(new_n569), .B2(new_n523), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n564), .A2(new_n552), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(new_n522), .A3(new_n568), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n258), .B1(new_n567), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(G71gat), .ZN(new_n577));
  INV_X1    g376(.A(G78gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n576), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n583), .A3(new_n576), .ZN(new_n584));
  AND2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT95), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G57gat), .ZN(new_n588));
  INV_X1    g387(.A(G64gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G57gat), .A2(G64gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT94), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(G57gat), .A2(G64gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(G57gat), .A2(G64gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n595), .B1(new_n598), .B2(KEYINPUT94), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n582), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n607), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n609), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n232), .B1(new_n601), .B2(new_n600), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT96), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT98), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G99gat), .B(G106gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT8), .ZN(new_n631));
  NAND2_X1  g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT99), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(G99gat), .A3(G106gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n625), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT8), .ZN(new_n639));
  INV_X1    g438(.A(new_n629), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n627), .B2(new_n626), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(new_n641), .A3(new_n624), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n222), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n218), .B2(new_n643), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n623), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n630), .A2(new_n636), .A3(new_n625), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n624), .B1(new_n639), .B2(new_n641), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n220), .B2(new_n221), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n653), .A2(new_n647), .A3(new_n622), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT97), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n649), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n644), .A2(new_n648), .A3(new_n623), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n622), .B1(new_n653), .B2(new_n647), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n621), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n656), .B1(new_n649), .B2(new_n654), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(new_n660), .A3(new_n658), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n620), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n618), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G230gat), .A2(G233gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n600), .B1(new_n650), .B2(new_n651), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n594), .B1(new_n580), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n673), .A2(new_n584), .A3(new_n592), .A4(new_n587), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(new_n582), .A3(new_n642), .A4(new_n637), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n600), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n652), .A2(new_n678), .A3(KEYINPUT10), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n670), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n671), .A2(new_n675), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n670), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(G120gat), .B(G148gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT100), .ZN(new_n686));
  XOR2_X1   g485(.A(G176gat), .B(G204gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n681), .A2(new_n683), .A3(new_n688), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n668), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n575), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n520), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT101), .B(G1gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1324gat));
  INV_X1    g497(.A(new_n490), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n700), .B(KEYINPUT102), .Z(new_n703));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(G8gat), .ZN(new_n705));
  OAI221_X1 g504(.A(new_n702), .B1(KEYINPUT42), .B2(new_n701), .C1(new_n703), .C2(new_n705), .ZN(G1325gat));
  INV_X1    g505(.A(new_n695), .ZN(new_n707));
  AOI21_X1  g506(.A(G15gat), .B1(new_n707), .B2(new_n571), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n562), .A2(new_n565), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G15gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT103), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n707), .B2(new_n711), .ZN(G1326gat));
  NOR2_X1   g511(.A1(new_n695), .A2(new_n568), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT43), .B(G22gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  NAND2_X1  g514(.A1(new_n523), .A2(new_n341), .ZN(new_n716));
  INV_X1    g515(.A(new_n519), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT87), .B1(new_n518), .B2(new_n491), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT104), .B1(new_n719), .B2(new_n709), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n516), .A2(new_n519), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n566), .A4(new_n716), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n720), .A2(new_n574), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n724), .B2(new_n666), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n567), .A2(new_n574), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n667), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n618), .A2(new_n693), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n257), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n520), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n575), .A2(new_n666), .A3(new_n732), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n203), .A3(new_n521), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(G1328gat));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n204), .A3(new_n490), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n739), .A2(new_n740), .A3(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n739), .B2(KEYINPUT46), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n741), .A2(new_n742), .B1(new_n739), .B2(KEYINPUT46), .ZN(new_n743));
  OAI21_X1  g542(.A(G36gat), .B1(new_n733), .B2(new_n699), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1329gat));
  NAND2_X1  g544(.A1(new_n709), .A2(G43gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n733), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(G43gat), .B1(new_n735), .B2(new_n571), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT47), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  INV_X1    g549(.A(new_n748), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n750), .B(new_n751), .C1(new_n733), .C2(new_n746), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1330gat));
  NAND2_X1  g552(.A1(new_n341), .A2(G50gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n733), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n735), .A2(new_n341), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(G50gat), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT48), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  OAI221_X1 g558(.A(new_n759), .B1(G50gat), .B2(new_n756), .C1(new_n733), .C2(new_n754), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1331gat));
  NOR2_X1   g560(.A1(new_n668), .A2(new_n257), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n724), .A2(new_n693), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n520), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n588), .ZN(G1332gat));
  INV_X1    g564(.A(new_n763), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n490), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  AND2_X1   g567(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n768), .B2(new_n767), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n763), .B2(new_n566), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n571), .A2(new_n577), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g574(.A1(new_n763), .A2(new_n568), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n578), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n618), .A2(new_n257), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n692), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n725), .A2(new_n730), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G85gat), .B1(new_n783), .B2(new_n520), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n723), .A2(new_n574), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n722), .B1(new_n524), .B2(new_n566), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n666), .B(new_n778), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n724), .A2(KEYINPUT51), .A3(new_n666), .A4(new_n778), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n520), .A2(G85gat), .A3(new_n692), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT106), .Z(new_n794));
  OAI21_X1  g593(.A(new_n784), .B1(new_n792), .B2(new_n794), .ZN(G1336gat));
  AND2_X1   g594(.A1(new_n490), .A2(G92gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n731), .A2(new_n780), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n699), .A2(new_n692), .ZN(new_n802));
  AOI21_X1  g601(.A(G92gat), .B1(new_n791), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n798), .A2(new_n799), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n804), .ZN(new_n806));
  INV_X1    g605(.A(new_n803), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n782), .A2(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n805), .A2(new_n809), .ZN(G1337gat));
  OAI21_X1  g609(.A(G99gat), .B1(new_n783), .B2(new_n566), .ZN(new_n811));
  INV_X1    g610(.A(new_n571), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n812), .A2(G99gat), .A3(new_n692), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT108), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n792), .B2(new_n814), .ZN(G1338gat));
  INV_X1    g614(.A(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n782), .B2(new_n341), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n568), .A2(G106gat), .A3(new_n692), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT109), .B1(new_n791), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n820));
  INV_X1    g619(.A(new_n818), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n820), .B(new_n821), .C1(new_n789), .C2(new_n790), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n817), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n724), .A2(new_n666), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n727), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n341), .A3(new_n729), .A4(new_n780), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n782), .A2(KEYINPUT110), .A3(new_n341), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n816), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n824), .B1(new_n792), .B2(new_n821), .ZN(new_n832));
  OAI22_X1  g631(.A1(new_n823), .A2(new_n824), .B1(new_n831), .B2(new_n832), .ZN(G1339gat));
  INV_X1    g632(.A(new_n617), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n615), .B(new_n834), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n677), .A2(new_n679), .A3(new_n670), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(new_n680), .A3(new_n837), .ZN(new_n838));
  AOI211_X1 g637(.A(KEYINPUT54), .B(new_n670), .C1(new_n677), .C2(new_n679), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT111), .B1(new_n839), .B2(new_n688), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n677), .A2(new_n679), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n837), .A3(new_n669), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n689), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n838), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n691), .B1(new_n845), .B2(KEYINPUT55), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n847), .B(new_n838), .C1(new_n844), .C2(new_n840), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT112), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n838), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n839), .A2(KEYINPUT111), .A3(new_n688), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n843), .B1(new_n842), .B2(new_n689), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n847), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n850), .B(KEYINPUT55), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n691), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n849), .A2(new_n257), .A3(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n244), .A2(new_n245), .A3(new_n243), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n234), .B1(new_n233), .B2(new_n237), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n252), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n693), .A2(new_n256), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n666), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n256), .A2(new_n861), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT113), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n256), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n865), .A2(new_n666), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(new_n849), .A3(new_n857), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n835), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n618), .A2(new_n258), .A3(new_n667), .A4(new_n692), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT114), .B1(new_n872), .B2(new_n568), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n874));
  AOI211_X1 g673(.A(new_n874), .B(new_n341), .C1(new_n870), .C2(new_n871), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n520), .A2(new_n490), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n812), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G113gat), .B1(new_n880), .B2(new_n258), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n878), .B1(new_n870), .B2(new_n871), .ZN(new_n882));
  INV_X1    g681(.A(new_n569), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n258), .A2(new_n359), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(G1340gat));
  INV_X1    g685(.A(new_n880), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n692), .A2(new_n350), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n883), .A3(new_n693), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n887), .A2(new_n888), .B1(new_n350), .B2(new_n889), .ZN(G1341gat));
  OAI21_X1  g689(.A(new_n348), .B1(new_n880), .B2(new_n835), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n835), .A2(new_n348), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n884), .B2(new_n892), .ZN(G1342gat));
  NAND4_X1  g692(.A1(new_n882), .A2(new_n357), .A3(new_n883), .A4(new_n666), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT115), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n887), .A2(new_n666), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(new_n357), .ZN(G1343gat));
  NOR2_X1   g698(.A1(new_n709), .A2(new_n568), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n882), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n262), .B1(new_n901), .B2(new_n258), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n862), .B(KEYINPUT116), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n258), .A2(new_n848), .A3(new_n846), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n667), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n869), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n618), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n871), .B1(new_n907), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n341), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT57), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n709), .A2(new_n878), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n872), .A2(new_n341), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n912), .B(new_n913), .C1(KEYINPUT57), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n257), .A2(G141gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n902), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g717(.A(new_n901), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n263), .A3(new_n693), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n915), .A2(new_n692), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(KEYINPUT59), .A3(new_n263), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n666), .A2(new_n691), .A3(new_n856), .A4(new_n854), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT118), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(KEYINPUT118), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n925), .A2(new_n865), .A3(new_n867), .A4(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n618), .B1(new_n905), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n871), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n568), .A2(KEYINPUT57), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n930), .A2(new_n931), .B1(new_n914), .B2(KEYINPUT57), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n693), .A3(new_n913), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n923), .B1(new_n933), .B2(G148gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n920), .B1(new_n922), .B2(new_n934), .ZN(G1345gat));
  OAI21_X1  g734(.A(G155gat), .B1(new_n915), .B2(new_n835), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n272), .A3(new_n618), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n915), .B2(new_n667), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n273), .A3(new_n666), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n521), .A2(new_n699), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n872), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(new_n883), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n419), .A3(new_n257), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT119), .Z(new_n946));
  AND2_X1   g745(.A1(new_n571), .A2(new_n942), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n876), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n258), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n946), .A2(new_n950), .ZN(G1348gat));
  OAI21_X1  g750(.A(G176gat), .B1(new_n949), .B2(new_n692), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n944), .A2(new_n420), .A3(new_n693), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  NAND2_X1  g753(.A1(new_n948), .A2(new_n618), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n618), .A2(new_n447), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n955), .A2(G183gat), .B1(new_n944), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g756(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n959), .B(new_n960), .Z(G1350gat));
  OAI211_X1 g760(.A(new_n666), .B(new_n947), .C1(new_n873), .C2(new_n875), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G190gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT121), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n966), .A3(G190gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n964), .A2(KEYINPUT122), .A3(new_n965), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n964), .A2(new_n967), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n944), .A2(new_n448), .A3(new_n666), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n974), .A2(KEYINPUT123), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1351gat));
  AND2_X1   g779(.A1(new_n566), .A2(new_n942), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n932), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(G197gat), .B1(new_n982), .B2(new_n258), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n900), .A2(new_n943), .ZN(new_n984));
  INV_X1    g783(.A(G197gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n984), .A2(new_n985), .A3(new_n257), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n983), .A2(new_n986), .ZN(G1352gat));
  INV_X1    g786(.A(G204gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n984), .A2(new_n988), .A3(new_n693), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n932), .A2(new_n693), .A3(new_n981), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G204gat), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(KEYINPUT125), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n991), .A2(new_n997), .A3(new_n993), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n996), .A2(new_n998), .ZN(G1353gat));
  NAND4_X1  g798(.A1(new_n984), .A2(new_n286), .A3(new_n287), .A4(new_n618), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n932), .A2(new_n1001), .A3(new_n618), .A4(new_n981), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1002), .A2(G211gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(KEYINPUT126), .B1(new_n982), .B2(new_n835), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT63), .ZN(new_n1006));
  OAI21_X1  g805(.A(KEYINPUT127), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n1006), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(G1354gat));
  OAI21_X1  g810(.A(G218gat), .B1(new_n982), .B2(new_n667), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n984), .A2(new_n285), .A3(new_n666), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1012), .A2(new_n1013), .ZN(G1355gat));
endmodule


