//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT65), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n466), .B1(new_n471), .B2(G2104), .ZN(new_n472));
  AOI211_X1 g047(.A(new_n465), .B(new_n463), .C1(new_n468), .C2(new_n470), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n462), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n478), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n479), .A2(new_n462), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  AOI21_X1  g057(.A(KEYINPUT66), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT65), .B(KEYINPUT3), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(new_n463), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n471), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n462), .B1(new_n485), .B2(new_n486), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT67), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(KEYINPUT67), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n467), .A2(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n464), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n462), .A3(G138), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n462), .A2(G138), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n478), .A2(KEYINPUT68), .A3(new_n502), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n506), .B1(new_n472), .B2(new_n473), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n510));
  OAI211_X1 g085(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n511));
  OAI21_X1  g086(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n512));
  INV_X1    g087(.A(G114), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(G2105), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n510), .A2(new_n516), .ZN(G164));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G651), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n519), .A2(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n521), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n523), .A2(G543), .A3(new_n524), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G50), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND2_X1  g109(.A1(new_n531), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n526), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n535), .B(new_n536), .C1(new_n540), .C2(KEYINPUT70), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n540), .A2(KEYINPUT70), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n527), .A2(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n521), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n531), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n527), .A2(G81), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n521), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT71), .B(G43), .Z(new_n553));
  NAND2_X1  g128(.A1(new_n531), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT72), .Z(G188));
  AOI22_X1  g137(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n563), .A2(KEYINPUT73), .A3(new_n521), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT73), .B1(new_n563), .B2(new_n521), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G91), .B2(new_n527), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n523), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n566), .A2(KEYINPUT74), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT74), .B1(new_n566), .B2(new_n568), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  NAND2_X1  g147(.A1(new_n527), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n531), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n521), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT75), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n523), .A2(G86), .A3(new_n524), .A4(new_n525), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n523), .A2(G48), .A3(G543), .A4(new_n524), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n577), .B2(new_n521), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n531), .A2(G47), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT76), .B(G85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n526), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT77), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n521), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n527), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT10), .Z(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(new_n525), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n531), .A2(G54), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  XOR2_X1   g183(.A(KEYINPUT78), .B(G559), .Z(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(G860), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT79), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n487), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n489), .A2(G123), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  INV_X1    g194(.A(G111), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(G2105), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n619), .B2(new_n618), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n616), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n478), .A2(new_n475), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT13), .B(G2100), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n625), .A3(new_n630), .ZN(G156));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n637), .A2(new_n641), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OR3_X1    g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n651), .A2(new_n652), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n659), .B(new_n663), .Z(G227));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OR3_X1    g252(.A1(new_n667), .A2(new_n670), .A3(new_n674), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G229));
  NAND2_X1  g262(.A1(new_n489), .A2(G119), .ZN(new_n688));
  OR2_X1    g263(.A1(G95), .A2(G2105), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n689), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n487), .A2(G131), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT87), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G25), .B2(new_n696), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  MUX2_X1   g276(.A(G24), .B(G290), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G23), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT88), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G288), .B2(new_n705), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT33), .B(G1976), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G6), .B(G305), .S(G16), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n710), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n708), .A2(new_n709), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT34), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OR3_X1    g296(.A1(new_n719), .A2(KEYINPUT34), .A3(new_n720), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n704), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT36), .Z(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G35), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G162), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2090), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G4), .A2(G16), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n602), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT90), .B(G1348), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n705), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n705), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G171), .A2(new_n705), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G5), .B2(new_n705), .ZN(new_n740));
  INV_X1    g315(.A(G1961), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G19), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n556), .B2(G16), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n740), .A2(new_n741), .B1(G1341), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G1341), .B2(new_n743), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT93), .B(G28), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(new_n696), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n746), .B1(new_n748), .B2(new_n750), .C1(new_n623), .C2(new_n696), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n740), .B2(new_n741), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n696), .A2(G33), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n487), .A2(G139), .ZN(new_n754));
  NAND2_X1  g329(.A1(G115), .A2(G2104), .ZN(new_n755));
  INV_X1    g330(.A(G127), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n501), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n758));
  NAND2_X1  g333(.A1(G103), .A2(G2104), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G2105), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n757), .A2(G2105), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n753), .B1(new_n764), .B2(new_n696), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G2072), .Z(new_n766));
  NAND3_X1  g341(.A1(new_n745), .A2(new_n752), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n696), .B1(KEYINPUT24), .B2(G34), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(KEYINPUT24), .B2(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n481), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G27), .A2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G164), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2078), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n738), .A2(new_n767), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n696), .A2(G26), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT28), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n487), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n489), .A2(G128), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n778), .B1(new_n789), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2067), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n489), .A2(G129), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT26), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n795), .A2(new_n796), .B1(G105), .B2(new_n475), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n487), .A2(G141), .ZN(new_n799));
  AOI21_X1  g374(.A(KEYINPUT92), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(KEYINPUT92), .A3(new_n799), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G32), .B(new_n803), .S(G29), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT27), .B(G1996), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n705), .A2(G20), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT23), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n606), .B2(new_n705), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT95), .B(G1956), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n729), .A2(new_n776), .A3(new_n791), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n724), .A2(new_n813), .ZN(G311));
  OR2_X1    g389(.A1(new_n724), .A2(new_n813), .ZN(G150));
  NAND2_X1  g390(.A1(G80), .A2(G543), .ZN(new_n816));
  INV_X1    g391(.A(G67), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n597), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT97), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(new_n816), .C1(new_n597), .C2(new_n817), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(G651), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT98), .B(G55), .ZN(new_n823));
  AOI22_X1  g398(.A1(G93), .A2(new_n527), .B1(new_n531), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n602), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n556), .A2(new_n822), .A3(new_n824), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n825), .A2(new_n555), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n830), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n827), .B1(new_n836), .B2(new_n838), .ZN(G145));
  INV_X1    g414(.A(G164), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n788), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(G164), .B1(new_n786), .B2(new_n787), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n763), .B1(new_n801), .B2(new_n802), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n798), .A2(new_n799), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n764), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n802), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n764), .B1(new_n847), .B2(new_n800), .ZN(new_n848));
  INV_X1    g423(.A(new_n845), .ZN(new_n849));
  INV_X1    g424(.A(new_n787), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n840), .B1(new_n850), .B2(new_n785), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n786), .A2(new_n787), .A3(G164), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n848), .B(new_n849), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n487), .A2(G142), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n489), .B2(G130), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n693), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n856), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n691), .A2(new_n862), .A3(new_n692), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n628), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n628), .B1(new_n861), .B2(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n855), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n854), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n477), .A2(KEYINPUT99), .A3(new_n480), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT99), .B1(new_n477), .B2(new_n480), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n497), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n495), .B(new_n496), .C1(new_n870), .C2(new_n871), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n623), .ZN(new_n876));
  INV_X1    g451(.A(new_n623), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n877), .A3(new_n874), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n864), .B(new_n865), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n880), .A2(new_n846), .A3(new_n855), .A4(new_n853), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n869), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT101), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n869), .A2(new_n879), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n866), .A2(new_n867), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n854), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n879), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g467(.A1(new_n825), .A2(G868), .ZN(new_n893));
  INV_X1    g468(.A(G288), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n589), .A2(new_n894), .A3(new_n591), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n589), .B2(new_n591), .ZN(new_n897));
  XNOR2_X1  g472(.A(G166), .B(G305), .ZN(new_n898));
  OR4_X1    g473(.A1(KEYINPUT103), .A2(new_n896), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT103), .B1(new_n896), .B2(new_n897), .ZN(new_n900));
  INV_X1    g475(.A(new_n897), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n895), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n903), .A3(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n569), .B2(new_n570), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n566), .A2(new_n568), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT74), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n566), .A2(KEYINPUT74), .A3(new_n568), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(KEYINPUT102), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n916), .A3(new_n602), .ZN(new_n917));
  NAND3_X1  g492(.A1(G299), .A2(KEYINPUT102), .A3(new_n601), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n612), .B(new_n833), .Z(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n919), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT105), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n909), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n925), .A2(KEYINPUT105), .A3(new_n927), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n893), .B1(new_n931), .B2(G868), .ZN(G295));
  AOI21_X1  g507(.A(new_n893), .B1(new_n931), .B2(G868), .ZN(G331));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n831), .A2(new_n832), .A3(G301), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G301), .B1(new_n831), .B2(new_n832), .ZN(new_n937));
  OAI21_X1  g512(.A(G286), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n937), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(G168), .A3(new_n935), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n921), .A2(new_n941), .A3(new_n922), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n926), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n945), .B2(new_n905), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n942), .A2(new_n899), .A3(new_n904), .A4(new_n944), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n947), .B1(new_n946), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n934), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n945), .A2(new_n905), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n948), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n949), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT106), .A3(new_n934), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n949), .A2(KEYINPUT107), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n946), .A2(new_n962), .A3(new_n947), .A4(new_n948), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n961), .A2(KEYINPUT44), .A3(new_n958), .A4(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n954), .A2(new_n960), .A3(new_n964), .ZN(G397));
  INV_X1    g540(.A(G2067), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n788), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n844), .A2(G1996), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n803), .B2(G1996), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n510), .B2(new_n516), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT109), .B(G40), .Z(new_n975));
  NAND4_X1  g550(.A1(new_n474), .A2(new_n480), .A3(new_n476), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n970), .A2(KEYINPUT111), .A3(new_n977), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n693), .B(new_n699), .Z(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n977), .ZN(new_n983));
  OR2_X1    g558(.A1(G290), .A2(G1986), .ZN(new_n984));
  NAND2_X1  g559(.A1(G290), .A2(G1986), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT110), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n977), .C1(KEYINPUT110), .C2(new_n985), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n980), .A2(new_n981), .A3(new_n983), .A4(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT112), .Z(new_n989));
  INV_X1    g564(.A(G1981), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT117), .B1(new_n580), .B2(new_n581), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n578), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n582), .A2(KEYINPUT117), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n990), .A2(new_n579), .A3(new_n582), .A4(new_n584), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT49), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(KEYINPUT49), .C1(new_n994), .C2(new_n995), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n504), .A2(new_n507), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n505), .B1(new_n485), .B2(new_n486), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n502), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n514), .B1(new_n489), .B2(G126), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n976), .ZN(new_n1007));
  AOI211_X1 g582(.A(KEYINPUT116), .B(new_n1001), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(G8), .ZN(new_n1011));
  OAI22_X1  g586(.A1(new_n998), .A2(new_n1000), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n894), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1014), .A2(new_n995), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n894), .A2(G1976), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n1011), .B2(new_n1008), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT52), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1016), .B(new_n1019), .C1(new_n1011), .C2(new_n1008), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1018), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1023), .A2(KEYINPUT115), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT45), .B(new_n971), .C1(new_n510), .C2(new_n516), .ZN(new_n1029));
  INV_X1    g604(.A(new_n973), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1029), .B(new_n1007), .C1(new_n1006), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1971), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(KEYINPUT113), .A3(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n972), .A2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n971), .C1(new_n510), .C2(new_n516), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n972), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n1043));
  AOI211_X1 g618(.A(G2090), .B(new_n976), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(G8), .B(new_n1028), .C1(new_n1037), .C2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1015), .B1(new_n1022), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n976), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n771), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n976), .B1(new_n972), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1006), .A2(new_n1030), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n736), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1054), .A2(G8), .A3(G168), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT63), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1028), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1057), .A2(new_n1045), .A3(new_n1021), .A4(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1007), .B1(new_n1006), .B2(new_n1040), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1041), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1062), .A2(new_n1063), .A3(G2090), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1059), .B1(new_n1065), .B2(new_n1001), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1021), .A2(new_n1045), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1056), .B1(new_n1067), .B2(new_n1055), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1046), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n974), .A2(new_n1007), .A3(new_n1029), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n976), .B1(new_n972), .B2(KEYINPUT50), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1956), .B1(new_n1073), .B2(new_n1041), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT120), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1956), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n1071), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n912), .A2(KEYINPUT57), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n566), .B2(new_n568), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1075), .A2(new_n1079), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT121), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1075), .A2(new_n1079), .A3(new_n1087), .A4(new_n1084), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1006), .A2(new_n1007), .A3(new_n966), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1047), .B2(G1348), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n602), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1077), .A2(new_n1071), .A3(new_n1083), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1077), .A2(new_n1083), .A3(KEYINPUT119), .A4(new_n1071), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1089), .A2(new_n1092), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1996), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n974), .A2(new_n1098), .A3(new_n1007), .A4(new_n1029), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1010), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(KEYINPUT122), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT122), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n556), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT59), .B(new_n556), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1083), .B1(new_n1077), .B2(new_n1071), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1106), .B(new_n1107), .C1(new_n1109), .C2(KEYINPUT61), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n602), .B1(new_n1091), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1041), .A2(new_n1039), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1006), .A2(new_n1040), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1043), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1007), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1348), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n601), .A4(new_n1090), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1112), .A2(new_n1120), .B1(new_n1111), .B2(new_n1091), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1110), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1089), .A2(KEYINPUT61), .A3(new_n1093), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1097), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1117), .A2(new_n741), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1031), .B2(G2078), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n477), .A2(KEYINPUT124), .ZN(new_n1128));
  INV_X1    g703(.A(G2078), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n480), .A2(KEYINPUT53), .A3(G40), .A4(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n477), .A2(KEYINPUT124), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n974), .A3(new_n1029), .A4(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1125), .A2(G301), .A3(new_n1127), .A4(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1050), .A2(KEYINPUT53), .A3(new_n1129), .A4(new_n1051), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(new_n1127), .C1(new_n1047), .C2(G1961), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT54), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n1067), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1031), .A2(G2078), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1117), .A2(new_n741), .B1(new_n1140), .B2(new_n1126), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1141), .A2(KEYINPUT125), .A3(G301), .A4(new_n1135), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1136), .B2(G171), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n1133), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G171), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(KEYINPUT54), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  AOI211_X1 g724(.A(G2084), .B(new_n976), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1053), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1048), .A2(KEYINPUT123), .A3(new_n1053), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G168), .A2(new_n1001), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1152), .A2(new_n1153), .A3(G168), .ZN(new_n1157));
  AND2_X1   g732(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1054), .A2(G8), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1155), .A2(KEYINPUT51), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1157), .A2(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1139), .B(new_n1148), .C1(new_n1156), .C2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1069), .B1(new_n1124), .B2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1067), .A2(new_n1137), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1161), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1156), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(KEYINPUT62), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1161), .B2(new_n1156), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1164), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n989), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n977), .B1(new_n967), .B2(new_n844), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT126), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n977), .A2(new_n1098), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT46), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT47), .ZN(new_n1177));
  AND4_X1   g752(.A1(new_n695), .A2(new_n980), .A3(new_n699), .A4(new_n981), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n789), .A2(G2067), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n977), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n984), .A2(new_n976), .A3(new_n974), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT48), .Z(new_n1182));
  NAND4_X1  g757(.A1(new_n1182), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1177), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1171), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1187));
  NOR3_X1   g761(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1188), .B1(new_n685), .B2(new_n686), .ZN(new_n1189));
  AOI21_X1  g763(.A(new_n1189), .B1(new_n886), .B2(new_n890), .ZN(new_n1190));
  OAI211_X1 g764(.A(new_n1187), .B(new_n1190), .C1(new_n950), .C2(new_n951), .ZN(new_n1191));
  INV_X1    g765(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1187), .B1(new_n959), .B2(new_n1190), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n1192), .A2(new_n1193), .ZN(G308));
  NAND2_X1  g768(.A1(new_n959), .A2(new_n1190), .ZN(G225));
endmodule


