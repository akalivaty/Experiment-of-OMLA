

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U553 ( .A1(n777), .A2(n778), .ZN(n725) );
  NOR2_X1 U554 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U555 ( .A(n725), .B(KEYINPUT92), .ZN(n692) );
  NOR2_X1 U556 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U557 ( .A1(n875), .A2(G137), .ZN(n520) );
  INV_X1 U558 ( .A(n725), .ZN(n679) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n708) );
  XNOR2_X1 U560 ( .A(n709), .B(n708), .ZN(n733) );
  OR2_X1 U561 ( .A1(n724), .A2(n723), .ZN(n740) );
  INV_X1 U562 ( .A(KEYINPUT17), .ZN(n518) );
  NOR2_X1 U563 ( .A1(G651), .A2(n632), .ZN(n639) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n527), .Z(n643) );
  AND2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U566 ( .A1(n883), .A2(G113), .ZN(n517) );
  XNOR2_X1 U567 ( .A(n517), .B(KEYINPUT64), .ZN(n521) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XNOR2_X2 U569 ( .A(n519), .B(n518), .ZN(n875) );
  NAND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U571 ( .A(n522), .B(KEYINPUT65), .ZN(n524) );
  INV_X1 U572 ( .A(G2104), .ZN(n525) );
  AND2_X1 U573 ( .A1(n525), .A2(G2105), .ZN(n882) );
  NAND2_X1 U574 ( .A1(G125), .A2(n882), .ZN(n523) );
  AND2_X1 U575 ( .A1(n524), .A2(n523), .ZN(n672) );
  NOR2_X2 U576 ( .A1(G2105), .A2(n525), .ZN(n877) );
  NAND2_X1 U577 ( .A1(G101), .A2(n877), .ZN(n526) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n526), .Z(n671) );
  AND2_X1 U579 ( .A1(n672), .A2(n671), .ZN(G160) );
  XOR2_X1 U580 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  NAND2_X1 U581 ( .A1(G52), .A2(n639), .ZN(n529) );
  INV_X1 U582 ( .A(G651), .ZN(n530) );
  NOR2_X1 U583 ( .A1(G543), .A2(n530), .ZN(n527) );
  NAND2_X1 U584 ( .A1(G64), .A2(n643), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n635) );
  NAND2_X1 U587 ( .A1(G90), .A2(n635), .ZN(n532) );
  NOR2_X1 U588 ( .A1(n632), .A2(n530), .ZN(n636) );
  NAND2_X1 U589 ( .A1(G77), .A2(n636), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U591 ( .A(KEYINPUT9), .B(n533), .Z(n534) );
  NOR2_X1 U592 ( .A1(n535), .A2(n534), .ZN(G171) );
  INV_X1 U593 ( .A(G57), .ZN(G237) );
  INV_X1 U594 ( .A(G82), .ZN(G220) );
  NAND2_X1 U595 ( .A1(G138), .A2(n875), .ZN(n537) );
  NAND2_X1 U596 ( .A1(G102), .A2(n877), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G126), .A2(n882), .ZN(n539) );
  NAND2_X1 U599 ( .A1(G114), .A2(n883), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U602 ( .A1(n636), .A2(G76), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT76), .B(n542), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n635), .A2(G89), .ZN(n543) );
  XNOR2_X1 U605 ( .A(KEYINPUT4), .B(n543), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G51), .A2(n639), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G63), .A2(n643), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U613 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U614 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U615 ( .A1(G94), .A2(G452), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n553), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U617 ( .A1(G7), .A2(G661), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U619 ( .A(G223), .ZN(n822) );
  NAND2_X1 U620 ( .A1(n822), .A2(G567), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  NAND2_X1 U622 ( .A1(n643), .A2(G56), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT14), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G43), .A2(n639), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n635), .A2(G81), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U628 ( .A1(G68), .A2(n636), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(KEYINPUT71), .B(n562), .ZN(n563) );
  XNOR2_X1 U631 ( .A(KEYINPUT13), .B(n563), .ZN(n564) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n923) );
  NAND2_X1 U633 ( .A1(n923), .A2(G860), .ZN(G153) );
  XOR2_X1 U634 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  INV_X1 U635 ( .A(G868), .ZN(n593) );
  NOR2_X1 U636 ( .A1(G301), .A2(n593), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G54), .A2(n639), .ZN(n567) );
  NAND2_X1 U638 ( .A1(G79), .A2(n636), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n567), .A2(n566), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G92), .A2(n635), .ZN(n569) );
  NAND2_X1 U641 ( .A1(G66), .A2(n643), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U643 ( .A(n570), .B(KEYINPUT73), .Z(n571) );
  NOR2_X1 U644 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U645 ( .A(KEYINPUT15), .B(n573), .Z(n574) );
  XOR2_X1 U646 ( .A(KEYINPUT74), .B(n574), .Z(n687) );
  INV_X1 U647 ( .A(n687), .ZN(n605) );
  INV_X1 U648 ( .A(n605), .ZN(n934) );
  NOR2_X1 U649 ( .A1(n934), .A2(G868), .ZN(n575) );
  NOR2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U651 ( .A(KEYINPUT75), .B(n577), .Z(G284) );
  NAND2_X1 U652 ( .A1(G91), .A2(n635), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G78), .A2(n636), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n584) );
  NAND2_X1 U655 ( .A1(G53), .A2(n639), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G65), .A2(n643), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U658 ( .A(KEYINPUT68), .B(n582), .ZN(n583) );
  NOR2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U660 ( .A(n585), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U661 ( .A1(G286), .A2(G868), .ZN(n587) );
  NAND2_X1 U662 ( .A1(G299), .A2(n593), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(G297) );
  INV_X1 U664 ( .A(G860), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n588), .A2(G559), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n589), .A2(n605), .ZN(n590) );
  XNOR2_X1 U667 ( .A(n590), .B(KEYINPUT16), .ZN(n591) );
  XOR2_X1 U668 ( .A(KEYINPUT77), .B(n591), .Z(G148) );
  NAND2_X1 U669 ( .A1(G868), .A2(n605), .ZN(n592) );
  NOR2_X1 U670 ( .A1(G559), .A2(n592), .ZN(n595) );
  AND2_X1 U671 ( .A1(n593), .A2(n923), .ZN(n594) );
  NOR2_X1 U672 ( .A1(n595), .A2(n594), .ZN(G282) );
  XOR2_X1 U673 ( .A(G2100), .B(KEYINPUT78), .Z(n604) );
  NAND2_X1 U674 ( .A1(n882), .A2(G123), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT18), .ZN(n598) );
  NAND2_X1 U676 ( .A1(G111), .A2(n883), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G135), .A2(n875), .ZN(n600) );
  NAND2_X1 U679 ( .A1(G99), .A2(n877), .ZN(n599) );
  NAND2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n1011) );
  XNOR2_X1 U682 ( .A(n1011), .B(G2096), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(G156) );
  NAND2_X1 U684 ( .A1(n605), .A2(G559), .ZN(n606) );
  XOR2_X1 U685 ( .A(n923), .B(n606), .Z(n654) );
  NOR2_X1 U686 ( .A1(n654), .A2(G860), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G55), .A2(n639), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G67), .A2(n643), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G93), .A2(n635), .ZN(n610) );
  NAND2_X1 U691 ( .A1(G80), .A2(n636), .ZN(n609) );
  NAND2_X1 U692 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n652) );
  XNOR2_X1 U694 ( .A(n613), .B(n652), .ZN(G145) );
  NAND2_X1 U695 ( .A1(G73), .A2(n636), .ZN(n614) );
  XNOR2_X1 U696 ( .A(n614), .B(KEYINPUT2), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G86), .A2(n635), .ZN(n616) );
  NAND2_X1 U698 ( .A1(G61), .A2(n643), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G48), .A2(n639), .ZN(n617) );
  XNOR2_X1 U701 ( .A(KEYINPUT79), .B(n617), .ZN(n618) );
  NOR2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(G305) );
  NAND2_X1 U704 ( .A1(G85), .A2(n635), .ZN(n623) );
  NAND2_X1 U705 ( .A1(G72), .A2(n636), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U707 ( .A1(G47), .A2(n639), .ZN(n624) );
  XOR2_X1 U708 ( .A(KEYINPUT66), .B(n624), .Z(n625) );
  NOR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n643), .A2(G60), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(G290) );
  NAND2_X1 U712 ( .A1(G49), .A2(n639), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U715 ( .A1(n643), .A2(n631), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G88), .A2(n635), .ZN(n638) );
  NAND2_X1 U719 ( .A1(G75), .A2(n636), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n639), .A2(G50), .ZN(n640) );
  XOR2_X1 U722 ( .A(KEYINPUT80), .B(n640), .Z(n641) );
  NOR2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n643), .A2(G62), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(G303) );
  NOR2_X1 U726 ( .A1(G868), .A2(n652), .ZN(n646) );
  XOR2_X1 U727 ( .A(n646), .B(KEYINPUT82), .Z(n657) );
  XOR2_X1 U728 ( .A(G290), .B(G299), .Z(n647) );
  XNOR2_X1 U729 ( .A(G305), .B(n647), .ZN(n648) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(n648), .ZN(n650) );
  XNOR2_X1 U731 ( .A(G288), .B(KEYINPUT81), .ZN(n649) );
  XNOR2_X1 U732 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(n653), .B(G303), .ZN(n898) );
  XNOR2_X1 U735 ( .A(n898), .B(n654), .ZN(n655) );
  NAND2_X1 U736 ( .A1(G868), .A2(n655), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n658) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U744 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U745 ( .A1(G219), .A2(G220), .ZN(n662) );
  XOR2_X1 U746 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U747 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U748 ( .A1(G96), .A2(n664), .ZN(n828) );
  NAND2_X1 U749 ( .A1(n828), .A2(G2106), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G69), .A2(G120), .ZN(n665) );
  NOR2_X1 U751 ( .A1(G237), .A2(n665), .ZN(n666) );
  NAND2_X1 U752 ( .A1(G108), .A2(n666), .ZN(n829) );
  NAND2_X1 U753 ( .A1(n829), .A2(G567), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n668), .A2(n667), .ZN(n830) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n669) );
  NOR2_X1 U756 ( .A1(n830), .A2(n669), .ZN(n827) );
  NAND2_X1 U757 ( .A1(n827), .A2(G36), .ZN(n670) );
  XOR2_X1 U758 ( .A(KEYINPUT83), .B(n670), .Z(G176) );
  AND2_X1 U759 ( .A1(G40), .A2(n671), .ZN(n673) );
  AND2_X1 U760 ( .A1(n673), .A2(n672), .ZN(n777) );
  NOR2_X1 U761 ( .A1(G164), .A2(G1384), .ZN(n778) );
  INV_X1 U762 ( .A(G2067), .ZN(n674) );
  OR2_X1 U763 ( .A1(n692), .A2(n674), .ZN(n677) );
  NAND2_X1 U764 ( .A1(G1348), .A2(n725), .ZN(n675) );
  XOR2_X1 U765 ( .A(KEYINPUT93), .B(n675), .Z(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U767 ( .A(n678), .B(KEYINPUT94), .ZN(n686) );
  NAND2_X1 U768 ( .A1(n686), .A2(n687), .ZN(n685) );
  AND2_X1 U769 ( .A1(G1341), .A2(n725), .ZN(n683) );
  NAND2_X1 U770 ( .A1(n679), .A2(G1996), .ZN(n680) );
  XNOR2_X1 U771 ( .A(n680), .B(KEYINPUT26), .ZN(n681) );
  NAND2_X1 U772 ( .A1(n681), .A2(n923), .ZN(n682) );
  NOR2_X1 U773 ( .A1(n683), .A2(n682), .ZN(n684) );
  AND2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U776 ( .A(n690), .B(KEYINPUT95), .ZN(n696) );
  INV_X1 U777 ( .A(n692), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n703), .A2(G2072), .ZN(n691) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(n691), .Z(n694) );
  NAND2_X1 U780 ( .A1(n692), .A2(G1956), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U782 ( .A1(G299), .A2(n698), .ZN(n695) );
  NOR2_X1 U783 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U784 ( .A(n697), .B(KEYINPUT96), .ZN(n701) );
  NAND2_X1 U785 ( .A1(G299), .A2(n698), .ZN(n699) );
  XOR2_X1 U786 ( .A(KEYINPUT28), .B(n699), .Z(n700) );
  XNOR2_X1 U787 ( .A(n702), .B(KEYINPUT29), .ZN(n707) );
  XNOR2_X1 U788 ( .A(G2078), .B(KEYINPUT25), .ZN(n970) );
  NAND2_X1 U789 ( .A1(n703), .A2(n970), .ZN(n705) );
  INV_X1 U790 ( .A(G1961), .ZN(n949) );
  NAND2_X1 U791 ( .A1(n949), .A2(n725), .ZN(n704) );
  NAND2_X1 U792 ( .A1(n705), .A2(n704), .ZN(n714) );
  NAND2_X1 U793 ( .A1(G171), .A2(n714), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U795 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n719) );
  NAND2_X1 U796 ( .A1(G8), .A2(n725), .ZN(n762) );
  NOR2_X1 U797 ( .A1(G1966), .A2(n762), .ZN(n721) );
  NOR2_X1 U798 ( .A1(G2084), .A2(n725), .ZN(n720) );
  NOR2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n710) );
  NAND2_X1 U800 ( .A1(G8), .A2(n710), .ZN(n711) );
  XNOR2_X1 U801 ( .A(KEYINPUT30), .B(n711), .ZN(n712) );
  NOR2_X1 U802 ( .A1(G168), .A2(n712), .ZN(n713) );
  XOR2_X1 U803 ( .A(KEYINPUT98), .B(n713), .Z(n717) );
  NOR2_X1 U804 ( .A1(G171), .A2(n714), .ZN(n715) );
  XNOR2_X1 U805 ( .A(KEYINPUT99), .B(n715), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U807 ( .A(n719), .B(n718), .ZN(n731) );
  AND2_X1 U808 ( .A1(n733), .A2(n731), .ZN(n724) );
  AND2_X1 U809 ( .A1(G8), .A2(n720), .ZN(n722) );
  OR2_X1 U810 ( .A1(n722), .A2(n721), .ZN(n723) );
  INV_X1 U811 ( .A(G8), .ZN(n730) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n762), .ZN(n727) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n725), .ZN(n726) );
  NOR2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n728), .A2(G303), .ZN(n729) );
  OR2_X1 U816 ( .A1(n730), .A2(n729), .ZN(n734) );
  AND2_X1 U817 ( .A1(n731), .A2(n734), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n733), .A2(n732), .ZN(n737) );
  INV_X1 U819 ( .A(n734), .ZN(n735) );
  OR2_X1 U820 ( .A1(n735), .A2(G286), .ZN(n736) );
  NAND2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U822 ( .A(n738), .B(KEYINPUT32), .ZN(n739) );
  NAND2_X1 U823 ( .A1(n740), .A2(n739), .ZN(n757) );
  NOR2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n744) );
  NOR2_X1 U825 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U826 ( .A1(n744), .A2(n741), .ZN(n920) );
  NAND2_X1 U827 ( .A1(n757), .A2(n920), .ZN(n742) );
  XNOR2_X1 U828 ( .A(KEYINPUT101), .B(n742), .ZN(n751) );
  NAND2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n918) );
  INV_X1 U830 ( .A(n762), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n918), .A2(n743), .ZN(n749) );
  NAND2_X1 U832 ( .A1(n744), .A2(KEYINPUT33), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n745), .A2(n762), .ZN(n747) );
  XOR2_X1 U834 ( .A(G1981), .B(G305), .Z(n928) );
  INV_X1 U835 ( .A(n928), .ZN(n746) );
  NOR2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n752) );
  INV_X1 U837 ( .A(n752), .ZN(n748) );
  OR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n754) );
  AND2_X1 U840 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n766) );
  NOR2_X1 U842 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U843 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U845 ( .A(n758), .B(KEYINPUT102), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n759), .A2(n762), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XOR2_X1 U848 ( .A(n760), .B(KEYINPUT24), .Z(n761) );
  OR2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n804) );
  NAND2_X1 U852 ( .A1(G128), .A2(n882), .ZN(n768) );
  NAND2_X1 U853 ( .A1(G116), .A2(n883), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U855 ( .A(n769), .B(KEYINPUT35), .ZN(n774) );
  NAND2_X1 U856 ( .A1(G140), .A2(n875), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G104), .A2(n877), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U859 ( .A(KEYINPUT34), .B(n772), .Z(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U861 ( .A(n775), .B(KEYINPUT36), .Z(n892) );
  XNOR2_X1 U862 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  OR2_X1 U863 ( .A1(n892), .A2(n813), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT85), .ZN(n1007) );
  INV_X1 U865 ( .A(n777), .ZN(n779) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(KEYINPUT84), .ZN(n816) );
  NAND2_X1 U868 ( .A1(n1007), .A2(n816), .ZN(n811) );
  NAND2_X1 U869 ( .A1(G119), .A2(n882), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G107), .A2(n883), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n782), .A2(n781), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n875), .A2(G131), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(KEYINPUT86), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G95), .A2(n877), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U876 ( .A(KEYINPUT87), .B(n786), .Z(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U878 ( .A(KEYINPUT88), .B(n789), .Z(n891) );
  XOR2_X1 U879 ( .A(KEYINPUT89), .B(G1991), .Z(n976) );
  AND2_X1 U880 ( .A1(n891), .A2(n976), .ZN(n790) );
  XNOR2_X1 U881 ( .A(n790), .B(KEYINPUT90), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G141), .A2(n875), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G129), .A2(n882), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G117), .A2(n883), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n877), .A2(G105), .ZN(n793) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U889 ( .A(KEYINPUT91), .B(n796), .Z(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n869) );
  AND2_X1 U891 ( .A1(G1996), .A2(n869), .ZN(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n806) );
  XOR2_X1 U893 ( .A(G1986), .B(G290), .Z(n919) );
  NAND2_X1 U894 ( .A1(n806), .A2(n919), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n801), .A2(n816), .ZN(n802) );
  AND2_X1 U896 ( .A1(n811), .A2(n802), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n819) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n869), .ZN(n805) );
  XOR2_X1 U899 ( .A(KEYINPUT103), .B(n805), .Z(n997) );
  INV_X1 U900 ( .A(n806), .ZN(n1018) );
  NOR2_X1 U901 ( .A1(n891), .A2(n976), .ZN(n1010) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n1010), .A2(n807), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n1018), .A2(n808), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n997), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n813), .A2(n892), .ZN(n1008) );
  NAND2_X1 U909 ( .A1(n814), .A2(n1008), .ZN(n815) );
  XNOR2_X1 U910 ( .A(KEYINPUT104), .B(n815), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n821) );
  XOR2_X1 U913 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n820) );
  XNOR2_X1 U914 ( .A(n821), .B(n820), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n822), .ZN(G217) );
  NAND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n824) );
  INV_X1 U917 ( .A(G661), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n830), .ZN(G319) );
  XOR2_X1 U929 ( .A(G2100), .B(KEYINPUT43), .Z(n832) );
  XNOR2_X1 U930 ( .A(G2090), .B(G2678), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U932 ( .A(n833), .B(KEYINPUT108), .Z(n835) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2096), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n841) );
  XNOR2_X1 U940 ( .A(G1966), .B(G1956), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n842), .B(G2474), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT41), .B(G1981), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1961), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U949 ( .A1(G112), .A2(n883), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n849), .B(KEYINPUT110), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n851) );
  NAND2_X1 U952 ( .A1(G124), .A2(n882), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U955 ( .A1(G136), .A2(n875), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G100), .A2(n877), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U958 ( .A1(n857), .A2(n856), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n859) );
  XNOR2_X1 U960 ( .A(KEYINPUT116), .B(KEYINPUT114), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n868) );
  NAND2_X1 U962 ( .A1(G127), .A2(n882), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G115), .A2(n883), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n862), .B(KEYINPUT47), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G103), .A2(n877), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G139), .A2(n875), .ZN(n865) );
  XNOR2_X1 U969 ( .A(KEYINPUT115), .B(n865), .ZN(n866) );
  NOR2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n1000) );
  XOR2_X1 U971 ( .A(n868), .B(n1000), .Z(n871) );
  XOR2_X1 U972 ( .A(G164), .B(n869), .Z(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n872), .B(G162), .Z(n874) );
  XNOR2_X1 U975 ( .A(G160), .B(n1011), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n890) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n875), .A2(G142), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n876), .B(KEYINPUT112), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G106), .A2(n877), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G130), .A2(n882), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G118), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(KEYINPUT111), .B(n886), .Z(n887) );
  NOR2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(n890), .B(n889), .Z(n894) );
  XOR2_X1 U989 ( .A(n892), .B(n891), .Z(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G395) );
  XOR2_X1 U992 ( .A(G286), .B(n923), .Z(n897) );
  XNOR2_X1 U993 ( .A(G171), .B(n934), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U996 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2443), .B(G2451), .Z(n902) );
  XNOR2_X1 U998 ( .A(G2446), .B(G2454), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n903), .B(G2427), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1003 ( .A(G2435), .B(KEYINPUT106), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G2430), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1006 ( .A(n909), .B(n908), .Z(n910) );
  NAND2_X1 U1007 ( .A1(G14), .A2(n910), .ZN(n916) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G303), .ZN(G166) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n916), .ZN(G401) );
  XNOR2_X1 U1018 ( .A(G16), .B(KEYINPUT56), .ZN(n940) );
  NAND2_X1 U1019 ( .A1(G1971), .A2(G303), .ZN(n917) );
  NAND2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n927) );
  XOR2_X1 U1023 ( .A(n923), .B(G1341), .Z(n925) );
  XOR2_X1 U1024 ( .A(G171), .B(G1961), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G168), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT122), .ZN(n931) );
  XOR2_X1 U1030 ( .A(KEYINPUT57), .B(n931), .Z(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(G299), .B(G1956), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n934), .B(G1348), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n969) );
  INV_X1 U1037 ( .A(G16), .ZN(n967) );
  XNOR2_X1 U1038 ( .A(G1986), .B(G24), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(G1971), .B(G22), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(KEYINPUT124), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(G23), .B(G1976), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(KEYINPUT125), .B(n944), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(KEYINPUT126), .B(n947), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT58), .ZN(n964) );
  XOR2_X1 U1047 ( .A(G1966), .B(G21), .Z(n951) );
  XNOR2_X1 U1048 ( .A(n949), .B(G5), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n962) );
  XNOR2_X1 U1050 ( .A(G1956), .B(G20), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(n952), .B(G4), .ZN(n953) );
  XNOR2_X1 U1053 ( .A(n953), .B(G1348), .ZN(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G1341), .B(G19), .ZN(n957) );
  XNOR2_X1 U1056 ( .A(G1981), .B(G6), .ZN(n956) );
  NOR2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(KEYINPUT60), .B(n960), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1062 ( .A(KEYINPUT61), .B(n965), .Z(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n993) );
  XOR2_X1 U1065 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n990) );
  XNOR2_X1 U1066 ( .A(G2090), .B(G35), .ZN(n985) );
  XNOR2_X1 U1067 ( .A(n970), .B(G27), .ZN(n972) );
  XOR2_X1 U1068 ( .A(G1996), .B(G32), .Z(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(G2067), .B(G26), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(G33), .B(G2072), .ZN(n973) );
  NOR2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(KEYINPUT120), .B(n975), .ZN(n980) );
  XOR2_X1 U1074 ( .A(n976), .B(G25), .Z(n977) );
  NAND2_X1 U1075 ( .A1(n977), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(n978), .B(KEYINPUT119), .ZN(n979) );
  NAND2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT53), .B(n983), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1081 ( .A(G2084), .B(G34), .Z(n986) );
  XNOR2_X1 U1082 ( .A(KEYINPUT54), .B(n986), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(n990), .B(n989), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(G29), .A2(n991), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(G11), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(n995), .B(KEYINPUT127), .ZN(n1024) );
  XOR2_X1 U1089 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1091 ( .A(KEYINPUT118), .B(n998), .Z(n999) );
  XNOR2_X1 U1092 ( .A(KEYINPUT51), .B(n999), .ZN(n1016) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1000), .Z(n1002) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(G160), .B(G2084), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(KEYINPUT117), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1019), .ZN(n1021) );
  INV_X1 U1107 ( .A(KEYINPUT55), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(G29), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

