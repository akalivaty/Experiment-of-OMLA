//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G50), .ZN(new_n205));
  INV_X1    g0005(.A(G226), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G116), .A2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n207), .B(new_n212), .C1(G107), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n219), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n227), .A2(G1), .A3(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G50), .B1(G58), .B2(G68), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n224), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n226), .A2(new_n228), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n214), .A2(KEYINPUT8), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT69), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT69), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n258), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n231), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n231), .A2(new_n265), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G58), .A2(G68), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n231), .B1(new_n268), .B2(new_n205), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n255), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n254), .B1(G1), .B2(new_n231), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G50), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n270), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G169), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT68), .A4(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G223), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n283), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G222), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n288), .B(new_n292), .C1(new_n293), .C2(new_n290), .ZN(new_n294));
  AND2_X1   g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n230), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT66), .B(G41), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n274), .B(G274), .C1(new_n298), .C2(G45), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n295), .A2(new_n225), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  XOR2_X1   g0104(.A(KEYINPUT67), .B(G226), .Z(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n297), .A2(new_n299), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n279), .B1(new_n280), .B2(new_n307), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n307), .A2(KEYINPUT70), .A3(G179), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT70), .B1(new_n307), .B2(G179), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n286), .A2(G238), .A3(new_n287), .ZN(new_n312));
  INV_X1    g0112(.A(G107), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n290), .A2(new_n291), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n312), .B1(new_n313), .B2(new_n290), .C1(new_n215), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n296), .ZN(new_n316));
  INV_X1    g0116(.A(G244), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n299), .C1(new_n317), .C2(new_n303), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G200), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n271), .A2(new_n293), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT72), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n275), .A2(G77), .ZN(new_n322));
  OR2_X1    g0122(.A1(KEYINPUT15), .A2(G87), .ZN(new_n323));
  NAND2_X1  g0123(.A1(KEYINPUT15), .A2(G87), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(KEYINPUT71), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(new_n263), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n256), .A2(new_n260), .ZN(new_n331));
  INV_X1    g0131(.A(new_n266), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(new_n332), .B1(G20), .B2(G77), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n254), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n321), .A2(new_n322), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n319), .B(new_n335), .C1(new_n336), .C2(new_n318), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n307), .A2(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT73), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT73), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n307), .A2(new_n340), .A3(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n278), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n270), .A2(KEYINPUT9), .A3(new_n273), .A4(new_n277), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n307), .A2(new_n336), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n342), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n349), .B1(new_n342), .B2(new_n348), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n311), .B(new_n337), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n282), .A2(new_n283), .A3(G232), .A4(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n314), .B2(new_n206), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n354), .B2(KEYINPUT74), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n296), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n299), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT75), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT75), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n304), .A2(G238), .B1(new_n299), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n359), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n359), .A2(new_n366), .A3(new_n361), .A4(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OR3_X1    g0168(.A1(new_n368), .A2(KEYINPUT76), .A3(new_n336), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n263), .A2(new_n293), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n266), .A2(new_n205), .B1(new_n231), .B2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n255), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  XOR2_X1   g0172(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n373));
  XNOR2_X1  g0173(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n275), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n216), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT12), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n216), .B2(new_n271), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n368), .B2(G200), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT76), .B1(new_n368), .B2(new_n336), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n369), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT78), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n368), .A2(G169), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n368), .A2(new_n387), .B1(new_n384), .B2(new_n385), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(new_n385), .ZN(new_n389));
  AOI211_X1 g0189(.A(new_n280), .B(new_n389), .C1(new_n365), .C2(new_n367), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n380), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n383), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n353), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n262), .A2(new_n275), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n272), .B2(new_n262), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n290), .A2(new_n399), .A3(G20), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n289), .B2(new_n231), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(G58), .B(G68), .ZN(new_n403));
  AOI22_X1  g0203(.A1(G20), .A2(new_n403), .B1(new_n332), .B2(G159), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT16), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n404), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n265), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT79), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n281), .B2(G33), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n407), .B1(new_n282), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT7), .B1(new_n410), .B2(G20), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n281), .A3(G33), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT79), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(new_n399), .A3(new_n231), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(G68), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n411), .A2(KEYINPUT80), .A3(G68), .A4(new_n416), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n406), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n405), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n398), .B1(new_n422), .B2(new_n255), .ZN(new_n423));
  INV_X1    g0223(.A(G41), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n229), .B1(new_n265), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n206), .A2(G1698), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n410), .B(new_n426), .C1(G223), .C2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G87), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n303), .A2(new_n215), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n429), .A2(new_n430), .A3(new_n360), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G179), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n280), .B2(new_n431), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n395), .B1(new_n423), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n415), .A2(new_n399), .A3(new_n231), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n399), .B1(new_n415), .B2(new_n231), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT80), .B1(new_n438), .B2(G68), .ZN(new_n439));
  INV_X1    g0239(.A(new_n420), .ZN(new_n440));
  OAI211_X1 g0240(.A(KEYINPUT16), .B(new_n404), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n405), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n255), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n397), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .A3(new_n433), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  INV_X1    g0247(.A(new_n429), .ZN(new_n448));
  INV_X1    g0248(.A(new_n430), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(new_n336), .A3(new_n449), .A4(new_n299), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n431), .B2(G200), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT17), .B1(new_n423), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n443), .A2(KEYINPUT17), .A3(new_n397), .A4(new_n451), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n447), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n443), .A2(new_n397), .A3(new_n451), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT17), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(KEYINPUT81), .A3(new_n453), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n446), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT82), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n335), .B1(new_n280), .B2(new_n318), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n318), .A2(G179), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n394), .A2(new_n460), .A3(new_n461), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n311), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n342), .A2(new_n348), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT10), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(new_n350), .ZN(new_n470));
  INV_X1    g0270(.A(new_n386), .ZN(new_n471));
  INV_X1    g0271(.A(new_n390), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n380), .B1(new_n473), .B2(new_n388), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n470), .A2(new_n474), .A3(new_n383), .A4(new_n337), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n435), .A2(new_n445), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n458), .A2(KEYINPUT81), .A3(new_n453), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT81), .B1(new_n458), .B2(new_n453), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n465), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT82), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n466), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n410), .A2(KEYINPUT22), .A3(new_n231), .A4(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G116), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G20), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT90), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n282), .A2(new_n283), .A3(new_n231), .A4(G87), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT23), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n231), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n313), .A2(KEYINPUT23), .A3(G20), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n486), .A2(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT24), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n482), .A2(KEYINPUT24), .A3(new_n485), .A4(new_n491), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n255), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n275), .A2(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n211), .A2(new_n291), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n410), .B(new_n500), .C1(G257), .C2(new_n291), .ZN(new_n501));
  XOR2_X1   g0301(.A(KEYINPUT91), .B(G294), .Z(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G33), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n425), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT5), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n274), .B(G45), .C1(new_n505), .C2(G41), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n298), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n300), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G264), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(G274), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  INV_X1    g0314(.A(new_n512), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n504), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G190), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT83), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n265), .A2(G1), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n254), .A2(new_n518), .A3(new_n275), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n226), .A2(new_n228), .A3(new_n275), .A4(new_n253), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT83), .B1(new_n522), .B2(new_n519), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G107), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n499), .A2(new_n514), .A3(new_n517), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n409), .A2(new_n282), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n291), .A3(new_n412), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n529), .B2(new_n317), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n527), .A2(new_n317), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(new_n291), .A3(new_n282), .A4(new_n283), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n282), .A2(new_n283), .A3(G250), .A4(G1698), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n425), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n298), .A2(new_n505), .ZN(new_n537));
  INV_X1    g0337(.A(new_n506), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n301), .ZN(new_n540));
  INV_X1    g0340(.A(G257), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n512), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G190), .ZN(new_n544));
  INV_X1    g0344(.A(G97), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n521), .B2(new_n523), .ZN(new_n546));
  OAI21_X1  g0346(.A(G107), .B1(new_n400), .B2(new_n401), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n332), .A2(G77), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n313), .A2(KEYINPUT6), .A3(G97), .ZN(new_n549));
  XOR2_X1   g0349(.A(G97), .B(G107), .Z(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n550), .B2(KEYINPUT6), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G20), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n546), .B1(new_n553), .B2(new_n255), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n275), .A2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n536), .B2(new_n542), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n544), .A2(new_n554), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT84), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n556), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n530), .A2(new_n535), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n296), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n515), .B1(G257), .B2(new_n508), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(G179), .ZN(new_n564));
  OAI21_X1  g0364(.A(G169), .B1(new_n536), .B2(new_n542), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n546), .B(new_n555), .C1(new_n553), .C2(new_n255), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n544), .A4(new_n557), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n526), .A2(new_n559), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n541), .A2(new_n291), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n410), .B(new_n573), .C1(G264), .C2(new_n291), .ZN(new_n574));
  INV_X1    g0374(.A(G303), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n290), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n296), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n539), .A2(G270), .A3(new_n301), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n578), .A2(KEYINPUT88), .A3(new_n512), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT88), .B1(new_n578), .B2(new_n512), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n533), .B(new_n231), .C1(G33), .C2(new_n545), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n255), .B(new_n582), .C1(new_n231), .C2(G116), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT89), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT20), .ZN(new_n585));
  INV_X1    g0385(.A(G116), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n254), .B1(G20), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(KEYINPUT20), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n584), .A2(KEYINPUT20), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n582), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n376), .A2(new_n586), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n226), .A2(new_n228), .A3(new_n275), .A4(new_n253), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(G116), .A3(new_n520), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n585), .A2(new_n590), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n581), .A2(G169), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n581), .A2(G200), .ZN(new_n598));
  INV_X1    g0398(.A(new_n594), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n577), .B(G190), .C1(new_n579), .C2(new_n580), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n581), .A2(new_n387), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n594), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n581), .A2(KEYINPUT21), .A3(new_n594), .A4(G169), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n597), .A2(new_n601), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n217), .A2(new_n291), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n317), .A2(G1698), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n483), .B1(new_n415), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n296), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n274), .A2(G45), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(G250), .C1(new_n295), .C2(new_n225), .ZN(new_n612));
  INV_X1    g0412(.A(G274), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT85), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n617), .B(new_n614), .C1(new_n609), .C2(new_n296), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n387), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n329), .A2(KEYINPUT86), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT86), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n327), .A2(new_n621), .A3(new_n328), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n620), .A2(new_n622), .B1(new_n521), .B2(new_n523), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT19), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n231), .B1(new_n357), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(G87), .B2(new_n203), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n625), .B1(new_n263), .B2(new_n545), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n231), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n216), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n630), .A2(new_n255), .B1(new_n329), .B2(new_n376), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n619), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n528), .A2(new_n412), .A3(new_n607), .A4(new_n606), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n425), .B1(new_n634), .B2(new_n483), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n617), .B1(new_n635), .B2(new_n614), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n610), .A2(KEYINPUT85), .A3(new_n615), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(G169), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n513), .A2(new_n280), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n496), .A2(new_n525), .A3(new_n498), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n516), .A2(new_n387), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(G190), .B1(new_n616), .B2(new_n618), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n518), .B1(new_n592), .B2(new_n520), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n522), .A2(KEYINPUT83), .A3(new_n519), .ZN(new_n647));
  OAI21_X1  g0447(.A(G87), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n524), .A2(KEYINPUT87), .A3(G87), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n636), .A2(new_n637), .A3(G200), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n645), .A2(new_n652), .A3(new_n631), .A4(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n640), .A2(new_n644), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n605), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n481), .A2(new_n572), .A3(new_n656), .ZN(G372));
  INV_X1    g0457(.A(KEYINPUT94), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n566), .A2(KEYINPUT93), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n564), .A2(new_n565), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n560), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT87), .B1(new_n524), .B2(G87), .ZN(new_n663));
  AOI211_X1 g0463(.A(new_n649), .B(new_n210), .C1(new_n521), .C2(new_n523), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n631), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n336), .B1(new_n636), .B2(new_n637), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n610), .A2(new_n615), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G200), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(G179), .B1(new_n636), .B2(new_n637), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n630), .A2(new_n255), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n329), .A2(new_n376), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n623), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n635), .A2(new_n614), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G169), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n671), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT92), .B1(new_n670), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n645), .A2(new_n652), .A3(new_n631), .A4(new_n668), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT92), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n667), .A2(new_n280), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n619), .A2(new_n632), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n662), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n658), .B1(new_n685), .B2(KEYINPUT26), .ZN(new_n686));
  INV_X1    g0486(.A(new_n567), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n654), .ZN(new_n688));
  INV_X1    g0488(.A(new_n661), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n660), .B1(new_n564), .B2(new_n565), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n689), .A2(new_n690), .A3(new_n568), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n681), .B1(new_n680), .B2(new_n683), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(KEYINPUT94), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n686), .A2(new_n688), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n597), .A2(new_n603), .A3(new_n604), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n698), .A2(new_n644), .B1(new_n684), .B2(new_n679), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n678), .B1(new_n699), .B2(new_n572), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n481), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n465), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n383), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n474), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n455), .A2(new_n459), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n476), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n351), .A2(new_n352), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n467), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n702), .A2(new_n711), .ZN(G369));
  INV_X1    g0512(.A(G13), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n715), .A2(KEYINPUT27), .A3(G1), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT27), .B1(new_n715), .B2(G1), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G213), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G343), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n594), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT95), .Z(new_n722));
  NAND3_X1  g0522(.A1(new_n597), .A2(new_n603), .A3(new_n604), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n605), .B2(new_n722), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  INV_X1    g0526(.A(new_n644), .ZN(new_n727));
  INV_X1    g0527(.A(new_n720), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n642), .A2(new_n720), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n526), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n729), .B1(new_n731), .B2(new_n727), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n731), .A2(new_n644), .A3(new_n723), .A4(new_n728), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n729), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n733), .A2(new_n735), .ZN(G399));
  INV_X1    g0536(.A(new_n222), .ZN(new_n737));
  OR3_X1    g0537(.A1(new_n737), .A2(new_n298), .A3(KEYINPUT96), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT96), .B1(new_n737), .B2(new_n298), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(G1), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n233), .B2(new_n740), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n602), .A2(new_n543), .A3(new_n511), .A4(new_n638), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n676), .A2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n513), .A2(new_n581), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n543), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(new_n746), .B2(new_n747), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n728), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n656), .A2(new_n572), .A3(new_n728), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(KEYINPUT31), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n752), .A2(KEYINPUT97), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n748), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n752), .A2(KEYINPUT97), .ZN(new_n759));
  OAI211_X1 g0559(.A(KEYINPUT31), .B(new_n720), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n745), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n723), .A2(new_n727), .B1(new_n692), .B2(new_n693), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n683), .B1(new_n763), .B2(new_n571), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n687), .A2(new_n640), .A3(new_n695), .A4(new_n654), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n685), .B2(new_n695), .ZN(new_n766));
  OAI211_X1 g0566(.A(KEYINPUT29), .B(new_n728), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n720), .B1(new_n697), .B2(new_n700), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n744), .B1(new_n773), .B2(G1), .ZN(G364));
  OR2_X1    g0574(.A1(new_n725), .A2(G330), .ZN(new_n775));
  INV_X1    g0575(.A(new_n740), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n274), .B1(new_n714), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n775), .A2(new_n726), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n231), .A2(new_n336), .ZN(new_n782));
  INV_X1    g0582(.A(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G179), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n575), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n782), .A2(G179), .A3(new_n783), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n231), .A2(G190), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(G179), .A3(new_n783), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n787), .A2(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G179), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n786), .B(new_n792), .C1(G329), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n387), .A2(new_n783), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT102), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n789), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(new_n797), .B2(new_n789), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n789), .A2(new_n784), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n803), .A2(new_n804), .B1(G283), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n231), .B1(new_n793), .B2(G190), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n502), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n796), .A2(new_n289), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n782), .A2(new_n797), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(G326), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n803), .A2(G68), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n808), .A2(new_n545), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n289), .B(new_n816), .C1(G50), .C2(new_n813), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n805), .A2(new_n313), .ZN(new_n818));
  INV_X1    g0618(.A(new_n787), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(G58), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n790), .ZN(new_n821));
  INV_X1    g0621(.A(new_n785), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n821), .A2(G77), .B1(new_n822), .B2(G87), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n815), .A2(new_n817), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT100), .B(G159), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n795), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT101), .B(KEYINPUT32), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n811), .A2(new_n814), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n230), .B1(G20), .B2(new_n280), .ZN(new_n830));
  INV_X1    g0630(.A(G45), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n234), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n410), .A2(new_n737), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n251), .C2(new_n831), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n290), .A2(G355), .A3(new_n222), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(G116), .C2(new_n222), .ZN(new_n836));
  NOR2_X1   g0636(.A1(G13), .A2(G33), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(G20), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n830), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT99), .Z(new_n841));
  AOI22_X1  g0641(.A1(new_n829), .A2(new_n830), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n839), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n725), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n781), .B1(new_n780), .B2(new_n844), .ZN(G396));
  NAND2_X1  g0645(.A1(new_n701), .A2(new_n728), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n335), .A2(new_n728), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n465), .A2(KEYINPUT103), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT103), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n462), .B2(new_n464), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n337), .B(new_n847), .C1(new_n848), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n703), .A2(new_n720), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT104), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n337), .B1(new_n848), .B2(new_n850), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(new_n761), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n780), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n837), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n289), .B1(new_n802), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G107), .B2(new_n822), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n812), .A2(new_n575), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n816), .B(new_n865), .C1(G294), .C2(new_n819), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n821), .A2(G116), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n805), .A2(new_n210), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G311), .B2(new_n795), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G143), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n787), .A2(new_n871), .B1(new_n812), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n825), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n790), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(new_n803), .C2(G150), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT34), .Z(new_n877));
  AOI22_X1  g0677(.A1(G50), .A2(new_n822), .B1(new_n806), .B2(G68), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n415), .B1(G132), .B2(new_n795), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n808), .A2(new_n214), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n830), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n830), .A2(new_n837), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n293), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n861), .A2(new_n779), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n860), .A2(new_n886), .ZN(G384));
  AND2_X1   g0687(.A1(new_n753), .A2(KEYINPUT31), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n755), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n481), .A2(G330), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n392), .A2(new_n728), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n393), .A2(new_n891), .B1(new_n474), .B2(new_n728), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n853), .C1(new_n755), .C2(new_n888), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(KEYINPUT109), .A2(KEYINPUT40), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n404), .B1(new_n439), .B2(new_n440), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT16), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT105), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n421), .A2(new_n900), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n255), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n397), .ZN(new_n905));
  INV_X1    g0705(.A(new_n718), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT106), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT106), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n908), .B(new_n718), .C1(new_n904), .C2(new_n397), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n706), .B2(new_n476), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n444), .B1(new_n433), .B2(new_n906), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n456), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n419), .A2(new_n420), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n900), .B1(new_n915), .B2(new_n404), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n406), .B(new_n901), .C1(new_n419), .C2(new_n420), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n398), .B1(new_n918), .B2(new_n255), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n908), .B1(new_n919), .B2(new_n718), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n905), .A2(KEYINPUT106), .A3(new_n906), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n905), .A2(new_n433), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n920), .A2(new_n456), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n914), .B1(new_n923), .B2(KEYINPUT37), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n897), .B1(new_n911), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n914), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n456), .B1(new_n919), .B2(new_n434), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n927), .A2(new_n907), .A3(new_n909), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT37), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n931));
  INV_X1    g0731(.A(new_n910), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT38), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n894), .A2(new_n896), .B1(new_n925), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n893), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n718), .B1(new_n443), .B2(new_n397), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT37), .B1(new_n938), .B2(KEYINPUT107), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n913), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT107), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n423), .B2(new_n718), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n942), .A2(KEYINPUT37), .B1(new_n912), .B2(new_n456), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n458), .A2(new_n453), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n938), .B1(new_n446), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n897), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n934), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n894), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n935), .A2(new_n937), .B1(new_n950), .B2(KEYINPUT40), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n890), .B1(new_n951), .B2(new_n745), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(KEYINPUT40), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n925), .A2(new_n934), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n954), .B(new_n937), .C1(new_n893), .C2(new_n895), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n481), .A3(new_n889), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT108), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n466), .A2(new_n480), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n960), .B2(new_n771), .ZN(new_n961));
  INV_X1    g0761(.A(new_n767), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n846), .B2(new_n769), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(KEYINPUT108), .A3(new_n481), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n711), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n958), .B(new_n966), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n720), .B(new_n857), .C1(new_n697), .C2(new_n700), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n848), .A2(new_n720), .A3(new_n850), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n892), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n971), .A2(new_n954), .B1(new_n446), .B2(new_n718), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT39), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n949), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n474), .A2(new_n720), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n925), .A2(new_n934), .A3(KEYINPUT39), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n972), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n967), .B(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n274), .B2(new_n714), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n586), .B1(new_n551), .B2(KEYINPUT35), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n232), .C1(KEYINPUT35), .C2(new_n551), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT36), .ZN(new_n983));
  OAI21_X1  g0783(.A(G77), .B1(new_n214), .B2(new_n216), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n984), .A2(new_n233), .B1(G50), .B2(new_n216), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(G1), .A3(new_n713), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n983), .A3(new_n986), .ZN(G367));
  NAND2_X1  g0787(.A1(new_n679), .A2(new_n684), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n665), .A2(new_n720), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT110), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n683), .A2(new_n989), .ZN(new_n991));
  MUX2_X1   g0791(.A(new_n990), .B(KEYINPUT110), .S(new_n991), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n839), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n410), .B1(new_n803), .B2(new_n502), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n785), .B2(new_n586), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n805), .A2(new_n545), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G283), .B2(new_n821), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT115), .B(G311), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n813), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n994), .A2(new_n996), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G317), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n794), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n822), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n575), .B2(new_n787), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n808), .A2(new_n313), .ZN(new_n1006));
  NOR4_X1   g0806(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n819), .A2(G150), .B1(new_n806), .B2(G77), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n872), .B2(new_n794), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n808), .A2(new_n216), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n289), .B(new_n1010), .C1(new_n803), .C2(new_n825), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n205), .B2(new_n790), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(G143), .C2(new_n813), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n822), .A2(G58), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1007), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT47), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n830), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n833), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n840), .B1(new_n222), .B2(new_n329), .C1(new_n244), .C2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n993), .A2(new_n1017), .A3(new_n779), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT114), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n691), .A2(new_n720), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n560), .A2(new_n720), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n559), .A2(new_n570), .A3(new_n567), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n734), .A2(new_n729), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT45), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n726), .A2(KEYINPUT112), .A3(new_n732), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1025), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1031));
  NAND3_X1  g0831(.A1(new_n735), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1025), .B1(new_n734), .B2(new_n729), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(new_n1031), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n732), .B1(new_n698), .B2(new_n720), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n734), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1037), .A2(G330), .A3(new_n725), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n726), .A3(new_n734), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n762), .A3(new_n771), .A4(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1034), .A2(new_n1032), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1029), .B1(new_n1042), .B2(new_n1028), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n772), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n740), .B(KEYINPUT41), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1021), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1047), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n773), .B1(new_n1051), .B2(new_n1045), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1049), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(KEYINPUT114), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n778), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1030), .A2(new_n734), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT42), .Z(new_n1057));
  NAND2_X1  g0857(.A1(new_n1025), .A2(new_n727), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n720), .B1(new_n1058), .B2(new_n567), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT43), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1057), .A2(new_n1059), .B1(new_n1060), .B2(new_n992), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n992), .A2(new_n1060), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n726), .A2(new_n732), .A3(new_n1030), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1063), .B(new_n1064), .Z(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1020), .B1(new_n1055), .B2(new_n1066), .ZN(G387));
  AOI22_X1  g0867(.A1(new_n803), .A2(new_n999), .B1(G317), .B2(new_n819), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n575), .B2(new_n790), .C1(new_n788), .C2(new_n812), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT48), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n822), .A2(new_n502), .B1(new_n809), .B2(G283), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT117), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1070), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n795), .A2(G326), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n410), .B1(G116), .B2(new_n806), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n802), .A2(new_n262), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n620), .A2(new_n622), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n809), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n205), .B2(new_n787), .C1(new_n264), .C2(new_n794), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n997), .B(new_n1083), .C1(G68), .C2(new_n821), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G159), .A2(new_n813), .B1(new_n822), .B2(G77), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n410), .A3(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1079), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT118), .Z(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n830), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n732), .A2(new_n839), .ZN(new_n1090));
  OR3_X1    g0890(.A1(new_n741), .A2(new_n737), .A3(new_n289), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n331), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1092), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G68), .B2(G77), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT50), .B1(new_n1092), .B2(G50), .ZN(new_n1095));
  AOI21_X1  g0895(.A(G45), .B1(new_n741), .B2(KEYINPUT116), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n741), .A2(KEYINPUT116), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n833), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n241), .A2(new_n831), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1091), .B1(G107), .B2(new_n222), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n780), .B1(new_n1101), .B2(new_n841), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1089), .A2(new_n1090), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n773), .A2(new_n1040), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1040), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n740), .B1(new_n772), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1103), .B(new_n1107), .C1(new_n777), .C2(new_n1105), .ZN(G393));
  NAND2_X1  g0908(.A1(new_n1042), .A2(new_n1028), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(new_n733), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1046), .A2(new_n1047), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1111), .A2(new_n776), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1030), .A2(new_n839), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n840), .B1(new_n545), .B2(new_n222), .C1(new_n248), .C2(new_n1018), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n410), .B1(new_n216), .B2(new_n785), .C1(new_n1092), .C2(new_n790), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G77), .B2(new_n809), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n803), .A2(G50), .ZN(new_n1117));
  INV_X1    g0917(.A(G159), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n787), .A2(new_n1118), .B1(new_n812), .B2(new_n264), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT51), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n868), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1116), .A2(new_n1117), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G143), .B2(new_n795), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n787), .A2(new_n791), .B1(new_n812), .B2(new_n1002), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT52), .Z(new_n1126));
  INV_X1    g0926(.A(G294), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n289), .B1(new_n1127), .B2(new_n790), .C1(new_n802), .C2(new_n575), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n818), .B1(G116), .B2(new_n809), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n862), .B2(new_n785), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n794), .A2(new_n788), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n830), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1113), .A2(new_n779), .A3(new_n1114), .A4(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1110), .B2(new_n777), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1112), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G390));
  AOI21_X1  g0937(.A(KEYINPUT38), .B1(new_n944), .B2(new_n946), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n1140), .B2(KEYINPUT38), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n976), .B1(new_n1141), .B2(KEYINPUT39), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n837), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n290), .B1(new_n803), .B2(G107), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n293), .B2(new_n808), .C1(new_n545), .C2(new_n790), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n812), .A2(new_n862), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n785), .A2(new_n210), .B1(new_n805), .B2(new_n216), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n787), .A2(new_n586), .B1(new_n794), .B2(new_n1127), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n803), .A2(G137), .B1(G125), .B2(new_n795), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n290), .C1(new_n1151), .C2(new_n812), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT54), .B(G143), .Z(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n790), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n822), .A2(G150), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n819), .A2(G132), .B1(new_n806), .B2(G50), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1118), .B2(new_n808), .ZN(new_n1159));
  NOR4_X1   g0959(.A1(new_n1152), .A2(new_n1155), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n830), .B1(new_n1149), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n884), .A2(new_n262), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1143), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n779), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n975), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n970), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n969), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n728), .B1(new_n764), .B2(new_n766), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n857), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n892), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n975), .B1(new_n934), .B2(new_n948), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1142), .A2(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n893), .A2(new_n745), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT119), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n761), .A2(new_n853), .A3(new_n892), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT119), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n974), .A2(new_n976), .B1(new_n970), .B2(new_n1165), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1171), .A2(new_n1170), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1173), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1164), .B1(new_n1182), .B2(new_n777), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n960), .A2(new_n771), .A3(new_n959), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT108), .B1(new_n963), .B2(new_n481), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n711), .B(new_n890), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT120), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n965), .A2(KEYINPUT120), .A3(new_n711), .A4(new_n890), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n892), .B1(new_n761), .B2(new_n853), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1190), .A2(new_n1173), .B1(new_n968), .B2(new_n969), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1169), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n889), .A2(G330), .A3(new_n853), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1176), .B(new_n1192), .C1(new_n1193), .C2(new_n892), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1188), .A2(new_n1189), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1182), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n740), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1182), .A2(new_n1196), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1183), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(G378));
  NAND2_X1  g1001(.A1(new_n278), .A2(new_n906), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n470), .B(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n837), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n410), .B(new_n298), .C1(new_n803), .C2(G97), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n293), .B2(new_n785), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1081), .B2(new_n821), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n787), .A2(new_n313), .B1(new_n812), .B2(new_n586), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1010), .B(new_n1210), .C1(G283), .C2(new_n795), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(new_n214), .C2(new_n805), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT121), .Z(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT58), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n205), .B1(G33), .B2(G41), .C1(new_n410), .C2(new_n298), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n803), .A2(G132), .B1(G125), .B2(new_n813), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n787), .A2(new_n1151), .B1(new_n790), .B2(new_n872), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G150), .B2(new_n809), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(new_n785), .C2(new_n1154), .ZN(new_n1219));
  XOR2_X1   g1019(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1220));
  XOR2_X1   g1020(.A(new_n1219), .B(new_n1220), .Z(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n805), .B2(new_n874), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1215), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n830), .B1(new_n1214), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n884), .A2(new_n205), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1206), .A2(new_n779), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1205), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n956), .B2(G330), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n745), .B(new_n1205), .C1(new_n953), .C2(new_n955), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n978), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1205), .B1(new_n951), .B2(new_n745), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n956), .A2(G330), .A3(new_n1229), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n977), .A4(new_n972), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1228), .B1(new_n1236), .B2(new_n778), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1195), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1239), .B1(new_n1182), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1236), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT57), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n740), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(KEYINPUT57), .A3(new_n1236), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1238), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(G375));
  AOI21_X1  g1047(.A(new_n1195), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n1053), .A3(new_n1196), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT123), .Z(new_n1251));
  OR2_X1    g1051(.A1(new_n892), .A2(new_n838), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n819), .A2(G137), .B1(new_n809), .B2(G50), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1151), .B2(new_n794), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G58), .B2(new_n806), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n813), .A2(G132), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n415), .B1(new_n803), .B2(new_n1153), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n821), .A2(G150), .B1(new_n822), .B2(G159), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1127), .A2(new_n812), .B1(new_n790), .B2(new_n313), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n803), .B2(G116), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT124), .Z(new_n1262));
  AOI22_X1  g1062(.A1(G97), .A2(new_n822), .B1(new_n806), .B2(G77), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n289), .A3(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1082), .B1(new_n862), .B2(new_n787), .C1(new_n575), .C2(new_n794), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1259), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n830), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n884), .A2(new_n216), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1252), .A2(new_n779), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1240), .B2(new_n777), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT125), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1251), .A2(new_n1271), .ZN(G381));
  OAI211_X1 g1072(.A(new_n1020), .B(new_n1136), .C1(new_n1055), .C2(new_n1066), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(G381), .A2(G396), .A3(G393), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1246), .A2(new_n1200), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1274), .A2(new_n860), .A3(new_n886), .A4(new_n1276), .ZN(G407));
  OAI211_X1 g1077(.A(G407), .B(G213), .C1(G343), .C2(new_n1275), .ZN(G409));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G343), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1241), .A2(new_n1053), .A3(new_n1236), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1282), .A2(new_n1237), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(new_n1200), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1246), .B2(new_n1200), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1196), .B1(new_n1248), .B2(KEYINPUT60), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT126), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n740), .B1(new_n1248), .B2(KEYINPUT60), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1289), .B(new_n1196), .C1(new_n1248), .C2(KEYINPUT60), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1271), .ZN(new_n1292));
  INV_X1    g1092(.A(G384), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1291), .A2(G384), .A3(new_n1271), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT62), .B1(new_n1285), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1281), .A2(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1291), .A2(G384), .A3(new_n1271), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G384), .B1(new_n1291), .B2(new_n1271), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1294), .A2(new_n1295), .A3(new_n1298), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1285), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1245), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT57), .B1(new_n1241), .B2(new_n1236), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1306), .A2(new_n1307), .A3(new_n740), .ZN(new_n1308));
  OAI21_X1  g1108(.A(G378), .B1(new_n1308), .B2(new_n1238), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1305), .A2(new_n1309), .A3(new_n1310), .A4(new_n1284), .ZN(new_n1311));
  AND4_X1   g1111(.A1(new_n1279), .A2(new_n1297), .A3(new_n1304), .A4(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(G393), .B(G396), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1054), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT114), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n777), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1065), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1136), .B1(new_n1318), .B2(new_n1020), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1273), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1314), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G387), .A2(G390), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1273), .A3(new_n1313), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1200), .B1(new_n1326), .B2(new_n1237), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1282), .A2(new_n1237), .ZN(new_n1328));
  OAI22_X1  g1128(.A1(G378), .A2(new_n1328), .B1(new_n1280), .B2(G343), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1304), .A2(KEYINPUT63), .B1(new_n1330), .B2(new_n1305), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1305), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1325), .A3(new_n1279), .ZN(new_n1333));
  OAI22_X1  g1133(.A1(new_n1312), .A2(new_n1325), .B1(new_n1331), .B2(new_n1333), .ZN(G405));
  NAND3_X1  g1134(.A1(new_n1324), .A2(new_n1275), .A3(new_n1309), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1321), .B(new_n1323), .C1(new_n1276), .C2(new_n1327), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1335), .A2(new_n1336), .A3(new_n1305), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1305), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


