//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(KEYINPUT64), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(G567), .B2(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT64), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n463), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(new_n465), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(KEYINPUT65), .A3(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n477), .A2(KEYINPUT66), .A3(new_n463), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT66), .B1(new_n477), .B2(new_n463), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n483), .B1(G124), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT67), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n463), .A2(KEYINPUT68), .A3(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT68), .B1(new_n463), .B2(G114), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n493), .A3(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT69), .A3(new_n491), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n507), .B1(new_n464), .B2(new_n465), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n507), .B(new_n510), .C1(new_n465), .C2(new_n464), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n503), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n503), .B2(new_n512), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(G164));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  OAI211_X1 g100(.A(G50), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n527), .A2(new_n528), .B1(new_n524), .B2(new_n525), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n533), .B(new_n526), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n523), .B1(new_n532), .B2(new_n534), .ZN(G166));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  OR2_X1    g112(.A1(KEYINPUT6), .A2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT6), .A2(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n528), .A2(new_n527), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(G89), .ZN(new_n545));
  NAND2_X1  g120(.A1(G63), .A2(G651), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n522), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n541), .A2(new_n551), .B1(new_n529), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  AOI22_X1  g129(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n522), .ZN(new_n556));
  INV_X1    g131(.A(new_n529), .ZN(new_n557));
  INV_X1    g132(.A(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n538), .B2(new_n539), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n557), .A2(G81), .B1(G43), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g139(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n518), .B2(new_n519), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g149(.A(KEYINPUT73), .B(new_n572), .C1(new_n544), .C2(new_n570), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(G651), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n559), .A2(new_n577), .A3(G53), .ZN(new_n578));
  OAI211_X1 g153(.A(G53), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n557), .A2(G91), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  OR2_X1    g159(.A1(new_n543), .A2(new_n547), .ZN(G286));
  XNOR2_X1  g160(.A(G166), .B(KEYINPUT74), .ZN(G303));
  NAND2_X1  g161(.A1(new_n557), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n559), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  INV_X1    g165(.A(G73), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT75), .B1(new_n591), .B2(new_n558), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n593), .A2(G73), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n592), .B(new_n594), .C1(new_n544), .C2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G48), .B2(new_n559), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n557), .A2(G86), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n522), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n541), .A2(new_n602), .B1(new_n529), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n557), .A2(G92), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT10), .Z(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n544), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n559), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n607), .B1(new_n615), .B2(G868), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT76), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(G868), .B2(new_n620), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(G868), .B2(new_n620), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n561), .A2(G868), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n614), .A2(G559), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT77), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(G868), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(new_n481), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G135), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT78), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n463), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n487), .A2(G123), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n479), .A2(new_n470), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT80), .Z(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT81), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n662), .A3(G14), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(KEYINPUT17), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n669), .B1(new_n671), .B2(new_n667), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT82), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  OR2_X1    g250(.A1(new_n666), .A2(new_n667), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n675), .C1(new_n671), .C2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  INV_X1    g262(.A(new_n682), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n684), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n687), .B(new_n691), .C1(new_n688), .C2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G229));
  XOR2_X1   g273(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT85), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G22), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G166), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n703), .B1(new_n704), .B2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n705), .A2(G23), .ZN(new_n715));
  INV_X1    g290(.A(G288), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n705), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT33), .B(G1976), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G1971), .B2(new_n711), .ZN(new_n720));
  OR3_X1    g295(.A1(new_n713), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n714), .B1(new_n713), .B2(new_n720), .ZN(new_n722));
  AOI21_X1  g297(.A(KEYINPUT34), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT84), .B(G29), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n487), .A2(G119), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n630), .A2(G131), .ZN(new_n727));
  OR2_X1    g302(.A1(G95), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n724), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n605), .A2(new_n708), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G24), .B2(new_n708), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G1986), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(G1986), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n723), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n721), .A2(KEYINPUT34), .A3(new_n722), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n700), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n724), .ZN(new_n743));
  NAND2_X1  g318(.A1(G162), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G35), .B2(new_n743), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(G2090), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n562), .A2(new_n709), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G19), .B2(new_n709), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT88), .B(G1341), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT90), .B(G28), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n754), .B(new_n755), .C1(new_n757), .C2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G34), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n724), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G160), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n759), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n752), .A2(new_n753), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT25), .Z(new_n772));
  AOI22_X1  g347(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  INV_X1    g348(.A(G139), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n772), .B1(new_n463), .B2(new_n773), .C1(new_n481), .C2(new_n774), .ZN(new_n775));
  MUX2_X1   g350(.A(G33), .B(new_n775), .S(G29), .Z(new_n776));
  AOI22_X1  g351(.A1(new_n637), .A2(new_n743), .B1(G2072), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT26), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n780), .A2(new_n781), .B1(G105), .B2(new_n470), .ZN(new_n782));
  INV_X1    g357(.A(G141), .ZN(new_n783));
  INV_X1    g358(.A(G129), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n782), .B1(new_n481), .B2(new_n783), .C1(new_n486), .C2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G32), .B(new_n785), .S(G29), .Z(new_n786));
  XOR2_X1   g361(.A(KEYINPUT27), .B(G1996), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G5), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G171), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1961), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n762), .B2(new_n768), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n770), .A2(new_n777), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n630), .A2(G140), .ZN(new_n794));
  INV_X1    g369(.A(G128), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n463), .A2(G116), .ZN(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n794), .B1(new_n795), .B2(new_n486), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n724), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT28), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G2067), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n705), .A2(G4), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n615), .B2(new_n705), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(G1348), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n776), .A2(G2072), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(G1348), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n804), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n793), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n746), .A2(new_n747), .ZN(new_n812));
  INV_X1    g387(.A(G2090), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n743), .A2(G27), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G164), .B2(new_n743), .ZN(new_n816));
  INV_X1    g391(.A(G2078), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n705), .A2(G21), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G168), .B2(new_n705), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT89), .ZN(new_n821));
  INV_X1    g396(.A(G1966), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n709), .A2(G20), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT23), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n620), .B2(new_n705), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT92), .B(G1956), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n821), .A2(new_n822), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n786), .A2(new_n787), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n823), .A2(new_n828), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n811), .A2(new_n814), .A3(new_n818), .A4(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n742), .A2(new_n750), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n740), .A2(KEYINPUT87), .A3(KEYINPUT36), .A4(new_n741), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(G311));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n833), .B2(new_n834), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n750), .A2(new_n832), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n740), .A2(new_n741), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n699), .ZN(new_n840));
  AND4_X1   g415(.A1(new_n836), .A2(new_n838), .A3(new_n840), .A4(new_n834), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(G150));
  AOI22_X1  g417(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(new_n522), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT94), .B(G55), .Z(new_n845));
  XOR2_X1   g420(.A(KEYINPUT95), .B(G93), .Z(new_n846));
  OAI22_X1  g421(.A1(new_n541), .A2(new_n845), .B1(new_n529), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n561), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n562), .A2(KEYINPUT96), .A3(new_n848), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n615), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT97), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n849), .B1(new_n859), .B2(new_n860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n851), .B1(new_n862), .B2(new_n863), .ZN(G145));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n866));
  INV_X1    g441(.A(G118), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n865), .A2(new_n866), .B1(new_n867), .B2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n866), .B2(new_n865), .ZN(new_n869));
  INV_X1    g444(.A(G130), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n486), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(G142), .B2(new_n630), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n642), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n785), .B(new_n775), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n503), .A2(new_n512), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n798), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n730), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n875), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G162), .B(new_n767), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n637), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n881), .B2(new_n879), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n615), .A2(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n614), .A2(new_n620), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n614), .A2(KEYINPUT99), .A3(new_n620), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n885), .A2(new_n886), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n627), .B(new_n856), .ZN(new_n894));
  MUX2_X1   g469(.A(new_n889), .B(new_n893), .S(new_n894), .Z(new_n895));
  XNOR2_X1  g470(.A(G290), .B(G305), .ZN(new_n896));
  NAND2_X1  g471(.A1(G166), .A2(G288), .ZN(new_n897));
  OR2_X1    g472(.A1(G166), .A2(G288), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n897), .ZN(new_n900));
  XNOR2_X1  g475(.A(G305), .B(new_n605), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT100), .B1(new_n899), .B2(new_n902), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n907), .A2(KEYINPUT42), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT101), .B1(new_n903), .B2(KEYINPUT42), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n895), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n895), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g491(.A(new_n915), .B1(G868), .B2(new_n848), .ZN(G331));
  XNOR2_X1  g492(.A(G286), .B(G171), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n856), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n854), .A2(new_n918), .A3(new_n855), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n889), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n921), .A2(KEYINPUT103), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(KEYINPUT103), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n856), .A2(KEYINPUT102), .A3(new_n919), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT102), .B1(new_n856), .B2(new_n919), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n924), .B(new_n925), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n907), .B(new_n923), .C1(new_n929), .C2(new_n893), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n923), .B1(new_n929), .B2(new_n893), .ZN(new_n933));
  INV_X1    g508(.A(new_n907), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n928), .B(new_n892), .C1(new_n891), .C2(new_n889), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(KEYINPUT104), .A3(new_n907), .A4(new_n923), .ZN(new_n937));
  INV_X1    g512(.A(G37), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n932), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n930), .B2(new_n931), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n922), .B1(new_n890), .B2(new_n891), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n889), .B1(new_n928), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n891), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n934), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n942), .A2(new_n943), .A3(new_n937), .A4(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n940), .A2(new_n941), .A3(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n932), .A2(new_n938), .A3(new_n937), .A4(new_n947), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT43), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n949), .B1(new_n956), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT74), .ZN(new_n959));
  OR2_X1    g534(.A1(G166), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(G166), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(G8), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(G303), .A2(KEYINPUT108), .A3(KEYINPUT55), .A4(G8), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n963), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT107), .B(G40), .Z(new_n969));
  NOR3_X1   g544(.A1(new_n468), .A2(new_n472), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n503), .B2(new_n512), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT69), .B1(new_n501), .B2(new_n491), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n497), .B(new_n490), .C1(new_n499), .C2(new_n500), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n511), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n510), .B1(new_n479), .B2(new_n507), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n504), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT70), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n514), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n973), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n704), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n971), .B1(new_n972), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n813), .B(new_n985), .C1(new_n981), .C2(new_n984), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n968), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n967), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n970), .B1(new_n972), .B2(new_n984), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n984), .B2(new_n981), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n813), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n968), .B1(new_n991), .B2(new_n983), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n967), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n716), .A2(G1976), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n970), .B(new_n998), .C1(new_n976), .C2(new_n979), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n999), .A2(new_n1000), .A3(G8), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n999), .B2(G8), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n995), .B(new_n997), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n999), .A2(G8), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT109), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n999), .A2(new_n1000), .A3(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(KEYINPUT111), .A3(new_n995), .A4(new_n997), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n597), .A2(new_n1012), .A3(new_n598), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT112), .B(G86), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n557), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n597), .B2(new_n1017), .ZN(new_n1018));
  OR3_X1    g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n1009), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1011), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1024), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT110), .B1(new_n1024), .B2(KEYINPUT52), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n994), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1005), .A2(new_n1010), .B1(new_n1009), .B2(new_n1021), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1007), .A2(new_n1008), .B1(G1976), .B2(new_n716), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1029), .A2(new_n1035), .A3(KEYINPUT114), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n993), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n762), .B(new_n985), .C1(new_n981), .C2(new_n984), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n970), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(KEYINPUT45), .B2(new_n981), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1038), .B(G168), .C1(new_n1040), .C2(G1966), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT126), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1040), .B2(G1966), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  OAI211_X1 g620(.A(G8), .B(new_n1041), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1038), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT45), .B(new_n998), .C1(new_n515), .C2(new_n516), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n876), .A2(new_n998), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n971), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1966), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(G8), .B(G286), .C1(new_n1047), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT125), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1043), .A2(KEYINPUT125), .A3(G8), .A4(G286), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1041), .A2(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n822), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n968), .B1(new_n1060), .B2(new_n1038), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1058), .B(KEYINPUT51), .C1(new_n1061), .C2(new_n1042), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1046), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT62), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1046), .A2(new_n1057), .A3(new_n1065), .A4(new_n1062), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n982), .A2(G2078), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  INV_X1    g643(.A(G1961), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n985), .B1(new_n981), .B2(new_n984), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1067), .A2(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n817), .ZN(new_n1072));
  AOI21_X1  g647(.A(G301), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1064), .A2(new_n1066), .A3(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n973), .B(new_n1075), .C1(new_n981), .C2(KEYINPUT45), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT118), .B(G1956), .Z(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n990), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n581), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT119), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n576), .A2(new_n582), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n576), .A2(KEYINPUT120), .A3(new_n582), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT121), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1088), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT120), .B1(new_n576), .B2(new_n582), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1093), .B(new_n1090), .C1(new_n1096), .C2(new_n1084), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1092), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1079), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1079), .A2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT50), .B(G1384), .C1(new_n980), .C2(new_n514), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1077), .B1(new_n1102), .B2(new_n989), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(KEYINPUT123), .A3(new_n1076), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1098), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1348), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1070), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n999), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n972), .A2(KEYINPUT122), .A3(new_n970), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n803), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n615), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1099), .B1(new_n1105), .B2(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  NAND3_X1  g691(.A1(new_n1109), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G1996), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(new_n973), .C1(new_n981), .C2(KEYINPUT45), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1109), .A2(new_n1110), .A3(KEYINPUT124), .A4(new_n1116), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(KEYINPUT59), .A3(new_n562), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1112), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n615), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT60), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT59), .B1(new_n1123), .B2(new_n562), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n1099), .A2(new_n1131), .B1(new_n615), .B2(new_n1125), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1079), .A2(new_n1098), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1103), .A2(new_n1092), .A3(new_n1097), .A4(new_n1076), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT61), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1115), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1138));
  XNOR2_X1  g713(.A(G171), .B(KEYINPUT54), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT106), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT45), .B1(new_n1049), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1141), .B2(new_n1049), .ZN(new_n1143));
  NAND4_X1  g718(.A1(G160), .A2(KEYINPUT53), .A3(G40), .A4(new_n817), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(KEYINPUT127), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT127), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1147), .A2(new_n1140), .A3(new_n1148), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1138), .A2(new_n1140), .B1(new_n1149), .B2(new_n1071), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1063), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1137), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1037), .B1(new_n1074), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1061), .A2(G168), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G288), .A2(G1976), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1014), .B1(new_n1022), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT113), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1009), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n988), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1155), .B1(new_n1037), .B2(new_n1154), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1029), .A2(new_n1035), .A3(KEYINPUT63), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT116), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n987), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n987), .A2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n967), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1166), .B(new_n1167), .C1(new_n1168), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n988), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n992), .A2(new_n967), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1029), .A2(new_n1035), .A3(KEYINPUT114), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT114), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1178), .B(new_n1154), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1174), .B1(new_n1181), .B2(new_n1156), .ZN(new_n1182));
  OAI221_X1 g757(.A(new_n1157), .B1(new_n1164), .B2(new_n988), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT117), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1153), .A2(new_n1175), .A3(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n798), .B(new_n803), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n785), .B(new_n1120), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n730), .B(new_n733), .Z(new_n1189));
  NOR2_X1   g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n605), .B(G1986), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1143), .A2(new_n971), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1185), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1193), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1196), .A2(G1986), .A3(G290), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT48), .ZN(new_n1198));
  OAI22_X1  g773(.A1(new_n1197), .A2(new_n1198), .B1(new_n1196), .B2(new_n1190), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1199), .B1(new_n1198), .B2(new_n1197), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1186), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1193), .B1(new_n1201), .B2(new_n785), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1193), .A2(new_n1120), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1203), .A2(KEYINPUT46), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1203), .A2(KEYINPUT46), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1202), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT47), .Z(new_n1207));
  NAND2_X1  g782(.A1(new_n731), .A2(new_n733), .ZN(new_n1208));
  OAI22_X1  g783(.A1(new_n1188), .A2(new_n1208), .B1(G2067), .B2(new_n798), .ZN(new_n1209));
  AOI211_X1 g784(.A(new_n1200), .B(new_n1207), .C1(new_n1193), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1195), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g786(.A1(new_n940), .A2(new_n948), .ZN(new_n1213));
  NOR3_X1   g787(.A1(G229), .A2(new_n461), .A3(G227), .ZN(new_n1214));
  NAND4_X1  g788(.A1(new_n1213), .A2(new_n883), .A3(new_n663), .A4(new_n1214), .ZN(G225));
  INV_X1    g789(.A(G225), .ZN(G308));
endmodule


