//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(G101), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n193), .A2(new_n194), .A3(KEYINPUT75), .A4(G101), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT0), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n205), .B2(new_n206), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n193), .A2(G101), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n188), .A2(new_n191), .A3(new_n214), .A4(new_n192), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n199), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n190), .A2(G104), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n187), .A2(G107), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n224), .A2(new_n201), .A3(new_n203), .ZN(new_n225));
  AOI21_X1  g039(.A(G128), .B1(new_n201), .B2(new_n203), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n202), .A2(KEYINPUT1), .A3(G146), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT10), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT76), .B1(new_n229), .B2(new_n221), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n215), .A2(new_n220), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT76), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n201), .A3(new_n203), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n237), .B(new_n227), .C1(G128), .C2(new_n210), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n233), .B1(new_n240), .B2(new_n230), .ZN(new_n241));
  AOI211_X1 g055(.A(KEYINPUT77), .B(KEYINPUT10), .C1(new_n234), .C2(new_n239), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n217), .B(new_n232), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT79), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR3_X1   g059(.A1(new_n229), .A2(KEYINPUT76), .A3(new_n221), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n236), .B1(new_n235), .B2(new_n238), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n230), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT77), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n240), .A2(new_n233), .A3(new_n230), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n251), .A2(KEYINPUT79), .A3(new_n217), .A4(new_n232), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n255), .A2(new_n258), .A3(new_n261), .A4(new_n256), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n245), .A2(new_n252), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G110), .B(G140), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(G227), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n265), .B(new_n267), .Z(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n217), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n223), .A2(new_n231), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n270), .B(new_n271), .C1(new_n249), .C2(new_n250), .ZN(new_n272));
  INV_X1    g086(.A(new_n263), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n234), .A2(new_n239), .B1(new_n221), .B2(new_n229), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT12), .ZN(new_n276));
  OR3_X1    g090(.A1(new_n275), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n275), .B2(new_n273), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n243), .B2(new_n263), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n264), .A2(new_n274), .B1(new_n280), .B2(new_n269), .ZN(new_n281));
  OAI21_X1  g095(.A(G469), .B1(new_n281), .B2(G902), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n272), .A2(new_n273), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n268), .B1(new_n264), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n279), .A3(new_n268), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n283), .B(new_n286), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n284), .A2(new_n285), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n282), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G221), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT9), .B(G234), .Z(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n283), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G116), .B(G119), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT2), .B(G113), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n302), .B(new_n303), .Z(new_n304));
  NAND3_X1  g118(.A1(new_n199), .A2(new_n304), .A3(new_n216), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT81), .ZN(new_n306));
  INV_X1    g120(.A(new_n302), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n303), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n309));
  INV_X1    g123(.A(G116), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(new_n310), .A3(G119), .ZN(new_n311));
  INV_X1    g125(.A(G113), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n302), .A2(new_n309), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n223), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n199), .A2(new_n317), .A3(new_n304), .A4(new_n216), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n306), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G122), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n306), .A2(new_n320), .A3(new_n316), .A4(new_n318), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT6), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n325), .A3(new_n321), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n209), .A2(new_n211), .A3(G125), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n327), .A2(KEYINPUT83), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(KEYINPUT83), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n229), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G224), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G953), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n334), .B(KEYINPUT84), .Z(new_n335));
  XNOR2_X1  g149(.A(new_n332), .B(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n324), .A2(new_n326), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT7), .B1(new_n333), .B2(G953), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n328), .A2(new_n339), .A3(new_n329), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n332), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n315), .A2(new_n221), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n320), .B(KEYINPUT8), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n302), .A2(KEYINPUT5), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n308), .B1(new_n313), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n342), .B(new_n343), .C1(new_n221), .C2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n341), .B1(KEYINPUT85), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n332), .A2(new_n340), .A3(new_n338), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n346), .A2(KEYINPUT85), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n323), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(new_n283), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G210), .B1(G237), .B2(G902), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n337), .A2(new_n283), .A3(new_n350), .A4(new_n352), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n301), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT87), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n356), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(KEYINPUT87), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n299), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n266), .A3(G214), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G143), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n202), .A2(KEYINPUT88), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G237), .A2(G953), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n368), .A2(KEYINPUT88), .A3(new_n202), .A4(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n261), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT17), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n367), .A2(G131), .A3(new_n369), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G125), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT69), .B1(new_n376), .B2(KEYINPUT16), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT69), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT16), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n375), .A4(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n330), .A2(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n377), .B(new_n380), .C1(new_n382), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n200), .ZN(new_n384));
  XNOR2_X1  g198(.A(G125), .B(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT16), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(G146), .A3(new_n377), .A4(new_n380), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n367), .A2(KEYINPUT17), .A3(G131), .A4(new_n369), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n374), .A2(new_n384), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G113), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n187), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT18), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n370), .B1(new_n392), .B2(new_n261), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n382), .A2(G146), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n385), .A2(new_n200), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n393), .B(new_n396), .C1(new_n392), .C2(new_n373), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n389), .A2(KEYINPUT90), .A3(new_n391), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n371), .A2(new_n373), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT89), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n371), .A2(new_n405), .A3(new_n373), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n387), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n385), .B(KEYINPUT19), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n408), .A2(new_n200), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n397), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n391), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G475), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n283), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT20), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n413), .A2(new_n417), .A3(new_n414), .A4(new_n283), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(KEYINPUT91), .A3(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n418), .A2(KEYINPUT91), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n391), .B1(new_n389), .B2(new_n397), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n400), .B2(new_n401), .ZN(new_n422));
  OAI21_X1  g236(.A(G475), .B1(new_n422), .B2(G902), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n266), .A2(G952), .ZN(new_n425));
  NAND2_X1  g239(.A1(G234), .A2(G237), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT21), .B(G898), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(G902), .A3(G953), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G116), .B(G122), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n190), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n434), .A2(new_n190), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT92), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT13), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n206), .B2(G143), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n206), .A2(G143), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n202), .A2(G128), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT93), .A3(new_n439), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n444), .A2(new_n439), .ZN(new_n447));
  OAI21_X1  g261(.A(G134), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n444), .A2(new_n443), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n254), .ZN(new_n450));
  INV_X1    g264(.A(new_n434), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G107), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n435), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n438), .A2(new_n448), .A3(new_n450), .A4(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n449), .B(new_n254), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n310), .A2(KEYINPUT14), .A3(G122), .ZN(new_n457));
  OAI211_X1 g271(.A(G107), .B(new_n457), .C1(new_n451), .C2(KEYINPUT14), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n435), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n295), .A2(G217), .A3(new_n266), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(KEYINPUT94), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n466), .A3(new_n461), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n283), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G478), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n468), .B(new_n474), .Z(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n424), .A2(new_n433), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT96), .B1(new_n361), .B2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n360), .A2(new_n358), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT96), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n477), .A4(new_n299), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT23), .B1(new_n206), .B2(G119), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT67), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n206), .A2(G119), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT67), .B(KEYINPUT23), .C1(new_n206), .C2(G119), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G119), .B(G128), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT24), .B(G110), .Z(new_n494));
  OAI22_X1  g308(.A1(new_n492), .A2(G110), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n395), .A3(new_n387), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n492), .B2(G110), .ZN(new_n499));
  INV_X1    g313(.A(G110), .ZN(new_n500));
  AOI211_X1 g314(.A(KEYINPUT68), .B(new_n500), .C1(new_n485), .C2(new_n491), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n384), .A2(new_n387), .B1(new_n493), .B2(new_n494), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n492), .A2(G110), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n492), .A2(new_n498), .A3(G110), .ZN(new_n507));
  AND4_X1   g321(.A1(new_n497), .A2(new_n506), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n496), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT22), .B(G137), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n496), .B(new_n512), .C1(new_n504), .C2(new_n508), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n283), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n514), .A2(KEYINPUT71), .A3(new_n283), .A4(new_n515), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT72), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n516), .A2(new_n519), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT72), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n518), .A2(new_n524), .A3(new_n519), .A4(new_n520), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G217), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(G234), .B2(new_n283), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n514), .A2(new_n515), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT73), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n528), .A2(G902), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n263), .A2(new_n212), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT64), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n254), .B2(G137), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n257), .A2(KEYINPUT64), .A3(G134), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n256), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G131), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n238), .A2(new_n262), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT30), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n541), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n535), .A2(KEYINPUT65), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n263), .A2(new_n547), .A3(new_n212), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n545), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n304), .ZN(new_n552));
  INV_X1    g366(.A(new_n304), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n368), .A2(G210), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(new_n214), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n556), .B(new_n557), .Z(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n554), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n304), .B2(new_n551), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(KEYINPUT31), .A3(new_n558), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n542), .A2(new_n304), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n542), .B2(new_n304), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n565), .B(new_n567), .C1(new_n554), .C2(new_n566), .ZN(new_n568));
  INV_X1    g382(.A(new_n558), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n561), .A2(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(G472), .A2(G902), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(KEYINPUT32), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT32), .ZN(new_n574));
  INV_X1    g388(.A(new_n572), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n549), .B(new_n553), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT28), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n567), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n558), .A2(KEYINPUT29), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n283), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n563), .A2(new_n569), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n558), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT29), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(G472), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n573), .A2(new_n576), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n534), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n479), .A2(new_n482), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT97), .B(G101), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G3));
  NOR2_X1   g405(.A1(new_n570), .A2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(KEYINPUT98), .A2(G472), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n534), .A2(new_n298), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n462), .A2(KEYINPUT33), .A3(new_n464), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n465), .A2(new_n597), .A3(new_n467), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n596), .B1(new_n598), .B2(KEYINPUT99), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n596), .A2(KEYINPUT99), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n469), .A2(G902), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n468), .A2(new_n469), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n424), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n359), .A2(new_n605), .A3(new_n433), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n595), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  NAND2_X1  g423(.A1(new_n416), .A2(new_n418), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n423), .ZN(new_n611));
  NOR4_X1   g425(.A1(new_n359), .A2(new_n433), .A3(new_n475), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n595), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT35), .B(G107), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  INV_X1    g429(.A(new_n594), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n513), .A2(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n509), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n532), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n529), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n619), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n526), .B2(new_n528), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT100), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n479), .A2(new_n482), .A3(new_n616), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G12));
  OR3_X1    g443(.A1(new_n431), .A2(KEYINPUT101), .A3(G900), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT101), .B1(new_n431), .B2(G900), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n427), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n611), .A2(new_n475), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n634), .A2(KEYINPUT102), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n299), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n626), .A2(new_n637), .A3(new_n356), .A4(new_n586), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  XNOR2_X1  g453(.A(new_n632), .B(KEYINPUT39), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n299), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n299), .A2(KEYINPUT40), .A3(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n354), .A2(new_n355), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT38), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n563), .A2(new_n569), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n283), .B1(new_n577), .B2(new_n558), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n573), .A2(new_n576), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n424), .A2(new_n476), .A3(new_n300), .ZN(new_n653));
  OR3_X1    g467(.A1(new_n620), .A2(KEYINPUT103), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n620), .B2(new_n653), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n645), .A2(new_n652), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G143), .ZN(G45));
  AOI21_X1  g471(.A(new_n587), .B1(new_n622), .B2(new_n625), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n424), .A2(new_n604), .A3(new_n632), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n658), .A2(new_n356), .A3(new_n299), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  AOI22_X1  g476(.A1(new_n526), .A2(new_n528), .B1(new_n532), .B2(new_n531), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n288), .A2(new_n290), .ZN(new_n664));
  INV_X1    g478(.A(new_n292), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(new_n283), .A3(new_n665), .A4(new_n286), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n283), .B1(new_n288), .B2(new_n290), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n297), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n663), .A2(new_n670), .A3(new_n586), .A4(new_n606), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT41), .B(G113), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NOR3_X1   g487(.A1(new_n534), .A2(new_n587), .A3(new_n669), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n612), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G116), .ZN(G18));
  NAND4_X1  g490(.A1(new_n658), .A2(new_n477), .A3(new_n356), .A4(new_n670), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  NAND4_X1  g492(.A1(new_n424), .A2(new_n646), .A3(new_n476), .A4(new_n300), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n561), .A2(new_n564), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n579), .A2(new_n569), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n575), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n571), .A2(new_n283), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(G472), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n529), .A2(new_n533), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n663), .A2(KEYINPUT104), .A3(new_n684), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n679), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n669), .A2(new_n433), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  INV_X1    g506(.A(G472), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n680), .A2(new_n681), .ZN(new_n694));
  OAI22_X1  g508(.A1(new_n592), .A2(new_n693), .B1(new_n694), .B2(new_n575), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n624), .A2(new_n659), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n356), .A3(new_n670), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  NOR3_X1   g512(.A1(new_n285), .A2(KEYINPUT105), .A3(G902), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n282), .A2(KEYINPUT105), .B1(new_n281), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n291), .A2(new_n292), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n297), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n281), .A2(new_n699), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n264), .A2(new_n274), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n280), .A2(new_n269), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n285), .B1(new_n708), .B2(new_n283), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n705), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n666), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT106), .A3(new_n297), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n704), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n646), .A2(new_n301), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n533), .A2(new_n529), .A3(new_n586), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n660), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n659), .B1(new_n704), .B2(new_n713), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n716), .A3(new_n720), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  NAND4_X1  g541(.A1(new_n714), .A2(new_n636), .A3(new_n635), .A4(new_n716), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n708), .B(KEYINPUT45), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT108), .A3(G469), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n281), .A2(KEYINPUT45), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n281), .A2(KEYINPUT45), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(G469), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n732), .A2(new_n737), .B1(G469), .B2(G902), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n730), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g553(.A1(G469), .A2(G902), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT108), .B1(new_n731), .B2(G469), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n735), .A2(new_n736), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(KEYINPUT109), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n738), .A2(KEYINPUT46), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n739), .A2(new_n745), .A3(new_n666), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n604), .A2(new_n420), .A3(new_n419), .A4(new_n423), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n620), .A3(new_n594), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n747), .A2(new_n297), .A3(new_n640), .A4(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n750), .A2(new_n620), .A3(KEYINPUT44), .A4(new_n594), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n755), .A2(new_n756), .A3(new_n715), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n755), .B2(new_n715), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n257), .ZN(G39));
  INV_X1    g575(.A(new_n715), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n663), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n586), .A2(new_n659), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n747), .A2(new_n297), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n763), .B(new_n764), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  AND3_X1   g585(.A1(new_n573), .A2(new_n576), .A3(new_n650), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n297), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n773), .A2(new_n647), .A3(new_n301), .A4(new_n748), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n666), .A2(new_n668), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT49), .Z(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n776), .A3(new_n663), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n476), .A2(new_n424), .A3(new_n646), .A4(new_n300), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n712), .A2(new_n781), .A3(new_n297), .A4(new_n651), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n624), .A2(new_n632), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n772), .A2(new_n679), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n623), .B(new_n633), .C1(new_n526), .C2(new_n528), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n296), .B1(new_n711), .B2(new_n666), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n785), .A2(new_n786), .A3(KEYINPUT112), .A4(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n661), .A2(new_n789), .A3(new_n638), .A4(new_n697), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n696), .A2(new_n356), .A3(new_n670), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n624), .A2(KEYINPUT100), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n621), .B(new_n623), .C1(new_n526), .C2(new_n528), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n356), .B(new_n586), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n793), .B1(new_n797), .B2(new_n637), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT52), .A3(new_n661), .A4(new_n789), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n792), .A2(KEYINPUT113), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n661), .A2(new_n638), .A3(new_n697), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT52), .A4(new_n789), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n433), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n424), .A2(new_n475), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n805), .B(new_n806), .C1(new_n360), .C2(new_n358), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n595), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n605), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n595), .A2(new_n805), .A3(new_n480), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n627), .A2(new_n811), .A3(new_n589), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n724), .A2(new_n716), .A3(new_n720), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n724), .A2(new_n716), .B1(new_n721), .B2(new_n720), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n728), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n611), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n298), .A2(new_n476), .A3(new_n633), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n658), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n714), .A2(new_n696), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n762), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n675), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n796), .A2(new_n669), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n825), .B1(new_n826), .B2(new_n477), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n671), .B1(new_n689), .B2(new_n690), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT114), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(KEYINPUT114), .A2(new_n828), .A3(new_n675), .A4(new_n677), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n815), .B(new_n824), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT53), .B1(new_n804), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n820), .B(new_n586), .C1(new_n794), .C2(new_n795), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n822), .B1(new_n833), .B2(new_n611), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n715), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n726), .A3(new_n728), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n828), .A2(new_n675), .A3(new_n677), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n836), .A2(new_n814), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n792), .A2(new_n799), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n838), .A2(new_n839), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n800), .A2(new_n803), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n840), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n843), .A2(new_n844), .B1(new_n845), .B2(KEYINPUT53), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n779), .A2(new_n842), .B1(new_n846), .B2(KEYINPUT54), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT116), .B1(new_n768), .B2(new_n769), .ZN(new_n849));
  INV_X1    g663(.A(new_n769), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n767), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n666), .A2(new_n296), .A3(new_n668), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n427), .B1(new_n687), .B2(new_n688), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n750), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n762), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n669), .A2(new_n427), .A3(new_n762), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n663), .A3(new_n772), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n424), .A3(new_n604), .ZN(new_n861));
  INV_X1    g675(.A(new_n856), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n647), .A2(new_n669), .A3(new_n300), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT117), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n862), .A2(KEYINPUT50), .A3(new_n864), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n859), .A2(new_n750), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n620), .A3(new_n684), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n848), .B1(new_n858), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n862), .A2(new_n356), .A3(new_n670), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n875), .B(new_n425), .C1(new_n605), .C2(new_n860), .ZN(new_n876));
  INV_X1    g690(.A(new_n873), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n850), .A2(new_n767), .A3(new_n853), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n848), .B1(new_n878), .B2(new_n857), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n871), .A2(new_n588), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT48), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n847), .A2(new_n874), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n777), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NAND4_X1  g699(.A1(new_n832), .A2(G210), .A3(G902), .A4(new_n841), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n324), .A2(new_n326), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n336), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n266), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n837), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n827), .A2(KEYINPUT114), .A3(new_n828), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n836), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n815), .A3(new_n800), .A4(new_n803), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n896), .B1(KEYINPUT53), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(G210), .A4(G902), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n904), .A2(KEYINPUT119), .A3(new_n906), .A4(new_n905), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n895), .B1(new_n909), .B2(new_n910), .ZN(G51));
  XOR2_X1   g725(.A(new_n740), .B(KEYINPUT57), .Z(new_n912));
  NOR2_X1   g726(.A1(new_n842), .A2(new_n779), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n778), .B1(new_n832), .B2(new_n841), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n664), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n832), .A2(G902), .A3(new_n841), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n737), .A3(new_n732), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n893), .B1(new_n916), .B2(new_n918), .ZN(G54));
  AOI21_X1  g733(.A(KEYINPUT120), .B1(KEYINPUT58), .B2(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(KEYINPUT120), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n917), .A2(new_n413), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n413), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n832), .A2(G902), .A3(new_n841), .A4(new_n922), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n920), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n923), .A2(new_n894), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT121), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n923), .A2(new_n929), .A3(new_n926), .A4(new_n894), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(G60));
  NAND2_X1  g745(.A1(new_n599), .A2(new_n600), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n469), .A2(new_n283), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n932), .B1(new_n847), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n932), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n935), .C1(new_n913), .C2(new_n914), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n937), .A2(new_n894), .A3(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n902), .A2(new_n618), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n531), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n842), .B2(new_n942), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n946), .A3(new_n894), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(G953), .B1(new_n430), .B2(new_n333), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n814), .A2(new_n837), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n889), .B1(G898), .B2(new_n266), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  AOI21_X1  g768(.A(new_n266), .B1(G227), .B2(G900), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n551), .B(new_n408), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n716), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n812), .A2(new_n806), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n641), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n801), .A2(KEYINPUT62), .A3(new_n656), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n798), .A2(new_n656), .A3(new_n661), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n760), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n770), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n958), .B1(new_n968), .B2(G953), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n798), .A2(new_n661), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n760), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n801), .B(KEYINPUT123), .C1(new_n754), .C2(new_n759), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n534), .A2(new_n587), .A3(new_n679), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n747), .A2(new_n297), .A3(new_n640), .A4(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n976), .A2(new_n726), .A3(new_n728), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n974), .A2(new_n266), .A3(new_n770), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(G900), .A2(G953), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n957), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n969), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n969), .B2(new_n980), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n956), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n984), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n955), .A3(new_n982), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G72));
  NAND4_X1  g802(.A1(new_n974), .A2(new_n770), .A3(new_n951), .A4(new_n977), .ZN(new_n989));
  XNOR2_X1  g803(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n990));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n582), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n893), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n648), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n846), .A2(new_n582), .A3(new_n996), .A4(new_n992), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n966), .A2(new_n770), .A3(new_n967), .A4(new_n951), .ZN(new_n998));
  AOI211_X1 g812(.A(KEYINPUT126), .B(new_n996), .C1(new_n998), .C2(new_n992), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n992), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n648), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n995), .B(new_n997), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1001), .A2(new_n648), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(KEYINPUT126), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1001), .A2(new_n1000), .A3(new_n648), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1008), .A2(new_n1009), .A3(new_n997), .A4(new_n995), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1004), .A2(new_n1010), .ZN(G57));
endmodule


