

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739;

  INV_X2 U374 ( .A(G953), .ZN(n731) );
  XNOR2_X2 U375 ( .A(n468), .B(n440), .ZN(n507) );
  AND2_X2 U376 ( .A1(n394), .A2(n395), .ZN(n392) );
  XNOR2_X2 U377 ( .A(n389), .B(n439), .ZN(n468) );
  OR2_X2 U378 ( .A1(n643), .A2(G902), .ZN(n389) );
  XNOR2_X2 U379 ( .A(n464), .B(KEYINPUT94), .ZN(n728) );
  NOR2_X1 U380 ( .A1(n559), .A2(n658), .ZN(n545) );
  NOR2_X2 U381 ( .A1(n623), .A2(n589), .ZN(n352) );
  OR2_X1 U382 ( .A1(n635), .A2(G902), .ZN(n367) );
  AND2_X1 U383 ( .A1(n592), .A2(n591), .ZN(n602) );
  NOR2_X1 U384 ( .A1(n718), .A2(n593), .ZN(n603) );
  AND2_X1 U385 ( .A1(n501), .A2(n500), .ZN(n502) );
  AND2_X1 U386 ( .A1(n580), .A2(n706), .ZN(n556) );
  BUF_X1 U387 ( .A(n468), .Z(n559) );
  XNOR2_X1 U388 ( .A(n367), .B(n364), .ZN(n451) );
  XNOR2_X1 U389 ( .A(n387), .B(n385), .ZN(n437) );
  XNOR2_X1 U390 ( .A(n388), .B(G110), .ZN(n387) );
  XNOR2_X1 U391 ( .A(G107), .B(G104), .ZN(n388) );
  XNOR2_X2 U392 ( .A(n352), .B(n353), .ZN(n553) );
  NAND2_X1 U393 ( .A1(n416), .A2(G210), .ZN(n353) );
  BUF_X1 U394 ( .A(n709), .Z(n354) );
  XNOR2_X1 U395 ( .A(n467), .B(KEYINPUT31), .ZN(n709) );
  NOR2_X1 U396 ( .A1(n718), .A2(n593), .ZN(n355) );
  BUF_X1 U397 ( .A(n643), .Z(n356) );
  BUF_X1 U398 ( .A(n641), .Z(n357) );
  XNOR2_X1 U399 ( .A(n398), .B(n520), .ZN(n641) );
  AND2_X2 U400 ( .A1(n605), .A2(n604), .ZN(n358) );
  AND2_X2 U401 ( .A1(n605), .A2(n604), .ZN(n642) );
  XNOR2_X2 U402 ( .A(n432), .B(n431), .ZN(n464) );
  XNOR2_X1 U403 ( .A(n506), .B(n505), .ZN(n359) );
  XNOR2_X1 U404 ( .A(n390), .B(n393), .ZN(n360) );
  BUF_X1 U405 ( .A(n623), .Z(n361) );
  BUF_X1 U406 ( .A(n715), .Z(n362) );
  XNOR2_X1 U407 ( .A(n506), .B(n505), .ZN(n519) );
  XNOR2_X1 U408 ( .A(n390), .B(n393), .ZN(n718) );
  XNOR2_X2 U409 ( .A(n429), .B(KEYINPUT0), .ZN(n504) );
  NAND2_X1 U410 ( .A1(n641), .A2(n614), .ZN(n535) );
  NOR2_X1 U411 ( .A1(n674), .A2(n377), .ZN(n376) );
  INV_X1 U412 ( .A(KEYINPUT68), .ZN(n377) );
  NAND2_X1 U413 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X1 U414 ( .A1(n579), .A2(n578), .ZN(n382) );
  XNOR2_X1 U415 ( .A(n563), .B(KEYINPUT46), .ZN(n381) );
  NAND2_X1 U416 ( .A1(n363), .A2(KEYINPUT44), .ZN(n395) );
  AND2_X1 U417 ( .A1(n513), .A2(n694), .ZN(n394) );
  INV_X1 U418 ( .A(KEYINPUT4), .ZN(n399) );
  AND2_X1 U419 ( .A1(n545), .A2(n544), .ZN(n550) );
  NOR2_X1 U420 ( .A1(n662), .A2(n371), .ZN(n370) );
  INV_X1 U421 ( .A(n558), .ZN(n371) );
  NAND2_X1 U422 ( .A1(n374), .A2(n703), .ZN(n568) );
  XNOR2_X1 U423 ( .A(n375), .B(KEYINPUT47), .ZN(n374) );
  AND2_X1 U424 ( .A1(n704), .A2(n376), .ZN(n375) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n379) );
  INV_X1 U426 ( .A(KEYINPUT8), .ZN(n383) );
  NAND2_X1 U427 ( .A1(n731), .A2(G234), .ZN(n384) );
  OR2_X1 U428 ( .A1(n656), .A2(n655), .ZN(n658) );
  INV_X1 U429 ( .A(G902), .ZN(n538) );
  INV_X1 U430 ( .A(KEYINPUT45), .ZN(n393) );
  XNOR2_X1 U431 ( .A(n386), .B(G101), .ZN(n385) );
  INV_X1 U432 ( .A(KEYINPUT77), .ZN(n386) );
  NAND2_X1 U433 ( .A1(n656), .A2(n558), .ZN(n569) );
  XNOR2_X1 U434 ( .A(n552), .B(n551), .ZN(n567) );
  XNOR2_X1 U435 ( .A(n373), .B(n366), .ZN(n372) );
  NAND2_X1 U436 ( .A1(n609), .A2(G953), .ZN(n649) );
  NAND2_X1 U437 ( .A1(n519), .A2(n518), .ZN(n398) );
  OR2_X1 U438 ( .A1(n535), .A2(n615), .ZN(n363) );
  XOR2_X1 U439 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n364) );
  XOR2_X1 U440 ( .A(G113), .B(KEYINPUT3), .Z(n365) );
  XOR2_X1 U441 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n366) );
  XNOR2_X1 U442 ( .A(n728), .B(n438), .ZN(n643) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n378) );
  XNOR2_X2 U444 ( .A(n444), .B(n443), .ZN(n729) );
  XNOR2_X2 U445 ( .A(KEYINPUT40), .B(n556), .ZN(n739) );
  XNOR2_X1 U446 ( .A(n369), .B(n368), .ZN(n635) );
  XNOR2_X1 U447 ( .A(n729), .B(n442), .ZN(n368) );
  XNOR2_X1 U448 ( .A(n441), .B(n447), .ZN(n369) );
  NAND2_X1 U449 ( .A1(n370), .A2(n656), .ZN(n373) );
  NAND2_X1 U450 ( .A1(n560), .A2(n372), .ZN(n564) );
  NAND2_X1 U451 ( .A1(n378), .A2(n586), .ZN(n593) );
  XNOR2_X2 U452 ( .A(n384), .B(n383), .ZN(n493) );
  NAND2_X1 U453 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n396), .B(KEYINPUT70), .ZN(n391) );
  NAND2_X1 U455 ( .A1(n536), .A2(n537), .ZN(n396) );
  NOR2_X2 U456 ( .A1(n397), .A2(n428), .ZN(n429) );
  NOR2_X1 U457 ( .A1(n564), .A2(n397), .ZN(n704) );
  XNOR2_X2 U458 ( .A(n573), .B(n419), .ZN(n397) );
  XNOR2_X2 U459 ( .A(n492), .B(n399), .ZN(n432) );
  XNOR2_X2 U460 ( .A(n400), .B(n407), .ZN(n492) );
  XNOR2_X2 U461 ( .A(G143), .B(KEYINPUT64), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n533), .B(n532), .ZN(n615) );
  NOR2_X2 U463 ( .A1(n739), .A2(n738), .ZN(n563) );
  BUF_X1 U464 ( .A(n504), .Z(n526) );
  XOR2_X1 U465 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n401) );
  NOR2_X1 U466 ( .A1(n666), .A2(n665), .ZN(n402) );
  INV_X1 U467 ( .A(n674), .ZN(n500) );
  INV_X1 U468 ( .A(KEYINPUT86), .ZN(n534) );
  INV_X1 U469 ( .A(n711), .ZN(n578) );
  BUF_X1 U470 ( .A(n456), .Z(n462) );
  INV_X1 U471 ( .A(KEYINPUT78), .ZN(n551) );
  XNOR2_X1 U472 ( .A(G116), .B(G119), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n365), .B(n403), .ZN(n456) );
  XOR2_X1 U474 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n404) );
  XNOR2_X1 U475 ( .A(n404), .B(G122), .ZN(n405) );
  XNOR2_X1 U476 ( .A(n456), .B(n405), .ZN(n406) );
  XNOR2_X1 U477 ( .A(n437), .B(n406), .ZN(n715) );
  INV_X1 U478 ( .A(G128), .ZN(n407) );
  XNOR2_X2 U479 ( .A(G146), .B(G125), .ZN(n444) );
  XNOR2_X1 U480 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n408) );
  XNOR2_X1 U481 ( .A(n444), .B(n408), .ZN(n411) );
  NAND2_X1 U482 ( .A1(n731), .A2(G224), .ZN(n409) );
  XNOR2_X1 U483 ( .A(n409), .B(KEYINPUT90), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U485 ( .A(n432), .B(n412), .ZN(n413) );
  XNOR2_X1 U486 ( .A(n715), .B(n413), .ZN(n623) );
  XNOR2_X1 U487 ( .A(KEYINPUT89), .B(KEYINPUT15), .ZN(n414) );
  XNOR2_X1 U488 ( .A(n414), .B(n538), .ZN(n597) );
  INV_X1 U489 ( .A(n597), .ZN(n589) );
  INV_X1 U490 ( .A(G237), .ZN(n415) );
  NAND2_X1 U491 ( .A1(n538), .A2(n415), .ZN(n416) );
  NAND2_X1 U492 ( .A1(n416), .A2(G214), .ZN(n669) );
  NAND2_X1 U493 ( .A1(n553), .A2(n669), .ZN(n418) );
  INV_X1 U494 ( .A(KEYINPUT87), .ZN(n417) );
  XNOR2_X2 U495 ( .A(n418), .B(n417), .ZN(n573) );
  XNOR2_X1 U496 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n419) );
  XOR2_X1 U497 ( .A(KEYINPUT91), .B(KEYINPUT14), .Z(n421) );
  NAND2_X1 U498 ( .A1(G237), .A2(G234), .ZN(n420) );
  XNOR2_X1 U499 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U500 ( .A(KEYINPUT76), .B(n422), .Z(n423) );
  INV_X1 U501 ( .A(n423), .ZN(n542) );
  NAND2_X1 U502 ( .A1(G952), .A2(n542), .ZN(n681) );
  NOR2_X1 U503 ( .A1(n681), .A2(G953), .ZN(n427) );
  XOR2_X1 U504 ( .A(G898), .B(KEYINPUT92), .Z(n723) );
  NAND2_X1 U505 ( .A1(G953), .A2(n723), .ZN(n716) );
  NOR2_X1 U506 ( .A1(n423), .A2(n716), .ZN(n424) );
  NAND2_X1 U507 ( .A1(G902), .A2(n424), .ZN(n425) );
  XNOR2_X1 U508 ( .A(n425), .B(KEYINPUT93), .ZN(n426) );
  NOR2_X1 U509 ( .A1(n427), .A2(n426), .ZN(n428) );
  XNOR2_X1 U510 ( .A(G134), .B(G131), .ZN(n430) );
  XNOR2_X1 U511 ( .A(n430), .B(G137), .ZN(n431) );
  NAND2_X1 U512 ( .A1(n731), .A2(G227), .ZN(n433) );
  XNOR2_X1 U513 ( .A(n433), .B(G140), .ZN(n435) );
  XNOR2_X1 U514 ( .A(G146), .B(KEYINPUT79), .ZN(n434) );
  XNOR2_X1 U515 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U516 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U517 ( .A(KEYINPUT69), .B(G469), .ZN(n439) );
  XNOR2_X1 U518 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n440) );
  XOR2_X1 U519 ( .A(G119), .B(KEYINPUT24), .Z(n442) );
  NAND2_X1 U520 ( .A1(G221), .A2(n493), .ZN(n441) );
  XNOR2_X1 U521 ( .A(G140), .B(KEYINPUT10), .ZN(n443) );
  XOR2_X1 U522 ( .A(KEYINPUT23), .B(G137), .Z(n446) );
  XNOR2_X1 U523 ( .A(G128), .B(G110), .ZN(n445) );
  XNOR2_X1 U524 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U525 ( .A1(n597), .A2(G234), .ZN(n448) );
  XNOR2_X1 U526 ( .A(n448), .B(KEYINPUT20), .ZN(n452) );
  NAND2_X1 U527 ( .A1(n452), .A2(G217), .ZN(n449) );
  XNOR2_X1 U528 ( .A(KEYINPUT95), .B(n449), .ZN(n450) );
  XNOR2_X2 U529 ( .A(n451), .B(n450), .ZN(n656) );
  AND2_X1 U530 ( .A1(n452), .A2(G221), .ZN(n454) );
  XNOR2_X1 U531 ( .A(KEYINPUT97), .B(KEYINPUT21), .ZN(n453) );
  XNOR2_X1 U532 ( .A(n454), .B(n453), .ZN(n655) );
  INV_X1 U533 ( .A(n658), .ZN(n455) );
  NAND2_X1 U534 ( .A1(n507), .A2(n455), .ZN(n523) );
  XOR2_X1 U535 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n458) );
  XNOR2_X1 U536 ( .A(G101), .B(G146), .ZN(n457) );
  XNOR2_X1 U537 ( .A(n458), .B(n457), .ZN(n460) );
  NOR2_X1 U538 ( .A1(G953), .A2(G237), .ZN(n471) );
  NAND2_X1 U539 ( .A1(n471), .A2(G210), .ZN(n459) );
  XNOR2_X1 U540 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U541 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U542 ( .A(n464), .B(n463), .ZN(n618) );
  OR2_X1 U543 ( .A1(n618), .A2(G902), .ZN(n466) );
  INV_X1 U544 ( .A(G472), .ZN(n465) );
  XNOR2_X2 U545 ( .A(n466), .B(n465), .ZN(n662) );
  NOR2_X1 U546 ( .A1(n523), .A2(n662), .ZN(n665) );
  NAND2_X1 U547 ( .A1(n504), .A2(n665), .ZN(n467) );
  AND2_X1 U548 ( .A1(n545), .A2(n662), .ZN(n469) );
  AND2_X1 U549 ( .A1(n526), .A2(n469), .ZN(n696) );
  NOR2_X2 U550 ( .A1(n709), .A2(n696), .ZN(n470) );
  XNOR2_X1 U551 ( .A(n470), .B(KEYINPUT99), .ZN(n501) );
  XOR2_X1 U552 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n473) );
  NAND2_X1 U553 ( .A1(n471), .A2(G214), .ZN(n472) );
  XNOR2_X1 U554 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U555 ( .A(n474), .B(KEYINPUT101), .Z(n476) );
  XNOR2_X1 U556 ( .A(G143), .B(G131), .ZN(n475) );
  XNOR2_X1 U557 ( .A(n476), .B(n475), .ZN(n481) );
  XOR2_X1 U558 ( .A(KEYINPUT11), .B(G113), .Z(n478) );
  XNOR2_X1 U559 ( .A(G122), .B(G104), .ZN(n477) );
  XNOR2_X1 U560 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U561 ( .A(n729), .B(n479), .ZN(n480) );
  XNOR2_X1 U562 ( .A(n481), .B(n480), .ZN(n606) );
  NAND2_X1 U563 ( .A1(n606), .A2(n538), .ZN(n485) );
  XOR2_X1 U564 ( .A(KEYINPUT103), .B(KEYINPUT13), .Z(n483) );
  XNOR2_X1 U565 ( .A(KEYINPUT102), .B(G475), .ZN(n482) );
  XOR2_X1 U566 ( .A(n483), .B(n482), .Z(n484) );
  XNOR2_X1 U567 ( .A(n485), .B(n484), .ZN(n530) );
  XOR2_X1 U568 ( .A(G122), .B(G116), .Z(n487) );
  XNOR2_X1 U569 ( .A(G134), .B(G107), .ZN(n486) );
  XNOR2_X1 U570 ( .A(n487), .B(n486), .ZN(n491) );
  XOR2_X1 U571 ( .A(KEYINPUT7), .B(KEYINPUT104), .Z(n489) );
  XNOR2_X1 U572 ( .A(KEYINPUT9), .B(KEYINPUT105), .ZN(n488) );
  XNOR2_X1 U573 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U574 ( .A(n491), .B(n490), .Z(n496) );
  NAND2_X1 U575 ( .A1(G217), .A2(n493), .ZN(n494) );
  XNOR2_X1 U576 ( .A(n492), .B(n494), .ZN(n495) );
  XNOR2_X1 U577 ( .A(n496), .B(n495), .ZN(n630) );
  NAND2_X1 U578 ( .A1(n630), .A2(n538), .ZN(n498) );
  XNOR2_X1 U579 ( .A(KEYINPUT106), .B(G478), .ZN(n497) );
  XNOR2_X1 U580 ( .A(n498), .B(n497), .ZN(n529) );
  INV_X1 U581 ( .A(n529), .ZN(n499) );
  AND2_X1 U582 ( .A1(n530), .A2(n499), .ZN(n706) );
  NOR2_X1 U583 ( .A1(n530), .A2(n499), .ZN(n708) );
  NOR2_X1 U584 ( .A1(n706), .A2(n708), .ZN(n674) );
  XNOR2_X1 U585 ( .A(n502), .B(KEYINPUT107), .ZN(n513) );
  OR2_X1 U586 ( .A1(n530), .A2(n529), .ZN(n672) );
  NOR2_X1 U587 ( .A1(n672), .A2(n655), .ZN(n503) );
  NAND2_X1 U588 ( .A1(n503), .A2(n504), .ZN(n506) );
  XNOR2_X1 U589 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n505) );
  BUF_X1 U590 ( .A(n507), .Z(n508) );
  INV_X1 U591 ( .A(KEYINPUT108), .ZN(n509) );
  XNOR2_X1 U592 ( .A(n509), .B(KEYINPUT6), .ZN(n510) );
  XNOR2_X1 U593 ( .A(n662), .B(n510), .ZN(n514) );
  INV_X1 U594 ( .A(n656), .ZN(n515) );
  NAND2_X1 U595 ( .A1(n514), .A2(n515), .ZN(n511) );
  NOR2_X1 U596 ( .A1(n508), .A2(n511), .ZN(n512) );
  NAND2_X1 U597 ( .A1(n359), .A2(n512), .ZN(n694) );
  INV_X1 U598 ( .A(n514), .ZN(n571) );
  NOR2_X1 U599 ( .A1(n571), .A2(n515), .ZN(n516) );
  NAND2_X1 U600 ( .A1(n508), .A2(n516), .ZN(n517) );
  XNOR2_X1 U601 ( .A(n517), .B(KEYINPUT81), .ZN(n518) );
  XNOR2_X1 U602 ( .A(KEYINPUT80), .B(KEYINPUT32), .ZN(n520) );
  NAND2_X1 U603 ( .A1(n656), .A2(n662), .ZN(n521) );
  NOR2_X1 U604 ( .A1(n508), .A2(n521), .ZN(n522) );
  NAND2_X1 U605 ( .A1(n359), .A2(n522), .ZN(n614) );
  XNOR2_X1 U606 ( .A(n523), .B(KEYINPUT109), .ZN(n524) );
  NAND2_X1 U607 ( .A1(n524), .A2(n571), .ZN(n525) );
  XNOR2_X1 U608 ( .A(n525), .B(KEYINPUT33), .ZN(n668) );
  NAND2_X1 U609 ( .A1(n668), .A2(n526), .ZN(n528) );
  XNOR2_X1 U610 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n527) );
  XNOR2_X1 U611 ( .A(n528), .B(n527), .ZN(n531) );
  NAND2_X1 U612 ( .A1(n530), .A2(n529), .ZN(n565) );
  NOR2_X2 U613 ( .A1(n531), .A2(n565), .ZN(n533) );
  XNOR2_X1 U614 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n532) );
  NOR2_X1 U615 ( .A1(n615), .A2(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U616 ( .A(n535), .B(n534), .ZN(n536) );
  NOR2_X1 U617 ( .A1(G900), .A2(n538), .ZN(n539) );
  NOR2_X1 U618 ( .A1(n731), .A2(n539), .ZN(n541) );
  NOR2_X1 U619 ( .A1(G953), .A2(G952), .ZN(n540) );
  NOR2_X1 U620 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U621 ( .A1(n543), .A2(n542), .ZN(n557) );
  INV_X1 U622 ( .A(n557), .ZN(n544) );
  INV_X1 U623 ( .A(n662), .ZN(n546) );
  NAND2_X1 U624 ( .A1(n546), .A2(n669), .ZN(n548) );
  XOR2_X1 U625 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n547) );
  XNOR2_X1 U626 ( .A(n548), .B(n547), .ZN(n549) );
  NAND2_X1 U627 ( .A1(n550), .A2(n549), .ZN(n552) );
  INV_X1 U628 ( .A(KEYINPUT38), .ZN(n554) );
  XNOR2_X1 U629 ( .A(n554), .B(n553), .ZN(n670) );
  NAND2_X1 U630 ( .A1(n567), .A2(n670), .ZN(n555) );
  XNOR2_X1 U631 ( .A(n555), .B(n401), .ZN(n580) );
  NOR2_X1 U632 ( .A1(n655), .A2(n557), .ZN(n558) );
  XNOR2_X1 U633 ( .A(n559), .B(KEYINPUT111), .ZN(n560) );
  NAND2_X1 U634 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U635 ( .A1(n672), .A2(n673), .ZN(n561) );
  XNOR2_X1 U636 ( .A(n561), .B(KEYINPUT41), .ZN(n684) );
  NOR2_X1 U637 ( .A1(n564), .A2(n684), .ZN(n562) );
  XNOR2_X1 U638 ( .A(KEYINPUT42), .B(n562), .ZN(n738) );
  INV_X1 U639 ( .A(n553), .ZN(n584) );
  NOR2_X1 U640 ( .A1(n584), .A2(n565), .ZN(n566) );
  NAND2_X1 U641 ( .A1(n567), .A2(n566), .ZN(n703) );
  XNOR2_X1 U642 ( .A(n568), .B(KEYINPUT75), .ZN(n579) );
  INV_X1 U643 ( .A(n706), .ZN(n570) );
  NOR2_X1 U644 ( .A1(n570), .A2(n569), .ZN(n572) );
  AND2_X1 U645 ( .A1(n572), .A2(n571), .ZN(n581) );
  INV_X1 U646 ( .A(n573), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n581), .A2(n574), .ZN(n576) );
  INV_X1 U648 ( .A(KEYINPUT36), .ZN(n575) );
  XNOR2_X1 U649 ( .A(n576), .B(n575), .ZN(n577) );
  AND2_X1 U650 ( .A1(n577), .A2(n508), .ZN(n711) );
  AND2_X1 U651 ( .A1(n580), .A2(n708), .ZN(n714) );
  NAND2_X1 U652 ( .A1(n581), .A2(n669), .ZN(n582) );
  OR2_X1 U653 ( .A1(n582), .A2(n508), .ZN(n583) );
  XNOR2_X1 U654 ( .A(n583), .B(KEYINPUT43), .ZN(n585) );
  AND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n613) );
  NOR2_X1 U656 ( .A1(n714), .A2(n613), .ZN(n586) );
  INV_X1 U657 ( .A(KEYINPUT83), .ZN(n587) );
  AND2_X1 U658 ( .A1(n587), .A2(n589), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n603), .A2(n588), .ZN(n592) );
  NAND2_X1 U660 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n590) );
  OR2_X1 U661 ( .A1(n597), .A2(n590), .ZN(n591) );
  NOR2_X1 U662 ( .A1(n360), .A2(n597), .ZN(n595) );
  INV_X1 U663 ( .A(n593), .ZN(n730) );
  NAND2_X1 U664 ( .A1(n730), .A2(KEYINPUT83), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n600) );
  INV_X1 U666 ( .A(KEYINPUT2), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U668 ( .A1(n598), .A2(KEYINPUT66), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n355), .A2(KEYINPUT2), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n358), .A2(G475), .ZN(n608) );
  XOR2_X1 U673 ( .A(n606), .B(KEYINPUT59), .Z(n607) );
  XNOR2_X1 U674 ( .A(n608), .B(n607), .ZN(n610) );
  INV_X1 U675 ( .A(G952), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n610), .A2(n649), .ZN(n612) );
  INV_X1 U677 ( .A(KEYINPUT60), .ZN(n611) );
  XNOR2_X1 U678 ( .A(n612), .B(n611), .ZN(G60) );
  XOR2_X1 U679 ( .A(n613), .B(G140), .Z(G42) );
  XNOR2_X1 U680 ( .A(n614), .B(G110), .ZN(G12) );
  XNOR2_X1 U681 ( .A(G122), .B(KEYINPUT126), .ZN(n616) );
  XOR2_X1 U682 ( .A(n616), .B(n615), .Z(G24) );
  NAND2_X1 U683 ( .A1(n358), .A2(G472), .ZN(n620) );
  XOR2_X1 U684 ( .A(KEYINPUT88), .B(KEYINPUT62), .Z(n617) );
  XNOR2_X1 U685 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U686 ( .A(n620), .B(n619), .ZN(n621) );
  NAND2_X1 U687 ( .A1(n621), .A2(n649), .ZN(n622) );
  XNOR2_X1 U688 ( .A(n622), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U689 ( .A1(n642), .A2(G210), .ZN(n626) );
  XNOR2_X1 U690 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n624) );
  XNOR2_X1 U691 ( .A(n361), .B(n624), .ZN(n625) );
  XNOR2_X1 U692 ( .A(n626), .B(n625), .ZN(n627) );
  NAND2_X1 U693 ( .A1(n627), .A2(n649), .ZN(n629) );
  INV_X1 U694 ( .A(KEYINPUT56), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n629), .B(n628), .ZN(G51) );
  NAND2_X1 U696 ( .A1(n642), .A2(G478), .ZN(n631) );
  XNOR2_X1 U697 ( .A(n631), .B(n630), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n632), .A2(n649), .ZN(n634) );
  INV_X1 U699 ( .A(KEYINPUT120), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n634), .B(n633), .ZN(G63) );
  NAND2_X1 U701 ( .A1(n642), .A2(G217), .ZN(n637) );
  XNOR2_X1 U702 ( .A(n635), .B(KEYINPUT121), .ZN(n636) );
  XNOR2_X1 U703 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U704 ( .A1(n638), .A2(n649), .ZN(n640) );
  INV_X1 U705 ( .A(KEYINPUT122), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n640), .B(n639), .ZN(G66) );
  XNOR2_X1 U707 ( .A(n357), .B(G119), .ZN(G21) );
  NAND2_X1 U708 ( .A1(n358), .A2(G469), .ZN(n648) );
  XOR2_X1 U709 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n645) );
  XNOR2_X1 U710 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n644) );
  XOR2_X1 U711 ( .A(n645), .B(n644), .Z(n646) );
  XNOR2_X1 U712 ( .A(n356), .B(n646), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n648), .B(n647), .ZN(n651) );
  INV_X1 U714 ( .A(n649), .ZN(n650) );
  NOR2_X1 U715 ( .A1(n651), .A2(n650), .ZN(G54) );
  INV_X1 U716 ( .A(n355), .ZN(n652) );
  NAND2_X1 U717 ( .A1(n652), .A2(KEYINPUT82), .ZN(n654) );
  XNOR2_X1 U718 ( .A(KEYINPUT2), .B(KEYINPUT84), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n654), .B(n653), .ZN(n690) );
  NAND2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U721 ( .A(n657), .B(KEYINPUT49), .ZN(n664) );
  INV_X1 U722 ( .A(n508), .ZN(n659) );
  NAND2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U724 ( .A(n660), .B(KEYINPUT50), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n664), .A2(n663), .ZN(n666) );
  XOR2_X1 U727 ( .A(KEYINPUT51), .B(n402), .Z(n667) );
  NOR2_X1 U728 ( .A1(n684), .A2(n667), .ZN(n679) );
  INV_X1 U729 ( .A(n668), .ZN(n683) );
  NOR2_X1 U730 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U731 ( .A1(n672), .A2(n671), .ZN(n676) );
  NOR2_X1 U732 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U733 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U734 ( .A1(n683), .A2(n677), .ZN(n678) );
  NOR2_X1 U735 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U736 ( .A(n680), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U737 ( .A1(n682), .A2(n681), .ZN(n688) );
  NOR2_X1 U738 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U739 ( .A(n685), .B(KEYINPUT115), .ZN(n686) );
  NAND2_X1 U740 ( .A1(n686), .A2(n731), .ZN(n687) );
  NOR2_X1 U741 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U742 ( .A1(n690), .A2(n689), .ZN(n693) );
  XNOR2_X1 U743 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n691) );
  XNOR2_X1 U744 ( .A(n691), .B(KEYINPUT116), .ZN(n692) );
  XNOR2_X1 U745 ( .A(n693), .B(n692), .ZN(G75) );
  XNOR2_X1 U746 ( .A(G101), .B(n694), .ZN(G3) );
  NAND2_X1 U747 ( .A1(n696), .A2(n706), .ZN(n695) );
  XNOR2_X1 U748 ( .A(n695), .B(G104), .ZN(G6) );
  XOR2_X1 U749 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n698) );
  NAND2_X1 U750 ( .A1(n696), .A2(n708), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n698), .B(n697), .ZN(n700) );
  XOR2_X1 U752 ( .A(G107), .B(KEYINPUT27), .Z(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(G9) );
  XOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .Z(n702) );
  NAND2_X1 U755 ( .A1(n704), .A2(n708), .ZN(n701) );
  XNOR2_X1 U756 ( .A(n702), .B(n701), .ZN(G30) );
  XNOR2_X1 U757 ( .A(G143), .B(n703), .ZN(G45) );
  NAND2_X1 U758 ( .A1(n704), .A2(n706), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n705), .B(G146), .ZN(G48) );
  NAND2_X1 U760 ( .A1(n354), .A2(n706), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n707), .B(G113), .ZN(G15) );
  NAND2_X1 U762 ( .A1(n354), .A2(n708), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n710), .B(G116), .ZN(G18) );
  XNOR2_X1 U764 ( .A(n711), .B(KEYINPUT37), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n712), .B(KEYINPUT114), .ZN(n713) );
  XNOR2_X1 U766 ( .A(G125), .B(n713), .ZN(G27) );
  XOR2_X1 U767 ( .A(G134), .B(n714), .Z(G36) );
  XNOR2_X1 U768 ( .A(n362), .B(KEYINPUT125), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n727) );
  NOR2_X1 U770 ( .A1(n360), .A2(G953), .ZN(n725) );
  XOR2_X1 U771 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n720) );
  NAND2_X1 U772 ( .A1(G224), .A2(G953), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  XOR2_X1 U774 ( .A(KEYINPUT123), .B(n721), .Z(n722) );
  NOR2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U777 ( .A(n727), .B(n726), .ZN(G69) );
  XNOR2_X1 U778 ( .A(n728), .B(n729), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n730), .B(n733), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(n731), .ZN(n737) );
  XOR2_X1 U781 ( .A(G227), .B(n733), .Z(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(G900), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U785 ( .A(G137), .B(n738), .Z(G39) );
  XOR2_X1 U786 ( .A(n739), .B(G131), .Z(G33) );
endmodule

