//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1170, new_n1171,
    new_n1172, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n220), .A2(new_n221), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n217), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT69), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n205), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n213), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n206), .A2(G1), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT70), .B1(new_n254), .B2(new_n255), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G150), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n206), .A2(G33), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n260), .B1(new_n201), .B2(new_n206), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n263), .A2(new_n252), .B1(new_n250), .B2(new_n255), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT9), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT73), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n273), .A2(G222), .B1(G77), .B2(new_n272), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT67), .B(G223), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n269), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(new_n280), .B2(new_n279), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT66), .B(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  AOI211_X1 g0085(.A(G1), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n287), .B2(new_n285), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n268), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(G226), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n266), .B(new_n267), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT72), .B(G200), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(new_n291), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(new_n291), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n265), .B1(new_n297), .B2(G169), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n291), .A2(G179), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT78), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n276), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n304));
  INV_X1    g0104(.A(G223), .ZN(new_n305));
  OR2_X1    g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n275), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n304), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n268), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n286), .B1(G232), .B2(new_n289), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(G169), .B1(new_n311), .B2(new_n313), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n303), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n316), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT78), .A3(new_n314), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G58), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XOR2_X1   g0125(.A(new_n325), .B(KEYINPUT76), .Z(new_n326));
  INV_X1    g0126(.A(G159), .ZN(new_n327));
  INV_X1    g0127(.A(new_n259), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT7), .B1(new_n272), .B2(new_n206), .ZN(new_n331));
  AND4_X1   g0131(.A1(KEYINPUT7), .A2(new_n306), .A3(new_n206), .A4(new_n307), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n322), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n329), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n330), .B1(new_n329), .B2(new_n334), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n252), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n261), .A2(new_n254), .ZN(new_n338));
  XOR2_X1   g0138(.A(new_n338), .B(KEYINPUT77), .Z(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n253), .B1(new_n250), .B2(new_n261), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n320), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT18), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n317), .A2(new_n319), .B1(new_n337), .B2(new_n340), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT18), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n311), .B2(new_n313), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n311), .A2(new_n313), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(G190), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n337), .A2(new_n340), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n343), .A2(new_n346), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n262), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(KEYINPUT71), .A3(new_n358), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n359), .B1(new_n206), .B2(new_n202), .C1(new_n328), .C2(new_n261), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT71), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n252), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n254), .A2(new_n202), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n253), .A2(new_n363), .B1(new_n202), .B2(new_n250), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n276), .A2(G238), .B1(G107), .B2(new_n272), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n308), .A2(G232), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(G1698), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n268), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n286), .B1(G244), .B2(new_n289), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n292), .ZN(new_n372));
  AOI211_X1 g0172(.A(new_n365), .B(new_n372), .C1(new_n371), .C2(new_n294), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n312), .A3(new_n370), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(new_n365), .A3(new_n376), .ZN(new_n377));
  OR3_X1    g0177(.A1(new_n355), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n249), .A2(G68), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT12), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n328), .A2(new_n255), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n262), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n252), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g0183(.A(new_n383), .B(KEYINPUT11), .Z(new_n384));
  NOR2_X1   g0184(.A1(new_n254), .A2(new_n322), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n380), .B(new_n384), .C1(new_n253), .C2(new_n385), .ZN(new_n386));
  XOR2_X1   g0186(.A(new_n386), .B(KEYINPUT75), .Z(new_n387));
  NAND2_X1  g0187(.A1(new_n273), .A2(G226), .ZN(new_n388));
  NAND3_X1  g0188(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT74), .B1(G33), .B2(G97), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n388), .B(new_n392), .C1(new_n275), .C2(new_n367), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n268), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n286), .B1(G238), .B2(new_n289), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT13), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT14), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(G169), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n312), .B2(new_n397), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n398), .B1(new_n397), .B2(G169), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n387), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n397), .A2(new_n292), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n397), .A2(G200), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n386), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n302), .A2(new_n378), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT81), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT66), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G41), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT5), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n205), .A2(G45), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n413), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT81), .B(new_n415), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n268), .A2(new_n418), .A3(new_n283), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  OAI211_X1 g0220(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n421));
  OAI211_X1 g0221(.A(G257), .B(new_n275), .C1(new_n270), .C2(new_n271), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n306), .A2(G303), .A3(new_n307), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n268), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n415), .B(new_n417), .C1(new_n284), .C2(KEYINPUT5), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(G270), .A3(new_n269), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n420), .A2(G179), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G283), .ZN(new_n429));
  INV_X1    g0229(.A(G97), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n206), .C1(G33), .C2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT85), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G33), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G97), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(KEYINPUT85), .A3(new_n206), .A4(new_n429), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G116), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G20), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n252), .A2(KEYINPUT84), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n252), .A2(new_n439), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT84), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n437), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT20), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n252), .A2(KEYINPUT84), .A3(new_n439), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT84), .B1(new_n252), .B2(new_n439), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n437), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(G116), .B1(new_n247), .B2(new_n248), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n252), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n205), .A2(G33), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n249), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n453), .B1(new_n456), .B2(new_n438), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n428), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT20), .B1(new_n449), .B2(new_n437), .ZN(new_n459));
  AND4_X1   g0259(.A1(KEYINPUT20), .A2(new_n437), .A3(new_n440), .A4(new_n443), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n420), .A2(new_n425), .A3(new_n427), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(G169), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT21), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n249), .A2(new_n454), .A3(new_n455), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n452), .B1(new_n466), .B2(G116), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n446), .B2(new_n450), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n462), .A2(G169), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT86), .B1(new_n470), .B2(KEYINPUT21), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT86), .ZN(new_n472));
  NOR4_X1   g0272(.A1(new_n468), .A2(new_n469), .A3(new_n472), .A4(new_n464), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n465), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n462), .A2(G200), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n468), .B(new_n476), .C1(new_n292), .C2(new_n462), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  AND2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G97), .A2(G107), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(KEYINPUT6), .A2(G97), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(G107), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(G97), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n489), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n490));
  OAI21_X1  g0290(.A(G107), .B1(new_n331), .B2(new_n332), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n454), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n250), .A2(new_n430), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n466), .B2(new_n430), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g0296(.A(G244), .B(new_n275), .C1(new_n270), .C2(new_n271), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT80), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n496), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n308), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(new_n429), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n268), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n426), .A2(G257), .A3(new_n269), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n420), .A2(KEYINPUT82), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT82), .B1(new_n420), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n495), .B1(new_n508), .B2(G200), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n420), .A2(new_n505), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT83), .B1(new_n512), .B2(new_n292), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n502), .A2(new_n429), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n499), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n269), .B1(new_n515), .B2(new_n501), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n510), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT83), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(G190), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n509), .A2(new_n513), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n504), .B(new_n312), .C1(new_n506), .C2(new_n507), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n374), .B1(new_n516), .B2(new_n510), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n495), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n525));
  OAI211_X1 g0325(.A(G250), .B(new_n275), .C1(new_n270), .C2(new_n271), .ZN(new_n526));
  INV_X1    g0326(.A(G294), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n526), .C1(new_n434), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n268), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n426), .A2(G264), .A3(new_n269), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT88), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(G179), .A4(new_n420), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n420), .A2(new_n529), .A3(new_n530), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n534), .A2(G169), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT88), .B1(new_n534), .B2(new_n312), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n206), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n308), .A2(new_n540), .A3(new_n206), .A4(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n206), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n487), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n358), .A2(G116), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n543), .B1(new_n542), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n252), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT87), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT87), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n252), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT25), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n249), .B2(G107), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n487), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n556), .A2(new_n557), .B1(new_n456), .B2(G107), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n537), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n558), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n534), .A2(new_n347), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G190), .B2(new_n534), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NOR3_X1   g0364(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT19), .B1(new_n390), .B2(new_n391), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n206), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n308), .A2(new_n206), .A3(G68), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n262), .B2(new_n430), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n252), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n456), .A2(new_n357), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n249), .A2(new_n357), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G238), .B(new_n275), .C1(new_n270), .C2(new_n271), .ZN(new_n577));
  OAI211_X1 g0377(.A(G244), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(new_n434), .C2(new_n438), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n268), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n413), .A2(G250), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n268), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n374), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n583), .B1(new_n579), .B2(new_n268), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n312), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n576), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n456), .A2(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n572), .A2(new_n590), .A3(new_n575), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n587), .A2(new_n294), .ZN(new_n592));
  AOI211_X1 g0392(.A(G190), .B(new_n583), .C1(new_n579), .C2(new_n268), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n589), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n564), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n407), .A2(new_n479), .A3(new_n524), .A4(new_n598), .ZN(G372));
  NAND2_X1  g0399(.A1(new_n343), .A2(new_n346), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n405), .A2(new_n377), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n402), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n353), .A2(new_n354), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n300), .B1(new_n604), .B2(new_n296), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT91), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G97), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT74), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n389), .ZN(new_n612));
  AOI21_X1  g0412(.A(G20), .B1(new_n612), .B2(KEYINPUT19), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n568), .B(new_n570), .C1(new_n613), .C2(new_n565), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n574), .B1(new_n614), .B2(new_n252), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n573), .B1(new_n312), .B2(new_n587), .ZN(new_n616));
  OAI21_X1  g0416(.A(KEYINPUT89), .B1(new_n587), .B2(G169), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n587), .A2(KEYINPUT89), .A3(G169), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n474), .A2(new_n559), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n554), .A2(new_n558), .A3(new_n563), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n591), .A2(KEYINPUT90), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT90), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n615), .A2(new_n624), .A3(new_n590), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n592), .A2(new_n593), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT89), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n585), .B2(new_n374), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n618), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n626), .A2(new_n627), .B1(new_n630), .B2(new_n616), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n520), .A2(new_n622), .A3(new_n523), .A4(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n620), .B1(new_n621), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n523), .B2(new_n595), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n624), .B1(new_n615), .B2(new_n590), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n624), .A2(new_n572), .A3(new_n590), .A4(new_n575), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n627), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n492), .A2(new_n494), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n512), .B2(new_n374), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n637), .A2(new_n620), .A3(new_n639), .A4(new_n521), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n634), .B1(new_n640), .B2(KEYINPUT26), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n608), .B1(new_n407), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g0443(.A(new_n643), .B(KEYINPUT92), .Z(G369));
  NAND3_X1  g0444(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n461), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n479), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n475), .B2(new_n651), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  INV_X1    g0454(.A(new_n650), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n564), .B1(new_n561), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n559), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n655), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n475), .A2(new_n650), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n564), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n559), .B2(new_n655), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(G399));
  NAND2_X1  g0464(.A1(new_n209), .A2(new_n284), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n205), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n565), .A2(new_n438), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n667), .A2(new_n669), .B1(new_n216), .B2(new_n666), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT28), .Z(new_n671));
  NAND2_X1  g0471(.A1(new_n642), .A2(new_n655), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT29), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n523), .B2(new_n595), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n640), .B2(new_n675), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n620), .B(new_n677), .C1(new_n621), .C2(new_n632), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n678), .A2(KEYINPUT93), .A3(new_n655), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT93), .B1(new_n678), .B2(new_n655), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT29), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n598), .A2(new_n479), .A3(new_n524), .A4(new_n655), .ZN(new_n682));
  INV_X1    g0482(.A(new_n428), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n517), .A2(new_n683), .A3(new_n531), .A4(new_n587), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n312), .A2(new_n534), .A3(new_n462), .A4(new_n585), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n684), .A2(new_n685), .B1(new_n508), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n685), .B2(new_n684), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n650), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT31), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n674), .A2(new_n681), .B1(G330), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n671), .B1(new_n692), .B2(G1), .ZN(G364));
  NAND2_X1  g0493(.A1(new_n206), .A2(G13), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT94), .Z(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G45), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n667), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n654), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(G330), .B2(new_n653), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n209), .A2(new_n308), .ZN(new_n701));
  INV_X1    g0501(.A(G355), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n701), .A2(new_n702), .B1(G116), .B2(new_n209), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n240), .A2(new_n285), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n209), .A2(new_n272), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n285), .B2(new_n216), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n703), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(G20), .B1(KEYINPUT95), .B2(G169), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(KEYINPUT95), .A2(G169), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n213), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n698), .B1(new_n707), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n206), .A2(new_n292), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n312), .A2(G200), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G322), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n272), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n294), .A2(new_n312), .A3(new_n718), .ZN(new_n723));
  INV_X1    g0523(.A(G303), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n206), .A2(G190), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G179), .A2(G200), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n722), .B(new_n725), .C1(G329), .C2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G283), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n294), .A2(new_n312), .A3(new_n726), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n312), .A2(new_n347), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT97), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n733), .A2(new_n734), .A3(new_n726), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n734), .B1(new_n733), .B2(new_n726), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(KEYINPUT33), .B(G317), .Z(new_n738));
  OAI221_X1 g0538(.A(new_n730), .B1(new_n731), .B2(new_n732), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n718), .A2(new_n733), .ZN(new_n740));
  INV_X1    g0540(.A(G326), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n719), .A2(new_n726), .ZN(new_n742));
  INV_X1    g0542(.A(G311), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n740), .A2(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n206), .B1(new_n727), .B2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n744), .B1(G294), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT98), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n308), .B1(new_n742), .B2(new_n202), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n740), .A2(new_n255), .B1(new_n720), .B2(new_n321), .ZN(new_n750));
  INV_X1    g0550(.A(new_n723), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n749), .B(new_n750), .C1(G87), .C2(new_n751), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n752), .B1(new_n322), .B2(new_n737), .C1(new_n487), .C2(new_n732), .ZN(new_n753));
  XOR2_X1   g0553(.A(KEYINPUT96), .B(G159), .Z(new_n754));
  OR3_X1    g0554(.A1(new_n754), .A2(new_n728), .A3(KEYINPUT32), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT32), .B1(new_n754), .B2(new_n728), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n755), .B(new_n756), .C1(new_n430), .C2(new_n745), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n739), .A2(new_n748), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n717), .B1(new_n758), .B2(new_n711), .ZN(new_n759));
  INV_X1    g0559(.A(new_n714), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n653), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n700), .A2(new_n761), .ZN(G396));
  NAND2_X1  g0562(.A1(new_n377), .A2(new_n655), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n373), .B1(new_n365), .B2(new_n650), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n377), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n672), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n765), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n642), .A2(new_n767), .A3(new_n655), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n691), .A2(G330), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n698), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n711), .A2(new_n712), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n697), .B1(new_n202), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n711), .ZN(new_n775));
  INV_X1    g0575(.A(new_n732), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G87), .A2(new_n776), .B1(new_n751), .B2(G107), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n731), .B2(new_n737), .ZN(new_n778));
  INV_X1    g0578(.A(new_n720), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G294), .A2(new_n779), .B1(new_n729), .B2(G311), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n438), .B2(new_n742), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n272), .B1(new_n745), .B2(new_n430), .C1(new_n740), .C2(new_n724), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n778), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n740), .ZN(new_n784));
  INV_X1    g0584(.A(new_n754), .ZN(new_n785));
  INV_X1    g0585(.A(new_n742), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G137), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G143), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n720), .ZN(new_n789));
  INV_X1    g0589(.A(new_n737), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G150), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(KEYINPUT34), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G68), .A2(new_n776), .B1(new_n751), .B2(G50), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT99), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n308), .B1(new_n745), .B2(new_n321), .C1(new_n798), .C2(new_n728), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n791), .B2(KEYINPUT34), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n783), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n774), .B1(new_n775), .B2(new_n801), .C1(new_n767), .C2(new_n713), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n772), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G384));
  OR2_X1    g0604(.A1(new_n489), .A2(KEYINPUT35), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n489), .A2(KEYINPUT35), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n805), .A2(G116), .A3(new_n214), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT36), .Z(new_n808));
  OAI211_X1 g0608(.A(new_n216), .B(G77), .C1(new_n321), .C2(new_n322), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n255), .A2(G68), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n205), .B(G13), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT40), .ZN(new_n813));
  INV_X1    g0613(.A(new_n401), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n814), .B(new_n399), .C1(new_n312), .C2(new_n397), .ZN(new_n815));
  INV_X1    g0615(.A(new_n405), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n387), .B(new_n650), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n387), .A2(new_n650), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n402), .A2(new_n405), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n767), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n648), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n341), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n343), .A2(new_n346), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n603), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT38), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n342), .A2(new_n824), .A3(new_n351), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n342), .A2(new_n824), .A3(KEYINPUT37), .A4(new_n351), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n826), .A2(new_n827), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n832), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n355), .A2(new_n341), .A3(new_n823), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT38), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n822), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT102), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n691), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n682), .A2(new_n690), .A3(KEYINPUT102), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n813), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n827), .B1(new_n826), .B2(new_n832), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT38), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n821), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n846), .A3(KEYINPUT40), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n843), .A2(new_n407), .ZN(new_n849));
  OAI21_X1  g0649(.A(G330), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n833), .B2(new_n836), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n815), .A2(new_n387), .A3(new_n655), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT101), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n844), .A2(KEYINPUT39), .A3(new_n845), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n763), .B(KEYINPUT100), .Z(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n768), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n860), .B(new_n820), .C1(new_n833), .C2(new_n836), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n600), .A2(new_n648), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n857), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n407), .A2(new_n681), .A3(new_n674), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n607), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n863), .B(new_n865), .Z(new_n866));
  OAI22_X1  g0666(.A1(new_n851), .A2(new_n866), .B1(new_n205), .B2(new_n695), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n851), .A2(new_n866), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n812), .B1(new_n867), .B2(new_n868), .ZN(G367));
  OAI21_X1  g0669(.A(new_n524), .B1(new_n638), .B2(new_n655), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT103), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n523), .B2(new_n655), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n662), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n523), .B1(new_n871), .B2(new_n657), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(KEYINPUT42), .B1(new_n655), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(KEYINPUT104), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n875), .B2(KEYINPUT104), .ZN(new_n879));
  OR3_X1    g0679(.A1(new_n626), .A2(new_n620), .A3(new_n655), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n631), .B1(new_n626), .B2(new_n655), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n877), .A2(new_n879), .B1(KEYINPUT43), .B2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n654), .A2(new_n872), .A3(new_n658), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n665), .B(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n872), .A2(new_n663), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT45), .Z(new_n894));
  INV_X1    g0694(.A(KEYINPUT106), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(KEYINPUT44), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n872), .A2(new_n663), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(KEYINPUT44), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n894), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT107), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(new_n659), .Z(new_n904));
  OAI21_X1  g0704(.A(new_n661), .B1(new_n658), .B2(new_n660), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n654), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n692), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT108), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n892), .B1(new_n910), .B2(new_n692), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n696), .A2(G1), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n889), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n236), .A2(new_n705), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n715), .B1(new_n209), .B2(new_n356), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n698), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT109), .ZN(new_n917));
  INV_X1    g0717(.A(G317), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n720), .A2(new_n724), .B1(new_n728), .B2(new_n918), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n272), .B1(new_n745), .B2(new_n487), .C1(new_n740), .C2(new_n743), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(G283), .C2(new_n786), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n921), .B1(new_n430), .B2(new_n732), .C1(new_n527), .C2(new_n737), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n723), .A2(new_n438), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT46), .ZN(new_n924));
  INV_X1    g0724(.A(G137), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n308), .B1(new_n728), .B2(new_n925), .C1(new_n255), .C2(new_n742), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(G77), .B2(new_n776), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n321), .B2(new_n723), .C1(new_n737), .C2(new_n754), .ZN(new_n928));
  INV_X1    g0728(.A(G150), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n740), .A2(new_n788), .B1(new_n720), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n745), .A2(new_n322), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT110), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n922), .A2(new_n924), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT47), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n711), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n917), .B1(new_n882), .B2(new_n760), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n913), .A2(new_n939), .ZN(G387));
  OR2_X1    g0740(.A1(new_n658), .A2(new_n760), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n701), .A2(new_n669), .B1(G107), .B2(new_n209), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT111), .Z(new_n943));
  OR2_X1    g0743(.A1(new_n233), .A2(new_n285), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n261), .A2(G50), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT50), .ZN(new_n946));
  AOI211_X1 g0746(.A(G45), .B(new_n668), .C1(G68), .C2(G77), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n705), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n943), .B1(new_n944), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n698), .B1(new_n949), .B2(new_n716), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n308), .B1(new_n720), .B2(new_n255), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n742), .A2(new_n322), .B1(new_n728), .B2(new_n929), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n357), .C2(new_n746), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n784), .A2(G159), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT112), .ZN(new_n955));
  INV_X1    g0755(.A(new_n261), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n790), .A2(new_n956), .B1(G97), .B2(new_n776), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n751), .A2(G77), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n953), .A2(new_n955), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n308), .B1(new_n729), .B2(G326), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n723), .A2(new_n527), .B1(new_n731), .B2(new_n745), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT113), .B(G322), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n784), .A2(new_n963), .B1(new_n786), .B2(G303), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n918), .B2(new_n720), .C1(new_n737), .C2(new_n743), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT48), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n965), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT49), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n960), .B1(new_n438), .B2(new_n732), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n959), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n950), .B1(new_n972), .B2(new_n711), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n906), .A2(new_n912), .B1(new_n941), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n666), .B1(new_n906), .B2(new_n692), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n909), .B2(new_n975), .ZN(G393));
  XNOR2_X1  g0776(.A(new_n901), .B(new_n659), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n910), .B(new_n666), .C1(new_n909), .C2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n872), .A2(new_n760), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n243), .A2(new_n705), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n715), .B1(new_n430), .B2(new_n209), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n698), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n740), .A2(new_n929), .B1(new_n720), .B2(new_n327), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT51), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n308), .B1(new_n728), .B2(new_n788), .C1(new_n261), .C2(new_n742), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G77), .B2(new_n746), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n790), .A2(G50), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G87), .A2(new_n776), .B1(new_n751), .B2(G68), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n740), .A2(new_n918), .B1(new_n720), .B2(new_n743), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT52), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n728), .A2(new_n962), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n272), .B1(new_n742), .B2(new_n527), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G116), .C2(new_n746), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n790), .A2(G303), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G107), .A2(new_n776), .B1(new_n751), .B2(G283), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n991), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n989), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n982), .B1(new_n998), .B2(new_n711), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n977), .A2(new_n912), .B1(new_n979), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n978), .A2(new_n1000), .ZN(G390));
  NAND2_X1  g0801(.A1(new_n853), .A2(new_n856), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n855), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n860), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n820), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n691), .A2(G330), .A3(new_n767), .A4(new_n820), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n678), .A2(new_n655), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT93), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n678), .A2(KEYINPUT93), .A3(new_n655), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n765), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(KEYINPUT114), .B1(new_n1013), .B2(new_n858), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n767), .B1(new_n679), .B2(new_n680), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT114), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n859), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n820), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT115), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n855), .B1(new_n844), .B2(new_n845), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1019), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1007), .B(new_n1008), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(KEYINPUT115), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n839), .A2(G330), .A3(new_n767), .A4(new_n840), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n820), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1023), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n912), .ZN(new_n1033));
  OAI21_X1  g0833(.A(KEYINPUT117), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1007), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n820), .A3(new_n1030), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT117), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1036), .A2(new_n1037), .A3(new_n912), .A4(new_n1023), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1002), .A2(new_n712), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n773), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1040), .A2(new_n956), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n742), .A2(new_n430), .B1(new_n728), .B2(new_n527), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n272), .B1(new_n745), .B2(new_n202), .C1(new_n740), .C2(new_n731), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G116), .C2(new_n779), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G68), .A2(new_n776), .B1(new_n751), .B2(G87), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n487), .C2(new_n737), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n751), .A2(G150), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT53), .ZN(new_n1048));
  INV_X1    g0848(.A(G128), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n308), .B1(new_n740), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(G125), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n720), .A2(new_n798), .B1(new_n728), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G159), .C2(new_n746), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n790), .A2(G137), .B1(G50), .B2(new_n776), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(KEYINPUT54), .B(G143), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT118), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1053), .B(new_n1054), .C1(new_n742), .C2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1046), .B1(new_n1048), .B2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n697), .B(new_n1041), .C1(new_n1059), .C2(new_n711), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1034), .A2(new_n1038), .B1(new_n1039), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT116), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1005), .B1(new_n770), .B2(new_n765), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1029), .B2(new_n1005), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n860), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1029), .A2(new_n1005), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n1067), .A3(new_n1008), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n843), .A2(G330), .A3(new_n407), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n607), .A3(new_n864), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1032), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1071), .B1(new_n1068), .B2(new_n1065), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1023), .B(new_n1075), .C1(new_n1028), .C2(new_n1031), .ZN(new_n1076));
  AND4_X1   g0876(.A1(new_n1062), .A2(new_n1074), .A3(new_n666), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n665), .B1(new_n1032), .B2(new_n1073), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1062), .B1(new_n1078), .B2(new_n1076), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1061), .B1(new_n1077), .B2(new_n1079), .ZN(G378));
  NAND3_X1  g0880(.A1(new_n842), .A2(new_n847), .A3(G330), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n296), .A2(new_n301), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n265), .A2(new_n823), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  OR3_X1    g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1085), .B2(new_n1084), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1081), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1092), .A2(new_n842), .A3(G330), .A4(new_n847), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n863), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n863), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n912), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1090), .A2(new_n712), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n698), .B1(G50), .B2(new_n1040), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n732), .A2(new_n321), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT120), .Z(new_n1103));
  OAI22_X1  g0903(.A1(new_n740), .A2(new_n438), .B1(new_n742), .B2(new_n356), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n720), .A2(new_n487), .B1(new_n728), .B2(new_n731), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n272), .A2(new_n284), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n931), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n790), .A2(G97), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1103), .A2(new_n958), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT58), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1106), .B(new_n255), .C1(G33), .C2(G41), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT119), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n742), .A2(new_n925), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n740), .A2(new_n1051), .B1(new_n720), .B2(new_n1049), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(G150), .C2(new_n746), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1117), .B1(new_n798), .B2(new_n737), .C1(new_n723), .C2(new_n1057), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n776), .A2(new_n785), .ZN(new_n1120));
  AOI211_X1 g0920(.A(G33), .B(G41), .C1(new_n729), .C2(G124), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1114), .B1(new_n1110), .B2(new_n1109), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1101), .B1(new_n1124), .B2(new_n711), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1100), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1099), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1076), .A2(new_n1072), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1098), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT57), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n665), .B1(new_n1132), .B2(new_n1128), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1127), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(KEYINPUT121), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(G375));
  NOR2_X1   g0938(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1139), .A2(new_n1075), .A3(new_n892), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT122), .Z(new_n1141));
  INV_X1    g0941(.A(new_n1069), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT123), .B1(new_n1142), .B2(new_n1033), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT123), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1069), .A2(new_n1144), .A3(new_n912), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n698), .B1(G68), .B2(new_n1040), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n720), .A2(new_n731), .B1(new_n728), .B2(new_n724), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n272), .B1(new_n745), .B2(new_n356), .C1(new_n740), .C2(new_n527), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(G107), .C2(new_n786), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n790), .A2(G116), .B1(G77), .B2(new_n776), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n430), .C2(new_n723), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n308), .B1(new_n740), .B2(new_n798), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n720), .A2(new_n925), .B1(new_n728), .B2(new_n1049), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(G159), .C2(new_n751), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n742), .A2(new_n929), .B1(new_n745), .B2(new_n255), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT124), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(new_n737), .C2(new_n1057), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1103), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1151), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1146), .B1(new_n1159), .B2(new_n711), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n820), .B2(new_n713), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1143), .A2(new_n1145), .A3(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1141), .A2(new_n1162), .ZN(G381));
  OR3_X1    g0963(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1078), .A2(new_n1076), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1061), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1137), .A3(new_n1168), .ZN(G407));
  NAND2_X1  g0969(.A1(new_n649), .A2(G213), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1137), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(G407), .A2(G213), .A3(new_n1172), .ZN(G409));
  NOR2_X1   g0973(.A1(new_n1129), .A2(new_n892), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1099), .A2(KEYINPUT126), .A3(new_n1126), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT126), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1033), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1126), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1168), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT125), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1134), .A2(G378), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1134), .B2(G378), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1181), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1139), .B1(KEYINPUT60), .B2(new_n1073), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1071), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n666), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OR3_X1    g0989(.A1(new_n1189), .A2(new_n803), .A3(new_n1162), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n803), .B1(new_n1189), .B2(new_n1162), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1185), .A2(new_n1170), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT62), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT61), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1171), .A2(G2897), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1192), .B(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1134), .A2(G378), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT125), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1134), .A2(G378), .A3(new_n1182), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1180), .A2(new_n1174), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1200), .A2(new_n1201), .B1(new_n1168), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1198), .B1(new_n1203), .B2(new_n1171), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT62), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1185), .A2(new_n1205), .A3(new_n1193), .A4(new_n1170), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1195), .A2(new_n1196), .A3(new_n1204), .A4(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(G393), .B(G396), .Z(new_n1208));
  NAND2_X1  g1008(.A1(G390), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1208), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n978), .A3(new_n1000), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1212), .A2(G387), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(G387), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1207), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1185), .A2(new_n1170), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1198), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT63), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1194), .A2(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1185), .A2(KEYINPUT63), .A3(new_n1193), .A4(new_n1170), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1215), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1217), .A2(new_n1223), .ZN(G405));
  NAND2_X1  g1024(.A1(G375), .A2(new_n1168), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1225), .A2(KEYINPUT127), .A3(new_n1193), .A4(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1137), .B2(new_n1167), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1193), .A2(KEYINPUT127), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1193), .A2(KEYINPUT127), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1227), .A2(new_n1215), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1215), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(G402));
endmodule


