

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U547 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U548 ( .A1(n511), .A2(n510), .ZN(n802) );
  XOR2_X1 U549 ( .A(KEYINPUT1), .B(n524), .Z(n653) );
  OR2_X1 U550 ( .A1(n764), .A2(n763), .ZN(n510) );
  AND2_X1 U551 ( .A1(n761), .A2(n760), .ZN(n511) );
  AND2_X1 U552 ( .A1(n900), .A2(n812), .ZN(n512) );
  NOR2_X1 U553 ( .A1(n801), .A2(n512), .ZN(n513) );
  INV_X1 U554 ( .A(KEYINPUT31), .ZN(n724) );
  AND2_X1 U555 ( .A1(G160), .A2(n687), .ZN(n712) );
  INV_X1 U556 ( .A(n712), .ZN(n728) );
  NAND2_X1 U557 ( .A1(G8), .A2(n728), .ZN(n764) );
  AND2_X1 U558 ( .A1(n519), .A2(G2105), .ZN(n967) );
  NOR2_X1 U559 ( .A1(G2105), .A2(n519), .ZN(n959) );
  XOR2_X1 U560 ( .A(KEYINPUT17), .B(n518), .Z(n960) );
  NOR2_X1 U561 ( .A1(G651), .A2(n637), .ZN(n657) );
  NOR2_X1 U562 ( .A1(n523), .A2(n522), .ZN(G164) );
  AND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n966) );
  NAND2_X1 U564 ( .A1(G114), .A2(n966), .ZN(n514) );
  XNOR2_X1 U565 ( .A(n514), .B(KEYINPUT92), .ZN(n517) );
  INV_X1 U566 ( .A(G2104), .ZN(n519) );
  NAND2_X1 U567 ( .A1(G126), .A2(n967), .ZN(n515) );
  XOR2_X1 U568 ( .A(KEYINPUT91), .B(n515), .Z(n516) );
  NAND2_X1 U569 ( .A1(n517), .A2(n516), .ZN(n523) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  NAND2_X1 U571 ( .A1(G138), .A2(n960), .ZN(n521) );
  NAND2_X1 U572 ( .A1(G102), .A2(n959), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U574 ( .A(G651), .B(KEYINPUT66), .Z(n531) );
  NOR2_X1 U575 ( .A1(G543), .A2(n531), .ZN(n524) );
  NAND2_X1 U576 ( .A1(G63), .A2(n653), .ZN(n525) );
  XNOR2_X1 U577 ( .A(KEYINPUT79), .B(n525), .ZN(n528) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n637) );
  NAND2_X1 U579 ( .A1(n657), .A2(G51), .ZN(n526) );
  XOR2_X1 U580 ( .A(KEYINPUT80), .B(n526), .Z(n527) );
  NOR2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U582 ( .A(n529), .B(KEYINPUT6), .ZN(n536) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U584 ( .A1(n649), .A2(G89), .ZN(n530) );
  XNOR2_X1 U585 ( .A(n530), .B(KEYINPUT4), .ZN(n533) );
  NOR2_X1 U586 ( .A1(n637), .A2(n531), .ZN(n650) );
  NAND2_X1 U587 ( .A1(G76), .A2(n650), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(KEYINPUT5), .B(n534), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n537), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U592 ( .A1(G125), .A2(n967), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT64), .B(n538), .Z(n541) );
  NAND2_X1 U594 ( .A1(G101), .A2(n959), .ZN(n539) );
  XNOR2_X1 U595 ( .A(KEYINPUT23), .B(n539), .ZN(n540) );
  NOR2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n966), .A2(G113), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n547) );
  INV_X1 U599 ( .A(KEYINPUT65), .ZN(n545) );
  AND2_X1 U600 ( .A1(G137), .A2(n960), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n545), .B(n544), .ZN(n546) );
  NOR2_X2 U602 ( .A1(n547), .A2(n546), .ZN(G160) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U604 ( .A(G2443), .B(G2446), .Z(n549) );
  XNOR2_X1 U605 ( .A(G2427), .B(G2451), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n549), .B(n548), .ZN(n555) );
  XOR2_X1 U607 ( .A(G2430), .B(G2454), .Z(n551) );
  XNOR2_X1 U608 ( .A(G1341), .B(G1348), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U610 ( .A(G2435), .B(G2438), .Z(n552) );
  XNOR2_X1 U611 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U612 ( .A(n555), .B(n554), .Z(n556) );
  AND2_X1 U613 ( .A1(G14), .A2(n556), .ZN(G401) );
  NAND2_X1 U614 ( .A1(n653), .A2(G64), .ZN(n557) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(n557), .Z(n564) );
  NAND2_X1 U616 ( .A1(G90), .A2(n649), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G77), .A2(n650), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT9), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G52), .A2(n657), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U622 ( .A1(n564), .A2(n563), .ZN(G171) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  INV_X1 U624 ( .A(G69), .ZN(G235) );
  INV_X1 U625 ( .A(G108), .ZN(G238) );
  INV_X1 U626 ( .A(G120), .ZN(G236) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  NAND2_X1 U628 ( .A1(G94), .A2(G452), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT69), .ZN(G173) );
  XOR2_X1 U630 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n567) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G223) );
  XOR2_X1 U633 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n569) );
  INV_X1 U634 ( .A(G223), .ZN(n817) );
  NAND2_X1 U635 ( .A1(G567), .A2(n817), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G234) );
  XOR2_X1 U637 ( .A(G860), .B(KEYINPUT76), .Z(n600) );
  NAND2_X1 U638 ( .A1(n649), .A2(G81), .ZN(n570) );
  XNOR2_X1 U639 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G68), .A2(n650), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(n573), .Z(n577) );
  NAND2_X1 U643 ( .A1(n653), .A2(G56), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT75), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT14), .ZN(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n657), .A2(G43), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n882) );
  OR2_X1 U649 ( .A1(n600), .A2(n882), .ZN(G153) );
  NAND2_X1 U650 ( .A1(G66), .A2(n653), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G92), .A2(n649), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G54), .A2(n657), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G79), .A2(n650), .ZN(n582) );
  XNOR2_X1 U655 ( .A(KEYINPUT77), .B(n582), .ZN(n583) );
  NOR2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U658 ( .A(KEYINPUT15), .B(n587), .Z(n992) );
  INV_X1 U659 ( .A(G868), .ZN(n668) );
  NAND2_X1 U660 ( .A1(n992), .A2(n668), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n588), .B(KEYINPUT78), .ZN(n590) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G91), .A2(n649), .ZN(n592) );
  NAND2_X1 U665 ( .A1(G53), .A2(n657), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n650), .A2(G78), .ZN(n593) );
  XOR2_X1 U668 ( .A(KEYINPUT70), .B(n593), .Z(n594) );
  NOR2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G65), .A2(n653), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n668), .ZN(n599) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U674 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n600), .A2(G559), .ZN(n601) );
  INV_X1 U676 ( .A(n992), .ZN(n617) );
  NAND2_X1 U677 ( .A1(n601), .A2(n617), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n882), .ZN(n603) );
  XOR2_X1 U680 ( .A(KEYINPUT81), .B(n603), .Z(n606) );
  NAND2_X1 U681 ( .A1(G868), .A2(n617), .ZN(n604) );
  NOR2_X1 U682 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G99), .A2(n959), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G111), .A2(n966), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G135), .A2(n960), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n967), .A2(G123), .ZN(n609) );
  XOR2_X1 U689 ( .A(KEYINPUT18), .B(n609), .Z(n610) );
  NOR2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT82), .ZN(n972) );
  XOR2_X1 U693 ( .A(n972), .B(G2096), .Z(n616) );
  XNOR2_X1 U694 ( .A(G2100), .B(KEYINPUT83), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G559), .A2(n617), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n618), .B(KEYINPUT84), .ZN(n666) );
  XNOR2_X1 U698 ( .A(n666), .B(n882), .ZN(n619) );
  NOR2_X1 U699 ( .A1(n619), .A2(G860), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G93), .A2(n649), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G80), .A2(n650), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n657), .A2(G55), .ZN(n623) );
  NAND2_X1 U704 ( .A1(G67), .A2(n653), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U706 ( .A(KEYINPUT85), .B(n624), .Z(n625) );
  OR2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n669) );
  XOR2_X1 U708 ( .A(n627), .B(n669), .Z(G145) );
  NAND2_X1 U709 ( .A1(G86), .A2(n649), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G48), .A2(n657), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n650), .A2(G73), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n630), .B(KEYINPUT2), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n631), .B(KEYINPUT87), .ZN(n632) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G61), .A2(n653), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n636) );
  XNOR2_X1 U719 ( .A(n636), .B(KEYINPUT86), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G49), .A2(n657), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G87), .A2(n637), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U723 ( .A1(n653), .A2(n640), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U725 ( .A1(G88), .A2(n649), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G75), .A2(n650), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n657), .A2(G50), .ZN(n646) );
  NAND2_X1 U729 ( .A1(G62), .A2(n653), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U731 ( .A1(n648), .A2(n647), .ZN(G166) );
  NAND2_X1 U732 ( .A1(G85), .A2(n649), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G72), .A2(n650), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U735 ( .A1(G60), .A2(n653), .ZN(n654) );
  XNOR2_X1 U736 ( .A(KEYINPUT67), .B(n654), .ZN(n655) );
  NOR2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n657), .A2(G47), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(G290) );
  XOR2_X1 U740 ( .A(n669), .B(n882), .Z(n665) );
  XNOR2_X1 U741 ( .A(G288), .B(KEYINPUT19), .ZN(n661) );
  INV_X1 U742 ( .A(G299), .ZN(n694) );
  XNOR2_X1 U743 ( .A(G166), .B(n694), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U745 ( .A(n662), .B(G290), .Z(n663) );
  XNOR2_X1 U746 ( .A(G305), .B(n663), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n665), .B(n664), .ZN(n994) );
  XOR2_X1 U748 ( .A(n994), .B(n666), .Z(n667) );
  NOR2_X1 U749 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U750 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U751 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U758 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  XNOR2_X1 U759 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n677) );
  XNOR2_X1 U761 ( .A(KEYINPUT88), .B(KEYINPUT22), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n678), .A2(G96), .ZN(n679) );
  NOR2_X1 U764 ( .A1(G218), .A2(n679), .ZN(n680) );
  XNOR2_X1 U765 ( .A(KEYINPUT89), .B(n680), .ZN(n821) );
  NAND2_X1 U766 ( .A1(n821), .A2(G2106), .ZN(n685) );
  NOR2_X1 U767 ( .A1(G237), .A2(G236), .ZN(n682) );
  NOR2_X1 U768 ( .A1(G238), .A2(G235), .ZN(n681) );
  NAND2_X1 U769 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U770 ( .A(KEYINPUT90), .B(n683), .ZN(n822) );
  NAND2_X1 U771 ( .A1(G567), .A2(n822), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n938) );
  NAND2_X1 U773 ( .A1(G661), .A2(G483), .ZN(n686) );
  NOR2_X1 U774 ( .A1(n938), .A2(n686), .ZN(n820) );
  NAND2_X1 U775 ( .A1(n820), .A2(G36), .ZN(G176) );
  INV_X1 U776 ( .A(G166), .ZN(G303) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n766) );
  AND2_X1 U778 ( .A1(G40), .A2(n766), .ZN(n687) );
  NOR2_X1 U779 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NAND2_X1 U780 ( .A1(n749), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U781 ( .A1(n764), .A2(n688), .ZN(n754) );
  NAND2_X1 U782 ( .A1(n712), .A2(G2072), .ZN(n689) );
  XNOR2_X1 U783 ( .A(n689), .B(KEYINPUT27), .ZN(n691) );
  AND2_X1 U784 ( .A1(G1956), .A2(n728), .ZN(n690) );
  NOR2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n693) );
  XOR2_X1 U787 ( .A(KEYINPUT102), .B(KEYINPUT28), .Z(n692) );
  XNOR2_X1 U788 ( .A(n693), .B(n692), .ZN(n710) );
  NAND2_X1 U789 ( .A1(n695), .A2(n694), .ZN(n708) );
  AND2_X1 U790 ( .A1(n712), .A2(G1996), .ZN(n696) );
  XOR2_X1 U791 ( .A(n696), .B(KEYINPUT26), .Z(n698) );
  NAND2_X1 U792 ( .A1(n728), .A2(G1341), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U794 ( .A1(n882), .A2(n699), .ZN(n703) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n728), .ZN(n701) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n712), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n992), .A2(n704), .ZN(n702) );
  OR2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n992), .A2(n704), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U804 ( .A(n711), .B(KEYINPUT29), .Z(n717) );
  XOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .Z(n865) );
  NOR2_X1 U806 ( .A1(n865), .A2(n728), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n712), .A2(G1961), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U809 ( .A(KEYINPUT101), .B(n715), .ZN(n721) );
  NAND2_X1 U810 ( .A1(G171), .A2(n721), .ZN(n716) );
  NAND2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n727) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n764), .ZN(n742) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n728), .ZN(n739) );
  NOR2_X1 U814 ( .A1(n742), .A2(n739), .ZN(n718) );
  NAND2_X1 U815 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U816 ( .A(n719), .B(KEYINPUT30), .ZN(n720) );
  NOR2_X1 U817 ( .A1(n720), .A2(G168), .ZN(n723) );
  NOR2_X1 U818 ( .A1(G171), .A2(n721), .ZN(n722) );
  XNOR2_X1 U819 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n740) );
  NAND2_X1 U821 ( .A1(n740), .A2(G286), .ZN(n735) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n764), .ZN(n730) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U825 ( .A(KEYINPUT103), .B(n731), .Z(n732) );
  NAND2_X1 U826 ( .A1(n732), .A2(G303), .ZN(n733) );
  XNOR2_X1 U827 ( .A(n733), .B(KEYINPUT104), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n736), .A2(G8), .ZN(n738) );
  XOR2_X1 U830 ( .A(KEYINPUT32), .B(KEYINPUT105), .Z(n737) );
  XNOR2_X1 U831 ( .A(n738), .B(n737), .ZN(n746) );
  NAND2_X1 U832 ( .A1(G8), .A2(n739), .ZN(n744) );
  INV_X1 U833 ( .A(n740), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U837 ( .A(n747), .B(KEYINPUT106), .ZN(n757) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n894) );
  NAND2_X1 U840 ( .A1(n757), .A2(n894), .ZN(n750) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n890) );
  NAND2_X1 U842 ( .A1(n750), .A2(n890), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n751), .A2(n764), .ZN(n752) );
  NOR2_X1 U844 ( .A1(KEYINPUT33), .A2(n752), .ZN(n753) );
  NOR2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n886) );
  NAND2_X1 U847 ( .A1(n755), .A2(n886), .ZN(n761) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n756) );
  NAND2_X1 U849 ( .A1(G8), .A2(n756), .ZN(n758) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n759), .A2(n764), .ZN(n760) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U853 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  NAND2_X1 U854 ( .A1(G160), .A2(G40), .ZN(n765) );
  NOR2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n812) );
  NAND2_X1 U856 ( .A1(n959), .A2(G104), .ZN(n767) );
  XNOR2_X1 U857 ( .A(n767), .B(KEYINPUT94), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G140), .A2(n960), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n770), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G116), .A2(n966), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G128), .A2(n967), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n773), .Z(n774) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U866 ( .A(KEYINPUT36), .B(n776), .Z(n988) );
  XOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .Z(n803) );
  NAND2_X1 U868 ( .A1(n988), .A2(n803), .ZN(n777) );
  XNOR2_X1 U869 ( .A(KEYINPUT95), .B(n777), .ZN(n855) );
  NAND2_X1 U870 ( .A1(n812), .A2(n855), .ZN(n809) );
  NAND2_X1 U871 ( .A1(n967), .A2(G119), .ZN(n778) );
  XNOR2_X1 U872 ( .A(n778), .B(KEYINPUT96), .ZN(n780) );
  NAND2_X1 U873 ( .A1(G107), .A2(n966), .ZN(n779) );
  NAND2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U875 ( .A(KEYINPUT97), .B(n781), .ZN(n785) );
  NAND2_X1 U876 ( .A1(G131), .A2(n960), .ZN(n783) );
  NAND2_X1 U877 ( .A1(G95), .A2(n959), .ZN(n782) );
  AND2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n985) );
  AND2_X1 U880 ( .A1(n985), .A2(G1991), .ZN(n797) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(KEYINPUT100), .Z(n787) );
  NAND2_X1 U882 ( .A1(G105), .A2(n959), .ZN(n786) );
  XNOR2_X1 U883 ( .A(n787), .B(n786), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n967), .A2(G129), .ZN(n788) );
  XNOR2_X1 U885 ( .A(n788), .B(KEYINPUT98), .ZN(n790) );
  NAND2_X1 U886 ( .A1(G117), .A2(n966), .ZN(n789) );
  NAND2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U888 ( .A(KEYINPUT99), .B(n791), .Z(n792) );
  NOR2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n960), .A2(G141), .ZN(n794) );
  NAND2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n987) );
  AND2_X1 U892 ( .A1(n987), .A2(G1996), .ZN(n796) );
  NOR2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n849) );
  INV_X1 U894 ( .A(n812), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n849), .A2(n798), .ZN(n806) );
  INV_X1 U896 ( .A(n806), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n809), .A2(n799), .ZN(n801) );
  XOR2_X1 U898 ( .A(G1986), .B(KEYINPUT93), .Z(n800) );
  XNOR2_X1 U899 ( .A(G290), .B(n800), .ZN(n900) );
  NAND2_X1 U900 ( .A1(n802), .A2(n513), .ZN(n815) );
  OR2_X1 U901 ( .A1(n988), .A2(n803), .ZN(n843) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n987), .ZN(n831) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n985), .ZN(n847) );
  NOR2_X1 U905 ( .A1(n804), .A2(n847), .ZN(n805) );
  NOR2_X1 U906 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n831), .A2(n807), .ZN(n808) );
  XNOR2_X1 U908 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U910 ( .A1(n843), .A2(n811), .ZN(n813) );
  NAND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U913 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U916 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(G188) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(G325) );
  XNOR2_X1 U920 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  NAND2_X1 U922 ( .A1(G124), .A2(n967), .ZN(n823) );
  XNOR2_X1 U923 ( .A(n823), .B(KEYINPUT44), .ZN(n825) );
  NAND2_X1 U924 ( .A1(n966), .A2(G112), .ZN(n824) );
  NAND2_X1 U925 ( .A1(n825), .A2(n824), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G136), .A2(n960), .ZN(n827) );
  NAND2_X1 U927 ( .A1(G100), .A2(n959), .ZN(n826) );
  NAND2_X1 U928 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U929 ( .A1(n829), .A2(n828), .ZN(G162) );
  XOR2_X1 U930 ( .A(G2090), .B(G162), .Z(n830) );
  NOR2_X1 U931 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U932 ( .A(KEYINPUT51), .B(n832), .Z(n853) );
  NAND2_X1 U933 ( .A1(G139), .A2(n960), .ZN(n834) );
  NAND2_X1 U934 ( .A1(G103), .A2(n959), .ZN(n833) );
  NAND2_X1 U935 ( .A1(n834), .A2(n833), .ZN(n839) );
  NAND2_X1 U936 ( .A1(G115), .A2(n966), .ZN(n836) );
  NAND2_X1 U937 ( .A1(G127), .A2(n967), .ZN(n835) );
  NAND2_X1 U938 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(KEYINPUT47), .B(n837), .Z(n838) );
  NOR2_X1 U940 ( .A1(n839), .A2(n838), .ZN(n978) );
  XOR2_X1 U941 ( .A(G2072), .B(n978), .Z(n841) );
  XOR2_X1 U942 ( .A(G164), .B(G2078), .Z(n840) );
  NOR2_X1 U943 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n842), .B(KEYINPUT50), .ZN(n844) );
  NAND2_X1 U945 ( .A1(n844), .A2(n843), .ZN(n851) );
  XNOR2_X1 U946 ( .A(G160), .B(G2084), .ZN(n845) );
  NAND2_X1 U947 ( .A1(n845), .A2(n972), .ZN(n846) );
  NOR2_X1 U948 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U950 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U953 ( .A(KEYINPUT52), .B(n856), .ZN(n857) );
  INV_X1 U954 ( .A(KEYINPUT55), .ZN(n878) );
  NAND2_X1 U955 ( .A1(n857), .A2(n878), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n858), .A2(G29), .ZN(n909) );
  XNOR2_X1 U957 ( .A(G2090), .B(G35), .ZN(n873) );
  XOR2_X1 U958 ( .A(G1991), .B(G25), .Z(n859) );
  NAND2_X1 U959 ( .A1(n859), .A2(G28), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT119), .ZN(n864) );
  XNOR2_X1 U961 ( .A(G2067), .B(G26), .ZN(n862) );
  XNOR2_X1 U962 ( .A(G33), .B(G2072), .ZN(n861) );
  NOR2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n870) );
  XNOR2_X1 U965 ( .A(G1996), .B(G32), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n865), .B(G27), .ZN(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(KEYINPUT120), .B(n868), .Z(n869) );
  NOR2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U970 ( .A(KEYINPUT53), .B(n871), .ZN(n872) );
  NOR2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n876) );
  XOR2_X1 U972 ( .A(G2084), .B(G34), .Z(n874) );
  XNOR2_X1 U973 ( .A(KEYINPUT54), .B(n874), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n880) );
  INV_X1 U976 ( .A(G29), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G11), .A2(n881), .ZN(n907) );
  XNOR2_X1 U979 ( .A(G301), .B(G1961), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n882), .B(G1341), .ZN(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n902) );
  XOR2_X1 U982 ( .A(G1966), .B(G168), .Z(n885) );
  XNOR2_X1 U983 ( .A(KEYINPUT121), .B(n885), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n888), .B(KEYINPUT57), .ZN(n898) );
  NAND2_X1 U986 ( .A1(G1971), .A2(G303), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n896) );
  XNOR2_X1 U988 ( .A(G299), .B(G1956), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n992), .B(G1348), .ZN(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  NOR2_X1 U994 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U995 ( .A1(n902), .A2(n901), .ZN(n904) );
  XNOR2_X1 U996 ( .A(KEYINPUT56), .B(G16), .ZN(n903) );
  NAND2_X1 U997 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U998 ( .A(KEYINPUT122), .B(n905), .Z(n906) );
  NOR2_X1 U999 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1000 ( .A1(n909), .A2(n908), .ZN(n936) );
  XNOR2_X1 U1001 ( .A(G1961), .B(G5), .ZN(n910) );
  XNOR2_X1 U1002 ( .A(n910), .B(KEYINPUT123), .ZN(n918) );
  XOR2_X1 U1003 ( .A(G1986), .B(KEYINPUT126), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G24), .B(n911), .ZN(n915) );
  XNOR2_X1 U1005 ( .A(G1971), .B(G22), .ZN(n913) );
  XNOR2_X1 U1006 ( .A(G23), .B(G1976), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1009 ( .A(KEYINPUT58), .B(n916), .Z(n917) );
  NAND2_X1 U1010 ( .A1(n918), .A2(n917), .ZN(n932) );
  XNOR2_X1 U1011 ( .A(G1966), .B(G21), .ZN(n929) );
  XOR2_X1 U1012 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n927) );
  XOR2_X1 U1013 ( .A(G20), .B(G1956), .Z(n922) );
  XNOR2_X1 U1014 ( .A(G1341), .B(G19), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(G1981), .B(G6), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n925) );
  XOR2_X1 U1018 ( .A(KEYINPUT59), .B(G1348), .Z(n923) );
  XNOR2_X1 U1019 ( .A(G4), .B(n923), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1022 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1023 ( .A(n930), .B(KEYINPUT125), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1025 ( .A(KEYINPUT61), .B(n933), .Z(n934) );
  NOR2_X1 U1026 ( .A1(G16), .A2(n934), .ZN(n935) );
  NOR2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1028 ( .A(n937), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1029 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1030 ( .A(G96), .ZN(G221) );
  INV_X1 U1031 ( .A(n938), .ZN(G319) );
  XOR2_X1 U1032 ( .A(KEYINPUT41), .B(G2474), .Z(n940) );
  XNOR2_X1 U1033 ( .A(G1986), .B(G1976), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n940), .B(n939), .ZN(n941) );
  XOR2_X1 U1035 ( .A(n941), .B(KEYINPUT110), .Z(n943) );
  XNOR2_X1 U1036 ( .A(G1996), .B(G1956), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n943), .B(n942), .ZN(n947) );
  XOR2_X1 U1038 ( .A(KEYINPUT109), .B(G1971), .Z(n945) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G1961), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n945), .B(n944), .ZN(n946) );
  XOR2_X1 U1041 ( .A(n947), .B(n946), .Z(n949) );
  XNOR2_X1 U1042 ( .A(G1991), .B(G1981), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n949), .B(n948), .ZN(G229) );
  XOR2_X1 U1044 ( .A(G2100), .B(G2096), .Z(n951) );
  XNOR2_X1 U1045 ( .A(G2090), .B(KEYINPUT43), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(n951), .B(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(n952), .B(G2678), .Z(n954) );
  XNOR2_X1 U1048 ( .A(G2072), .B(KEYINPUT108), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n954), .B(n953), .ZN(n958) );
  XOR2_X1 U1050 ( .A(KEYINPUT42), .B(G2084), .Z(n956) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G2078), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(n956), .B(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n958), .B(n957), .ZN(G227) );
  XNOR2_X1 U1054 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n965) );
  NAND2_X1 U1055 ( .A1(n959), .A2(G106), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n960), .A2(G142), .ZN(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT111), .B(n961), .Z(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1059 ( .A(n965), .B(n964), .Z(n971) );
  NAND2_X1 U1060 ( .A1(G118), .A2(n966), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(G130), .A2(n967), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n972), .B(G160), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n974), .B(n973), .ZN(n982) );
  XOR2_X1 U1066 ( .A(KEYINPUT114), .B(KEYINPUT116), .Z(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(n977), .B(KEYINPUT46), .Z(n980) );
  XNOR2_X1 U1070 ( .A(n978), .B(KEYINPUT115), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n980), .B(n979), .ZN(n981) );
  XOR2_X1 U1072 ( .A(n982), .B(n981), .Z(n984) );
  XNOR2_X1 U1073 ( .A(G164), .B(G162), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n984), .B(n983), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n986), .B(n985), .ZN(n990) );
  XOR2_X1 U1076 ( .A(n988), .B(n987), .Z(n989) );
  XNOR2_X1 U1077 ( .A(n990), .B(n989), .ZN(n991) );
  NOR2_X1 U1078 ( .A1(G37), .A2(n991), .ZN(G395) );
  XNOR2_X1 U1079 ( .A(G286), .B(G301), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(n993), .B(n992), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(n995), .B(n994), .ZN(n996) );
  NOR2_X1 U1082 ( .A1(G37), .A2(n996), .ZN(G397) );
  NOR2_X1 U1083 ( .A1(G229), .A2(G227), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(n997), .B(KEYINPUT49), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(G401), .A2(n998), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(G319), .A2(n999), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT117), .B(n1000), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(G395), .A2(G397), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(KEYINPUT118), .B(n1003), .Z(G308) );
  INV_X1 U1091 ( .A(G308), .ZN(G225) );
endmodule

