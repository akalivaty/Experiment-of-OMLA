

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U551 ( .A1(n687), .A2(n686), .ZN(n704) );
  BUF_X2 U552 ( .A(n649), .Z(n650) );
  NOR2_X2 U553 ( .A1(n584), .A2(n536), .ZN(n788) );
  XNOR2_X2 U554 ( .A(n594), .B(KEYINPUT83), .ZN(n705) );
  NOR2_X1 U555 ( .A1(n649), .A2(n595), .ZN(n597) );
  NOR2_X1 U556 ( .A1(n604), .A2(n603), .ZN(n607) );
  AND2_X1 U557 ( .A1(n518), .A2(G2104), .ZN(n545) );
  XNOR2_X1 U558 ( .A(n519), .B(KEYINPUT64), .ZN(n520) );
  INV_X1 U559 ( .A(KEYINPUT23), .ZN(n519) );
  AND2_X2 U560 ( .A1(n522), .A2(G2105), .ZN(n886) );
  BUF_X1 U561 ( .A(n545), .Z(n889) );
  AND2_X1 U562 ( .A1(n744), .A2(n966), .ZN(n516) );
  XOR2_X1 U563 ( .A(n607), .B(n606), .Z(n517) );
  INV_X1 U564 ( .A(KEYINPUT26), .ZN(n596) );
  INV_X1 U565 ( .A(KEYINPUT94), .ZN(n620) );
  NOR2_X1 U566 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U567 ( .A1(n705), .A2(n707), .ZN(n649) );
  AND2_X1 U568 ( .A1(n677), .A2(n676), .ZN(n678) );
  INV_X1 U569 ( .A(KEYINPUT13), .ZN(n605) );
  XNOR2_X1 U570 ( .A(n605), .B(KEYINPUT72), .ZN(n606) );
  INV_X1 U571 ( .A(G2105), .ZN(n518) );
  NOR2_X1 U572 ( .A1(n739), .A2(n516), .ZN(n740) );
  INV_X1 U573 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n741), .A2(n740), .ZN(n743) );
  NOR2_X2 U575 ( .A1(G651), .A2(G543), .ZN(n787) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n584) );
  XNOR2_X1 U577 ( .A(n526), .B(n525), .ZN(n531) );
  NOR2_X2 U578 ( .A1(n531), .A2(n530), .ZN(G160) );
  NAND2_X1 U579 ( .A1(G101), .A2(n545), .ZN(n521) );
  XNOR2_X1 U580 ( .A(n521), .B(n520), .ZN(n524) );
  NAND2_X1 U581 ( .A1(G125), .A2(n886), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n526) );
  INV_X1 U583 ( .A(KEYINPUT65), .ZN(n525) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U585 ( .A1(G113), .A2(n885), .ZN(n529) );
  NOR2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X1 U587 ( .A(KEYINPUT17), .B(n527), .Z(n710) );
  NAND2_X1 U588 ( .A1(G137), .A2(n710), .ZN(n528) );
  NAND2_X1 U589 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n787), .A2(G89), .ZN(n532) );
  XNOR2_X1 U591 ( .A(n532), .B(KEYINPUT4), .ZN(n534) );
  INV_X1 U592 ( .A(G651), .ZN(n536) );
  NAND2_X1 U593 ( .A1(G76), .A2(n788), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U595 ( .A(n535), .B(KEYINPUT5), .ZN(n543) );
  NOR2_X1 U596 ( .A1(G543), .A2(n536), .ZN(n538) );
  XNOR2_X1 U597 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n537) );
  XNOR2_X1 U598 ( .A(n538), .B(n537), .ZN(n791) );
  NAND2_X1 U599 ( .A1(G63), .A2(n791), .ZN(n540) );
  NOR2_X2 U600 ( .A1(G651), .A2(n584), .ZN(n793) );
  NAND2_X1 U601 ( .A1(G51), .A2(n793), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(n541), .Z(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U605 ( .A(n544), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U606 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U607 ( .A1(G102), .A2(n889), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G138), .A2(n710), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G114), .A2(n885), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G126), .A2(n886), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n551), .A2(n550), .ZN(G164) );
  NAND2_X1 U614 ( .A1(G91), .A2(n787), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G53), .A2(n793), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G65), .A2(n791), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G78), .A2(n788), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n558), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U622 ( .A1(G64), .A2(n791), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G52), .A2(n793), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U625 ( .A1(G90), .A2(n787), .ZN(n562) );
  NAND2_X1 U626 ( .A1(G77), .A2(n788), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT68), .B(n566), .ZN(G171) );
  NAND2_X1 U631 ( .A1(G88), .A2(n787), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G75), .A2(n788), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G62), .A2(n791), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G50), .A2(n793), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(G166) );
  INV_X1 U638 ( .A(G166), .ZN(G303) );
  NAND2_X1 U639 ( .A1(G86), .A2(n787), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G61), .A2(n791), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n788), .A2(G73), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n575), .Z(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n793), .A2(G48), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(G305) );
  NAND2_X1 U647 ( .A1(G49), .A2(n793), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G74), .A2(G651), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n791), .A2(n582), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT79), .B(n583), .Z(n586) );
  NAND2_X1 U652 ( .A1(n584), .A2(G87), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U654 ( .A1(n793), .A2(G47), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n791), .A2(G60), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G85), .A2(n787), .ZN(n589) );
  XOR2_X1 U658 ( .A(KEYINPUT66), .B(n589), .Z(n590) );
  NOR2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n788), .A2(G72), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G290) );
  NAND2_X1 U662 ( .A1(G160), .A2(G40), .ZN(n594) );
  NOR2_X1 U663 ( .A1(G164), .A2(G1384), .ZN(n707) );
  INV_X1 U664 ( .A(G1996), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n597), .B(n596), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n650), .A2(G1341), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n611) );
  NAND2_X1 U668 ( .A1(n791), .A2(G56), .ZN(n600) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n600), .Z(n608) );
  NAND2_X1 U670 ( .A1(n788), .A2(G68), .ZN(n601) );
  XNOR2_X1 U671 ( .A(KEYINPUT71), .B(n601), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n787), .A2(G81), .ZN(n602) );
  XOR2_X1 U673 ( .A(n602), .B(KEYINPUT12), .Z(n603) );
  NOR2_X1 U674 ( .A1(n608), .A2(n517), .ZN(n610) );
  NAND2_X1 U675 ( .A1(n793), .A2(G43), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n610), .A2(n609), .ZN(n972) );
  NOR2_X2 U677 ( .A1(n611), .A2(n972), .ZN(n622) );
  NAND2_X1 U678 ( .A1(G79), .A2(n788), .ZN(n613) );
  NAND2_X1 U679 ( .A1(G54), .A2(n793), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U681 ( .A(KEYINPUT74), .B(n614), .ZN(n618) );
  NAND2_X1 U682 ( .A1(G92), .A2(n787), .ZN(n616) );
  NAND2_X1 U683 ( .A1(G66), .A2(n791), .ZN(n615) );
  NAND2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X2 U686 ( .A(KEYINPUT15), .B(n619), .Z(n963) );
  NOR2_X1 U687 ( .A1(n622), .A2(n963), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n621), .B(n620), .ZN(n628) );
  NAND2_X1 U689 ( .A1(n622), .A2(n963), .ZN(n626) );
  NOR2_X1 U690 ( .A1(G2067), .A2(n650), .ZN(n624) );
  INV_X1 U691 ( .A(n649), .ZN(n644) );
  NOR2_X1 U692 ( .A1(n644), .A2(G1348), .ZN(n623) );
  NOR2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n628), .A2(n627), .ZN(n633) );
  INV_X1 U696 ( .A(G299), .ZN(n983) );
  NAND2_X1 U697 ( .A1(n644), .A2(G2072), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n629), .B(KEYINPUT27), .ZN(n631) );
  INV_X1 U699 ( .A(G1956), .ZN(n1000) );
  NOR2_X1 U700 ( .A1(n1000), .A2(n644), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n636) );
  NAND2_X1 U702 ( .A1(n983), .A2(n636), .ZN(n632) );
  AND2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n635) );
  INV_X1 U704 ( .A(KEYINPUT95), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n640) );
  OR2_X1 U706 ( .A1(n983), .A2(n636), .ZN(n637) );
  XNOR2_X1 U707 ( .A(KEYINPUT28), .B(n637), .ZN(n638) );
  XNOR2_X1 U708 ( .A(KEYINPUT93), .B(n638), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n641), .B(KEYINPUT29), .ZN(n648) );
  XOR2_X1 U710 ( .A(G1961), .B(KEYINPUT90), .Z(n998) );
  NAND2_X1 U711 ( .A1(n998), .A2(n650), .ZN(n642) );
  XOR2_X1 U712 ( .A(KEYINPUT91), .B(n642), .Z(n646) );
  XNOR2_X1 U713 ( .A(G2078), .B(KEYINPUT25), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(KEYINPUT92), .ZN(n944) );
  NAND2_X1 U715 ( .A1(n644), .A2(n944), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n655) );
  NAND2_X1 U717 ( .A1(n655), .A2(G171), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n648), .A2(n647), .ZN(n661) );
  NAND2_X1 U719 ( .A1(G8), .A2(n649), .ZN(n696) );
  NOR2_X1 U720 ( .A1(G1966), .A2(n696), .ZN(n675) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n650), .ZN(n671) );
  NOR2_X1 U722 ( .A1(n675), .A2(n671), .ZN(n651) );
  NAND2_X1 U723 ( .A1(G8), .A2(n651), .ZN(n652) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n652), .ZN(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT96), .B(n653), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G168), .A2(n654), .ZN(n657) );
  NOR2_X1 U727 ( .A1(n655), .A2(G171), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT31), .B(n658), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n659), .B(KEYINPUT97), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n673) );
  NAND2_X1 U732 ( .A1(n673), .A2(G286), .ZN(n666) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n696), .ZN(n663) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n650), .ZN(n662) );
  NOR2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U736 ( .A1(n664), .A2(G303), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U738 ( .A(n667), .B(KEYINPUT98), .ZN(n668) );
  AND2_X1 U739 ( .A1(n668), .A2(G8), .ZN(n670) );
  INV_X1 U740 ( .A(KEYINPUT32), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n670), .B(n669), .ZN(n677) );
  NAND2_X1 U742 ( .A1(G8), .A2(n671), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  OR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n678), .B(KEYINPUT99), .ZN(n692) );
  NAND2_X1 U746 ( .A1(G8), .A2(G166), .ZN(n679) );
  NOR2_X1 U747 ( .A1(G2090), .A2(n679), .ZN(n682) );
  NOR2_X1 U748 ( .A1(G1981), .A2(G305), .ZN(n680) );
  XOR2_X1 U749 ( .A(n680), .B(KEYINPUT24), .Z(n681) );
  NOR2_X1 U750 ( .A1(n696), .A2(n681), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n682), .A2(n684), .ZN(n683) );
  AND2_X1 U752 ( .A1(n692), .A2(n683), .ZN(n687) );
  INV_X1 U753 ( .A(n684), .ZN(n685) );
  INV_X1 U754 ( .A(n696), .ZN(n694) );
  AND2_X1 U755 ( .A1(n685), .A2(n694), .ZN(n686) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n688) );
  NOR2_X1 U758 ( .A1(n981), .A2(n688), .ZN(n690) );
  INV_X1 U759 ( .A(KEYINPUT33), .ZN(n689) );
  AND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n702) );
  XOR2_X1 U762 ( .A(G1981), .B(G305), .Z(n968) );
  NAND2_X1 U763 ( .A1(G288), .A2(G1976), .ZN(n693) );
  XNOR2_X1 U764 ( .A(n693), .B(KEYINPUT100), .ZN(n978) );
  AND2_X1 U765 ( .A1(n694), .A2(n978), .ZN(n695) );
  NOR2_X1 U766 ( .A1(KEYINPUT33), .A2(n695), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n981), .A2(KEYINPUT33), .ZN(n697) );
  NOR2_X1 U768 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U769 ( .A1(n699), .A2(n698), .ZN(n700) );
  AND2_X1 U770 ( .A1(n968), .A2(n700), .ZN(n701) );
  NAND2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n741) );
  INV_X1 U773 ( .A(n705), .ZN(n706) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n744) );
  XNOR2_X1 U775 ( .A(KEYINPUT88), .B(n744), .ZN(n727) );
  NAND2_X1 U776 ( .A1(G105), .A2(n889), .ZN(n708) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n708), .Z(n709) );
  XNOR2_X1 U778 ( .A(n709), .B(KEYINPUT85), .ZN(n712) );
  BUF_X1 U779 ( .A(n710), .Z(n890) );
  NAND2_X1 U780 ( .A1(G141), .A2(n890), .ZN(n711) );
  NAND2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U782 ( .A1(G117), .A2(n885), .ZN(n714) );
  NAND2_X1 U783 ( .A1(G129), .A2(n886), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U786 ( .A(KEYINPUT86), .B(n717), .Z(n900) );
  NAND2_X1 U787 ( .A1(G1996), .A2(n900), .ZN(n718) );
  XOR2_X1 U788 ( .A(KEYINPUT87), .B(n718), .Z(n726) );
  NAND2_X1 U789 ( .A1(G95), .A2(n889), .ZN(n720) );
  NAND2_X1 U790 ( .A1(G107), .A2(n885), .ZN(n719) );
  NAND2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U792 ( .A1(G131), .A2(n890), .ZN(n722) );
  NAND2_X1 U793 ( .A1(G119), .A2(n886), .ZN(n721) );
  NAND2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n723) );
  OR2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n879) );
  NAND2_X1 U796 ( .A1(G1991), .A2(n879), .ZN(n725) );
  NAND2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n937) );
  NAND2_X1 U798 ( .A1(n727), .A2(n937), .ZN(n728) );
  XNOR2_X1 U799 ( .A(KEYINPUT89), .B(n728), .ZN(n749) );
  XNOR2_X1 U800 ( .A(G2067), .B(KEYINPUT37), .ZN(n729) );
  XOR2_X1 U801 ( .A(n729), .B(KEYINPUT84), .Z(n745) );
  NAND2_X1 U802 ( .A1(G104), .A2(n889), .ZN(n731) );
  NAND2_X1 U803 ( .A1(G140), .A2(n890), .ZN(n730) );
  NAND2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U805 ( .A(KEYINPUT34), .B(n732), .ZN(n737) );
  NAND2_X1 U806 ( .A1(G116), .A2(n885), .ZN(n734) );
  NAND2_X1 U807 ( .A1(G128), .A2(n886), .ZN(n733) );
  NAND2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U809 ( .A(KEYINPUT35), .B(n735), .Z(n736) );
  NOR2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U811 ( .A(KEYINPUT36), .B(n738), .Z(n903) );
  AND2_X1 U812 ( .A1(n745), .A2(n903), .ZN(n918) );
  AND2_X1 U813 ( .A1(n744), .A2(n918), .ZN(n753) );
  OR2_X1 U814 ( .A1(n749), .A2(n753), .ZN(n739) );
  XNOR2_X1 U815 ( .A(G1986), .B(G290), .ZN(n966) );
  INV_X1 U816 ( .A(KEYINPUT101), .ZN(n742) );
  XNOR2_X1 U817 ( .A(n743), .B(n742), .ZN(n759) );
  INV_X1 U818 ( .A(n744), .ZN(n756) );
  NOR2_X1 U819 ( .A1(n903), .A2(n745), .ZN(n917) );
  NOR2_X1 U820 ( .A1(G1996), .A2(n900), .ZN(n920) );
  NOR2_X1 U821 ( .A1(G1991), .A2(n879), .ZN(n925) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n746) );
  XNOR2_X1 U823 ( .A(KEYINPUT102), .B(n746), .ZN(n747) );
  NOR2_X1 U824 ( .A1(n925), .A2(n747), .ZN(n748) );
  NOR2_X1 U825 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U826 ( .A1(n920), .A2(n750), .ZN(n751) );
  XOR2_X1 U827 ( .A(KEYINPUT39), .B(n751), .Z(n752) );
  NOR2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U829 ( .A1(n917), .A2(n754), .ZN(n755) );
  NOR2_X1 U830 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U831 ( .A(KEYINPUT103), .B(n757), .ZN(n758) );
  NAND2_X1 U832 ( .A1(n759), .A2(n758), .ZN(n761) );
  XNOR2_X1 U833 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n761), .B(n760), .ZN(G329) );
  AND2_X1 U835 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U836 ( .A(G132), .ZN(G219) );
  INV_X1 U837 ( .A(G82), .ZN(G220) );
  INV_X1 U838 ( .A(G57), .ZN(G237) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n762) );
  XNOR2_X1 U840 ( .A(n762), .B(KEYINPUT70), .ZN(n763) );
  XNOR2_X1 U841 ( .A(KEYINPUT10), .B(n763), .ZN(G223) );
  INV_X1 U842 ( .A(G223), .ZN(n836) );
  NAND2_X1 U843 ( .A1(n836), .A2(G567), .ZN(n764) );
  XOR2_X1 U844 ( .A(KEYINPUT11), .B(n764), .Z(G234) );
  INV_X1 U845 ( .A(G860), .ZN(n769) );
  OR2_X1 U846 ( .A1(n972), .A2(n769), .ZN(G153) );
  XNOR2_X1 U847 ( .A(KEYINPUT73), .B(G171), .ZN(G301) );
  NAND2_X1 U848 ( .A1(G868), .A2(G301), .ZN(n766) );
  OR2_X1 U849 ( .A1(n963), .A2(G868), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n766), .A2(n765), .ZN(G284) );
  NAND2_X1 U851 ( .A1(G286), .A2(G868), .ZN(n768) );
  INV_X1 U852 ( .A(G868), .ZN(n809) );
  NAND2_X1 U853 ( .A1(G299), .A2(n809), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U855 ( .A1(n769), .A2(G559), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n770), .A2(n963), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U858 ( .A1(G868), .A2(n972), .ZN(n772) );
  XOR2_X1 U859 ( .A(KEYINPUT75), .B(n772), .Z(n775) );
  NAND2_X1 U860 ( .A1(G868), .A2(n963), .ZN(n773) );
  NOR2_X1 U861 ( .A1(G559), .A2(n773), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n775), .A2(n774), .ZN(G282) );
  NAND2_X1 U863 ( .A1(G123), .A2(n886), .ZN(n776) );
  XNOR2_X1 U864 ( .A(n776), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U865 ( .A1(G111), .A2(n885), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G135), .A2(n890), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n889), .A2(G99), .ZN(n779) );
  XOR2_X1 U869 ( .A(KEYINPUT76), .B(n779), .Z(n780) );
  NOR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n922) );
  XNOR2_X1 U872 ( .A(G2096), .B(n922), .ZN(n784) );
  NOR2_X1 U873 ( .A1(n784), .A2(G2100), .ZN(n785) );
  XNOR2_X1 U874 ( .A(n785), .B(KEYINPUT77), .ZN(G156) );
  NAND2_X1 U875 ( .A1(n963), .A2(G559), .ZN(n806) );
  XNOR2_X1 U876 ( .A(n972), .B(n806), .ZN(n786) );
  NOR2_X1 U877 ( .A1(n786), .A2(G860), .ZN(n798) );
  NAND2_X1 U878 ( .A1(G93), .A2(n787), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G80), .A2(n788), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n797) );
  NAND2_X1 U881 ( .A1(n791), .A2(G67), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(KEYINPUT78), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G55), .A2(n793), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n808) );
  XNOR2_X1 U886 ( .A(n798), .B(n808), .ZN(G145) );
  XNOR2_X1 U887 ( .A(n983), .B(n808), .ZN(n803) );
  XNOR2_X1 U888 ( .A(G166), .B(n972), .ZN(n801) );
  XNOR2_X1 U889 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n799), .B(G288), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U892 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n804), .B(G290), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n805), .B(G305), .ZN(n906) );
  XNOR2_X1 U895 ( .A(n906), .B(n806), .ZN(n807) );
  NOR2_X1 U896 ( .A1(n809), .A2(n807), .ZN(n811) );
  AND2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U898 ( .A1(n811), .A2(n810), .ZN(G295) );
  NAND2_X1 U899 ( .A1(G2078), .A2(G2084), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n812), .B(KEYINPUT81), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n813), .B(KEYINPUT20), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n814), .A2(G2090), .ZN(n815) );
  XNOR2_X1 U903 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U906 ( .A1(G69), .A2(G120), .ZN(n817) );
  NOR2_X1 U907 ( .A1(G237), .A2(n817), .ZN(n818) );
  NAND2_X1 U908 ( .A1(G108), .A2(n818), .ZN(n841) );
  NAND2_X1 U909 ( .A1(n841), .A2(G567), .ZN(n824) );
  NOR2_X1 U910 ( .A1(G220), .A2(G219), .ZN(n819) );
  XOR2_X1 U911 ( .A(KEYINPUT22), .B(n819), .Z(n820) );
  NOR2_X1 U912 ( .A1(G218), .A2(n820), .ZN(n821) );
  NAND2_X1 U913 ( .A1(G96), .A2(n821), .ZN(n840) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n840), .ZN(n822) );
  XNOR2_X1 U915 ( .A(KEYINPUT82), .B(n822), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n842) );
  NAND2_X1 U917 ( .A1(G483), .A2(G661), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n842), .A2(n825), .ZN(n839) );
  NAND2_X1 U919 ( .A1(n839), .A2(G36), .ZN(G176) );
  XOR2_X1 U920 ( .A(KEYINPUT105), .B(G2451), .Z(n827) );
  XNOR2_X1 U921 ( .A(G2446), .B(G2427), .ZN(n826) );
  XNOR2_X1 U922 ( .A(n827), .B(n826), .ZN(n834) );
  XOR2_X1 U923 ( .A(G2438), .B(G2435), .Z(n829) );
  XNOR2_X1 U924 ( .A(G2443), .B(G2430), .ZN(n828) );
  XNOR2_X1 U925 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U926 ( .A(n830), .B(G2454), .Z(n832) );
  XNOR2_X1 U927 ( .A(G1348), .B(G1341), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n835), .A2(G14), .ZN(n911) );
  XOR2_X1 U931 ( .A(KEYINPUT106), .B(n911), .Z(G401) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U934 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n842), .ZN(G319) );
  XOR2_X1 U944 ( .A(G2474), .B(G1961), .Z(n844) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1966), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n845), .B(KEYINPUT109), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1991), .B(G1996), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U950 ( .A(G1976), .B(G1981), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1956), .B(G1971), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U956 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n855) );
  XNOR2_X1 U957 ( .A(G2678), .B(KEYINPUT43), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U959 ( .A(KEYINPUT42), .B(G2072), .Z(n857) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2090), .ZN(n856) );
  XNOR2_X1 U961 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U962 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U963 ( .A(G2096), .B(G2100), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U965 ( .A(G2078), .B(G2084), .Z(n862) );
  XNOR2_X1 U966 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U967 ( .A1(G124), .A2(n886), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n889), .A2(G100), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G112), .A2(n885), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G136), .A2(n890), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U974 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G103), .A2(n889), .ZN(n872) );
  NAND2_X1 U976 ( .A1(G139), .A2(n890), .ZN(n871) );
  NAND2_X1 U977 ( .A1(n872), .A2(n871), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n885), .A2(G115), .ZN(n873) );
  XNOR2_X1 U979 ( .A(n873), .B(KEYINPUT112), .ZN(n875) );
  NAND2_X1 U980 ( .A1(G127), .A2(n886), .ZN(n874) );
  NAND2_X1 U981 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U983 ( .A1(n878), .A2(n877), .ZN(n928) );
  XNOR2_X1 U984 ( .A(n928), .B(n879), .ZN(n880) );
  XNOR2_X1 U985 ( .A(n880), .B(n922), .ZN(n884) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n882) );
  XNOR2_X1 U987 ( .A(KEYINPUT113), .B(KEYINPUT111), .ZN(n881) );
  XNOR2_X1 U988 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U989 ( .A(n884), .B(n883), .Z(n898) );
  NAND2_X1 U990 ( .A1(G118), .A2(n885), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G130), .A2(n886), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G106), .A2(n889), .ZN(n892) );
  NAND2_X1 U994 ( .A1(G142), .A2(n890), .ZN(n891) );
  NAND2_X1 U995 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U996 ( .A(KEYINPUT45), .B(n893), .Z(n894) );
  NOR2_X1 U997 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U998 ( .A(G160), .B(n896), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1000 ( .A(n899), .B(G162), .Z(n902) );
  XNOR2_X1 U1001 ( .A(n900), .B(G164), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n904), .B(n903), .Z(n905) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n905), .ZN(G395) );
  XOR2_X1 U1005 ( .A(KEYINPUT114), .B(n906), .Z(n908) );
  XNOR2_X1 U1006 ( .A(n963), .B(G286), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n909), .B(G171), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n910), .ZN(G397) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n911), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1018 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1029) );
  INV_X1 U1019 ( .A(KEYINPUT55), .ZN(n958) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n935) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n921), .Z(n927) );
  XNOR2_X1 U1024 ( .A(G160), .B(G2084), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1028 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n931), .Z(n932) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n958), .A2(n939), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(G29), .ZN(n1027) );
  XNOR2_X1 U1038 ( .A(G2090), .B(G35), .ZN(n953) );
  XOR2_X1 U1039 ( .A(G2067), .B(G26), .Z(n941) );
  NAND2_X1 U1040 ( .A1(n941), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(G1991), .B(G25), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n948) );
  XOR2_X1 U1044 ( .A(n944), .B(G27), .Z(n946) );
  XNOR2_X1 U1045 ( .A(G1996), .B(G32), .ZN(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n954) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n954), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n958), .B(n957), .ZN(n960) );
  INV_X1 U1055 ( .A(G29), .ZN(n959) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n961), .ZN(n1025) );
  INV_X1 U1058 ( .A(G16), .ZN(n1021) );
  XNOR2_X1 U1059 ( .A(KEYINPUT56), .B(KEYINPUT115), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(n1021), .B(n962), .ZN(n992) );
  XOR2_X1 U1061 ( .A(G1348), .B(n963), .Z(n964) );
  XNOR2_X1 U1062 ( .A(KEYINPUT118), .B(n964), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n990) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(n967), .B(KEYINPUT116), .ZN(n969) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n971) );
  XOR2_X1 U1067 ( .A(KEYINPUT57), .B(KEYINPUT117), .Z(n970) );
  XNOR2_X1 U1068 ( .A(n971), .B(n970), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G1341), .B(n972), .ZN(n974) );
  XOR2_X1 U1070 ( .A(G1961), .B(G171), .Z(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G303), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(KEYINPUT119), .B(n977), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1077 ( .A(KEYINPUT120), .B(n982), .Z(n985) );
  XOR2_X1 U1078 ( .A(n983), .B(G1956), .Z(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n986), .B(KEYINPUT121), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1023) );
  XOR2_X1 U1084 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n1019) );
  XOR2_X1 U1085 ( .A(G1976), .B(G23), .Z(n994) );
  XOR2_X1 U1086 ( .A(G1971), .B(G22), .Z(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G24), .B(G1986), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT58), .B(n997), .Z(n1016) );
  XOR2_X1 U1091 ( .A(n998), .B(G5), .Z(n1013) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(n999), .B(KEYINPUT122), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G20), .B(n1000), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1001) );
  NOR2_X1 U1097 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1099 ( .A(KEYINPUT59), .B(G1348), .Z(n1005) );
  XNOR2_X1 U1100 ( .A(G4), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1101 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1102 ( .A(KEYINPUT60), .B(n1008), .Z(n1009) );
  NOR2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1104 ( .A(KEYINPUT123), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1105 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1106 ( .A(KEYINPUT124), .B(n1014), .Z(n1015) );
  NOR2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(n1017), .B(KEYINPUT61), .ZN(n1018) );
  XNOR2_X1 U1109 ( .A(n1019), .B(n1018), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(n1029), .B(n1028), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

