//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G355));
  NOR2_X1   g0005(.A1(G58), .A2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n209), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G68), .A2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT66), .B2(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n214), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(KEYINPUT0), .ZN(new_n236));
  OR2_X1    g0036(.A1(new_n235), .A2(KEYINPUT0), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n211), .B(new_n233), .C1(new_n236), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n218), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G97), .B(G107), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT72), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G33), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n255), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT7), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(new_n209), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n258), .A2(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT72), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n257), .A2(new_n258), .A3(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(KEYINPUT7), .B1(new_n267), .B2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n268), .A3(G68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT73), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT73), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n263), .A2(new_n268), .A3(new_n271), .A4(G68), .ZN(new_n272));
  AND2_X1   g0072(.A1(G58), .A2(G68), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n273), .B2(new_n206), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G159), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT74), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n270), .A2(KEYINPUT16), .A3(new_n272), .A4(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n210), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n258), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n256), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT7), .B1(new_n284), .B2(new_n209), .ZN(new_n285));
  AOI211_X1 g0085(.A(new_n262), .B(G20), .C1(new_n256), .C2(new_n283), .ZN(new_n286));
  OAI21_X1  g0086(.A(G68), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n277), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT16), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n265), .A2(new_n266), .ZN(new_n293));
  INV_X1    g0093(.A(G223), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n222), .A2(G1698), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n293), .A2(new_n256), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G87), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G1), .A3(G13), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n305));
  INV_X1    g0105(.A(G274), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(G33), .A2(G41), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G41), .A2(G45), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n309), .A2(new_n210), .B1(new_n310), .B2(G1), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n308), .B1(new_n311), .B2(new_n227), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n292), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n302), .B1(new_n298), .B2(new_n299), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n315), .A2(new_n316), .A3(new_n312), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n281), .B1(new_n212), .B2(G20), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n318), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n314), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n291), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(KEYINPUT17), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT75), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n324), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(KEYINPUT17), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n291), .A2(new_n322), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n304), .B2(new_n313), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n315), .A2(new_n335), .A3(new_n312), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(new_n338), .A3(KEYINPUT18), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT18), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n323), .B1(new_n279), .B2(new_n290), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n284), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G238), .A2(G1698), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n345), .B(new_n346), .C1(new_n227), .C2(G1698), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n303), .C1(G107), .C2(new_n345), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n302), .A2(new_n350), .A3(new_n305), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G244), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(new_n308), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n335), .ZN(new_n356));
  INV_X1    g0156(.A(new_n318), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n275), .B1(G20), .B2(G77), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n209), .A2(G33), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT15), .B(G87), .Z(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n319), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n362), .A2(new_n281), .B1(new_n223), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n321), .A2(G77), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT71), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n354), .A2(new_n333), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n356), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n331), .A2(new_n344), .A3(new_n370), .ZN(new_n371));
  XOR2_X1   g0171(.A(KEYINPUT68), .B(G226), .Z(new_n372));
  AOI21_X1  g0172(.A(new_n307), .B1(new_n352), .B2(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n373), .A2(KEYINPUT70), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n295), .A2(G222), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n345), .B(new_n375), .C1(new_n294), .C2(new_n295), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n303), .C1(G77), .C2(new_n345), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(KEYINPUT70), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n333), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n275), .A2(G150), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n381), .B(new_n382), .C1(new_n359), .C2(new_n318), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n281), .B1(new_n221), .B2(new_n363), .ZN(new_n384));
  INV_X1    g0184(.A(new_n321), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n221), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n380), .B(new_n386), .C1(G179), .C2(new_n379), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n386), .B(KEYINPUT9), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n379), .A2(G200), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n316), .C2(new_n379), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n307), .B1(new_n352), .B2(G238), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n227), .A2(G1698), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G226), .B2(G1698), .ZN(new_n398));
  INV_X1    g0198(.A(G97), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n398), .A2(new_n284), .B1(new_n255), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n303), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n395), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n302), .A2(new_n350), .A3(new_n305), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n350), .B1(new_n302), .B2(new_n305), .ZN(new_n404));
  OAI21_X1  g0204(.A(G238), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND4_X1   g0205(.A1(new_n395), .A2(new_n401), .A3(new_n405), .A4(new_n308), .ZN(new_n406));
  OAI21_X1  g0206(.A(G169), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT14), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n402), .A2(new_n406), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G179), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(G169), .C1(new_n402), .C2(new_n406), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G68), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n275), .A2(G50), .B1(G20), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n223), .B2(new_n359), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n281), .ZN(new_n417));
  XOR2_X1   g0217(.A(new_n417), .B(KEYINPUT11), .Z(new_n418));
  INV_X1    g0218(.A(KEYINPUT12), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n363), .B2(new_n414), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n319), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n385), .A2(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n413), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n409), .A2(G190), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(new_n423), .C1(new_n292), .C2(new_n409), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n368), .B1(G190), .B2(new_n355), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n354), .A2(G200), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n371), .A2(new_n394), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G250), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n295), .ZN(new_n436));
  INV_X1    g0236(.A(G257), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G1698), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n293), .A2(new_n256), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G294), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n303), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n212), .A2(G45), .ZN(new_n443));
  OR2_X1    g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  NAND2_X1  g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n446), .A2(new_n303), .A3(new_n218), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(G274), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n442), .A2(new_n316), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n302), .B1(new_n439), .B2(new_n440), .ZN(new_n451));
  INV_X1    g0251(.A(new_n449), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n451), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n453), .B2(G200), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n212), .A2(G33), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n319), .A2(new_n455), .A3(new_n210), .A4(new_n280), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n456), .A2(KEYINPUT76), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(KEYINPUT76), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G107), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n319), .A2(G107), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT25), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT22), .ZN(new_n464));
  INV_X1    g0264(.A(G87), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n464), .A2(new_n465), .A3(G20), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n293), .A2(new_n256), .A3(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n256), .A2(new_n283), .A3(new_n209), .A4(G87), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n464), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n217), .A2(G20), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n467), .A2(new_n469), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT24), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n267), .A2(new_n466), .B1(new_n468), .B2(new_n464), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(KEYINPUT24), .A3(new_n472), .A4(new_n473), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n478), .A3(new_n281), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n454), .A2(new_n461), .A3(new_n463), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n461), .A3(new_n463), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n451), .A2(new_n447), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n449), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n333), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n453), .A2(new_n335), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT80), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n437), .A2(new_n295), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n218), .A2(G1698), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n293), .A2(new_n256), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n284), .A2(G303), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n303), .ZN(new_n494));
  INV_X1    g0294(.A(G45), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1), .ZN(new_n496));
  INV_X1    g0296(.A(new_n445), .ZN(new_n497));
  NOR2_X1   g0297(.A1(KEYINPUT5), .A2(G41), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(G270), .A3(new_n302), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n449), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n494), .A2(G179), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n363), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n282), .A2(G116), .A3(new_n455), .A4(new_n319), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n280), .A2(new_n210), .B1(G20), .B2(new_n504), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n508), .B(new_n209), .C1(G33), .C2(new_n399), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n507), .A2(KEYINPUT20), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT20), .B1(new_n507), .B2(new_n509), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n505), .B(new_n506), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n488), .B1(new_n503), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n501), .B1(new_n493), .B2(new_n303), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(KEYINPUT80), .A3(G179), .A4(new_n512), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(G190), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n513), .C1(new_n292), .C2(new_n515), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n512), .A2(G169), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(new_n515), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n494), .A2(new_n502), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(KEYINPUT21), .A3(G169), .A4(new_n512), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n517), .A2(new_n519), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n487), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(G107), .B1(new_n285), .B2(new_n286), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n275), .A2(G77), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n399), .A2(new_n217), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n202), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n217), .A2(G97), .ZN(new_n531));
  MUX2_X1   g0331(.A(new_n530), .B(new_n531), .S(KEYINPUT6), .Z(new_n532));
  OAI211_X1 g0332(.A(new_n527), .B(new_n528), .C1(new_n532), .C2(new_n209), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n281), .B1(G97), .B2(new_n460), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n363), .A2(new_n399), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G244), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n256), .A2(new_n283), .A3(G250), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT4), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G1698), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n538), .A2(G1698), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n543), .A2(new_n256), .A3(new_n283), .A4(G244), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n544), .A2(new_n508), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n539), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n303), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n446), .A2(new_n303), .A3(new_n437), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n452), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n316), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n536), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT4), .B1(new_n267), .B2(G244), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n544), .A2(new_n508), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n295), .B1(new_n540), .B2(KEYINPUT4), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT77), .B1(new_n556), .B2(new_n302), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT77), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n546), .A2(new_n558), .A3(new_n303), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n549), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n557), .A2(new_n335), .A3(new_n549), .A4(new_n559), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n534), .A2(new_n535), .B1(new_n550), .B2(new_n333), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n552), .A2(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G238), .A2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n224), .B2(G1698), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n267), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G116), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n302), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n443), .A2(G274), .ZN(new_n570));
  AOI211_X1 g0370(.A(new_n570), .B(new_n303), .C1(new_n435), .C2(new_n443), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n292), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(G190), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT79), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n576), .A3(G190), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n293), .A2(new_n209), .A3(G68), .A4(new_n256), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n359), .B2(new_n399), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n209), .B1(new_n255), .B2(new_n399), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT78), .B(G87), .ZN(new_n583));
  OAI211_X1 g0383(.A(KEYINPUT19), .B(new_n582), .C1(new_n583), .C2(new_n203), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n579), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(new_n281), .B1(new_n363), .B2(new_n361), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n457), .A2(G87), .A3(new_n458), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n572), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n460), .A2(new_n360), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n333), .A2(new_n589), .B1(new_n590), .B2(new_n586), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n572), .A2(new_n335), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n578), .A2(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n434), .A2(new_n526), .A3(new_n564), .A4(new_n593), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n594), .B(KEYINPUT81), .ZN(G372));
  INV_X1    g0395(.A(new_n573), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n586), .A2(KEYINPUT82), .A3(new_n587), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT82), .B1(new_n586), .B2(new_n587), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT83), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n575), .A2(new_n577), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT83), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n552), .A2(new_n561), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n486), .A2(new_n522), .A3(new_n524), .A4(new_n517), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n480), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n563), .A2(new_n562), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT26), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n578), .A2(new_n588), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n563), .A2(new_n562), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT26), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n591), .A2(new_n592), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n433), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n617), .B(KEYINPUT84), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n339), .A2(new_n342), .A3(KEYINPUT85), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT85), .B1(new_n339), .B2(new_n342), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n427), .A2(new_n370), .B1(new_n413), .B2(new_n424), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n331), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n392), .A2(new_n393), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n388), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n625), .ZN(G369));
  INV_X1    g0426(.A(G13), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(G20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n212), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n513), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n525), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n517), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n524), .A2(new_n522), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(KEYINPUT86), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(KEYINPUT86), .ZN(new_n643));
  INV_X1    g0443(.A(G330), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n481), .A2(new_n634), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n480), .A2(new_n486), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT87), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n480), .A2(new_n486), .A3(KEYINPUT87), .A4(new_n646), .ZN(new_n650));
  INV_X1    g0450(.A(new_n486), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n634), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT88), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n649), .A2(KEYINPUT88), .A3(new_n650), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n645), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n486), .A2(new_n634), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n658), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n234), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n583), .A2(G116), .A3(new_n203), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n208), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n635), .B1(new_n610), .B2(new_n615), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT90), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT29), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n674), .B(new_n635), .C1(new_n610), .C2(new_n615), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n611), .A2(new_n612), .ZN(new_n677));
  OAI221_X1 g0477(.A(new_n614), .B1(new_n677), .B2(KEYINPUT26), .C1(new_n607), .C2(new_n608), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n609), .A2(KEYINPUT26), .ZN(new_n679));
  OAI211_X1 g0479(.A(KEYINPUT29), .B(new_n635), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n526), .A2(new_n564), .A3(new_n593), .A4(new_n635), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n503), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n515), .A2(KEYINPUT89), .A3(G179), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n547), .A2(new_n572), .A3(new_n482), .A4(new_n549), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT89), .B1(new_n515), .B2(G179), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n302), .B1(new_n491), .B2(new_n492), .ZN(new_n691));
  NOR4_X1   g0491(.A1(new_n691), .A2(new_n501), .A3(new_n684), .A4(new_n335), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AND4_X1   g0493(.A1(new_n482), .A2(new_n547), .A3(new_n549), .A4(new_n572), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT30), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n572), .A2(G179), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n560), .A2(new_n483), .A3(new_n523), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n689), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n634), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n682), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n681), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n670), .B1(new_n706), .B2(G1), .ZN(G364));
  NAND2_X1  g0507(.A1(new_n628), .A2(G45), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT91), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n665), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n645), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n644), .B1(new_n642), .B2(new_n643), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n664), .A2(new_n284), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G355), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n250), .A2(G45), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT92), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n664), .A2(new_n267), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G45), .B2(new_n208), .ZN(new_n721));
  OAI221_X1 g0521(.A(new_n717), .B1(G116), .B2(new_n234), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n627), .A2(new_n255), .A3(KEYINPUT93), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G13), .B2(G33), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n210), .B1(G20), .B2(new_n333), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n335), .A2(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n209), .A2(G190), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G311), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR4_X1   g0536(.A1(new_n209), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT95), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT95), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G329), .ZN(new_n741));
  INV_X1    g0541(.A(G283), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n292), .A2(G179), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n733), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n740), .A2(new_n741), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n316), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n209), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n736), .B(new_n745), .C1(G294), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(G20), .A2(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G303), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n750), .A2(new_n335), .A3(new_n292), .A4(KEYINPUT94), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT94), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n335), .A2(new_n292), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(new_n751), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G326), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n732), .A2(new_n751), .ZN(new_n762));
  INV_X1    g0562(.A(G322), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n284), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n733), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n749), .A2(new_n754), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n765), .A2(new_n414), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n748), .A2(G97), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n223), .B2(new_n734), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n284), .B(new_n772), .C1(new_n760), .C2(G50), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n740), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n776));
  XNOR2_X1  g0576(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n753), .A2(new_n583), .ZN(new_n778));
  INV_X1    g0578(.A(new_n744), .ZN(new_n779));
  INV_X1    g0579(.A(new_n762), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n779), .A2(G107), .B1(new_n780), .B2(G58), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n773), .A2(new_n777), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n769), .B1(new_n770), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n729), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n637), .A2(new_n640), .A3(new_n728), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n731), .A2(new_n784), .A3(new_n785), .A4(new_n712), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n715), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n370), .A2(new_n635), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n430), .A2(new_n431), .B1(new_n368), .B2(new_n634), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n370), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n635), .B(new_n792), .C1(new_n610), .C2(new_n615), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n672), .A2(new_n675), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n791), .ZN(new_n796));
  INV_X1    g0596(.A(new_n704), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  INV_X1    g0599(.A(new_n712), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n726), .A2(new_n729), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n712), .B1(G77), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT97), .Z(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n729), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G150), .A2(new_n766), .B1(new_n780), .B2(G143), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n808), .B1(new_n774), .B2(new_n734), .C1(new_n759), .C2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT34), .Z(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G50), .B2(new_n753), .ZN(new_n812));
  INV_X1    g0612(.A(new_n740), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G132), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n748), .A2(G58), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n261), .B1(G68), .B2(new_n779), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n812), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n217), .A2(new_n752), .B1(new_n762), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G283), .B2(new_n766), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n771), .B(new_n820), .C1(new_n740), .C2(new_n735), .ZN(new_n821));
  INV_X1    g0621(.A(new_n734), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(G116), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n779), .A2(G87), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n760), .A2(G303), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n823), .A2(new_n284), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n807), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n806), .B(new_n827), .C1(new_n726), .C2(new_n791), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n801), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT98), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n801), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(G384));
  NAND3_X1  g0634(.A1(new_n676), .A2(new_n434), .A3(new_n680), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n625), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT39), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n324), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT75), .B1(new_n291), .B2(new_n324), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT17), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n326), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n619), .B2(new_n620), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n341), .A2(new_n632), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n332), .A2(new_n338), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n325), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT37), .B1(new_n847), .B2(new_n844), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n844), .A2(KEYINPUT37), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n330), .A2(new_n849), .A3(new_n846), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n270), .A2(new_n272), .A3(new_n278), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n289), .A2(KEYINPUT100), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n270), .A2(new_n272), .A3(new_n278), .A4(new_n854), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n281), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n632), .B1(new_n858), .B2(new_n322), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n322), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n338), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n862), .A3(new_n330), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n328), .A2(new_n329), .B1(new_n332), .B2(new_n338), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n863), .A2(KEYINPUT37), .B1(new_n849), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n860), .B1(new_n842), .B2(new_n343), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n837), .B1(new_n852), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n425), .A2(new_n634), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n838), .A2(new_n839), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n337), .B1(new_n858), .B2(new_n322), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n872), .A2(new_n859), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n850), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n859), .B1(new_n331), .B2(new_n344), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n871), .A2(new_n878), .A3(KEYINPUT39), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n869), .A2(new_n870), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n632), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n621), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT99), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n423), .B2(new_n635), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n424), .A2(KEYINPUT99), .A3(new_n634), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n425), .A2(new_n427), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n413), .A2(new_n424), .A3(new_n634), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n793), .B2(new_n789), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n871), .A2(new_n878), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n880), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n836), .B(new_n893), .Z(new_n894));
  NOR2_X1   g0694(.A1(new_n852), .A2(new_n868), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n791), .B1(new_n886), .B2(new_n887), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n703), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT101), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n703), .A2(new_n896), .A3(KEYINPUT101), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n897), .B1(new_n871), .B2(new_n878), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n895), .A2(new_n901), .B1(new_n902), .B2(KEYINPUT40), .ZN(new_n903));
  INV_X1    g0703(.A(new_n703), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n433), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(G330), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n894), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n212), .B2(new_n628), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT35), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n209), .B(new_n210), .C1(new_n532), .C2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n911), .B(G116), .C1(new_n910), .C2(new_n532), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT36), .ZN(new_n913));
  OAI21_X1  g0713(.A(G77), .B1(new_n226), .B2(new_n414), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n208), .A2(new_n914), .B1(G50), .B2(new_n414), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(G1), .A3(new_n627), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n913), .A3(new_n916), .ZN(G367));
  NAND2_X1  g0717(.A1(new_n536), .A2(new_n634), .ZN(new_n918));
  INV_X1    g0718(.A(new_n561), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n534), .B(new_n535), .C1(new_n316), .C2(new_n550), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n612), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n608), .A2(new_n634), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT103), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT103), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n658), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n660), .B1(new_n655), .B2(new_n656), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n921), .A2(new_n922), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT103), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n923), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n928), .A2(KEYINPUT42), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT42), .B1(new_n928), .B2(new_n932), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n608), .B1(new_n932), .B2(new_n651), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n933), .A2(new_n934), .B1(new_n634), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT43), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n597), .A2(new_n598), .A3(new_n635), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n614), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT102), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n604), .A2(new_n614), .A3(new_n942), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n946), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n939), .B2(new_n940), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n927), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n934), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n928), .A2(KEYINPUT42), .A3(new_n932), .ZN(new_n952));
  INV_X1    g0752(.A(new_n935), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n635), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT43), .B1(new_n954), .B2(KEYINPUT104), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n949), .B(new_n927), .C1(new_n957), .C2(new_n948), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n665), .B(KEYINPUT41), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n662), .A2(new_n932), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT105), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT105), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n662), .A2(new_n964), .A3(new_n932), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n963), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT45), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n928), .A2(new_n926), .A3(KEYINPUT105), .A4(new_n659), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n964), .B1(new_n662), .B2(new_n932), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n926), .B1(new_n928), .B2(new_n659), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n966), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n658), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n657), .A2(new_n661), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n928), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n645), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n705), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n966), .A2(new_n970), .A3(new_n973), .A4(new_n658), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n976), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n961), .B1(new_n982), .B2(new_n706), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n950), .A2(new_n959), .B1(new_n983), .B2(new_n711), .ZN(new_n984));
  INV_X1    g0784(.A(new_n720), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n730), .B1(new_n234), .B2(new_n361), .C1(new_n245), .C2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT106), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n712), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT107), .ZN(new_n989));
  INV_X1    g0789(.A(new_n728), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n760), .A2(G143), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n748), .A2(G68), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT108), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n765), .A2(new_n774), .B1(new_n734), .B2(new_n221), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .C1(new_n740), .C2(new_n809), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n991), .B(new_n995), .C1(new_n993), .C2(new_n994), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n780), .A2(G150), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n284), .B1(new_n779), .B2(G77), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n753), .A2(G58), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n997), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n813), .A2(G317), .B1(G303), .B2(new_n780), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n742), .B2(new_n734), .C1(new_n818), .C2(new_n765), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G107), .B2(new_n748), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n753), .A2(G116), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT46), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n744), .A2(new_n399), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(new_n267), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n759), .A2(new_n735), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1000), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n989), .B1(new_n990), .B2(new_n946), .C1(new_n1012), .C2(new_n807), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n984), .A2(new_n1013), .ZN(G387));
  INV_X1    g0814(.A(new_n980), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n705), .A2(new_n979), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n665), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n667), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n716), .A2(new_n1018), .B1(new_n217), .B2(new_n664), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT110), .Z(new_n1020));
  NOR2_X1   g0820(.A1(new_n414), .A2(new_n223), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n318), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT50), .B1(new_n318), .B2(G50), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1022), .A2(new_n667), .A3(new_n495), .A4(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n720), .B1(new_n1021), .B2(new_n1024), .C1(new_n242), .C2(new_n495), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n729), .B(new_n728), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n753), .A2(G77), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n414), .B2(new_n734), .C1(new_n759), .C2(new_n774), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n357), .B2(new_n766), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n762), .A2(new_n221), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1006), .B(new_n1030), .C1(new_n813), .C2(G150), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n748), .A2(new_n360), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n1031), .A3(new_n267), .A4(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G311), .A2(new_n766), .B1(new_n780), .B2(G317), .ZN(new_n1034));
  INV_X1    g0834(.A(G303), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n734), .C1(new_n759), .C2(new_n763), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n742), .B2(new_n747), .C1(new_n818), .C2(new_n752), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n813), .A2(G326), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n779), .A2(G116), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1040), .A2(new_n261), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n800), .B(new_n1026), .C1(new_n1045), .C2(new_n729), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n655), .A2(new_n656), .A3(new_n728), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n711), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1017), .B(new_n1048), .C1(new_n1049), .C2(new_n979), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n976), .A2(new_n981), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n976), .A2(KEYINPUT111), .A3(new_n981), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n711), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1051), .A2(new_n1015), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(new_n665), .A3(new_n982), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n800), .B1(new_n926), .B2(new_n728), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n730), .B1(new_n399), .B2(new_n234), .C1(new_n985), .C2(new_n253), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n760), .A2(G317), .B1(G311), .B2(new_n780), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n345), .B(new_n1061), .C1(G322), .C2(new_n813), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n742), .B2(new_n752), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n765), .A2(new_n1035), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n734), .A2(new_n818), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n747), .A2(new_n504), .B1(new_n217), .B2(new_n744), .ZN(new_n1066));
  NOR4_X1   g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(G150), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n759), .A2(new_n1068), .B1(new_n774), .B2(new_n762), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n748), .A2(G77), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n813), .A2(G143), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1070), .A2(new_n267), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n734), .A2(new_n318), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n752), .A2(new_n414), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n824), .B1(new_n221), .B2(new_n765), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n729), .B1(new_n1067), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1058), .A2(new_n1059), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1055), .A2(new_n1057), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(KEYINPUT112), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT112), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1055), .A2(new_n1057), .A3(new_n1082), .A4(new_n1079), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(G390));
  NAND2_X1  g0884(.A1(new_n845), .A2(new_n851), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n867), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n1086), .B2(new_n878), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n879), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n726), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n802), .A2(new_n318), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n760), .A2(G283), .B1(G107), .B2(new_n766), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n399), .B2(new_n734), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT113), .Z(new_n1093));
  OAI21_X1  g0893(.A(new_n284), .B1(new_n752), .B2(new_n465), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(KEYINPUT114), .A2(new_n1094), .B1(new_n748), .B2(G77), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n414), .C2(new_n744), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n762), .A2(new_n504), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1094), .A2(KEYINPUT114), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n740), .A2(new_n818), .ZN(new_n1099));
  NOR4_X1   g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n284), .B1(new_n813), .B2(G125), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  NAND2_X1  g0902(.A1(new_n822), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n774), .C2(new_n747), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n752), .B2(new_n1068), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n753), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G137), .A2(new_n766), .B1(new_n780), .B2(G132), .ZN(new_n1109));
  INV_X1    g0909(.A(G128), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(new_n1109), .C1(new_n1110), .C2(new_n759), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G50), .B2(new_n779), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n729), .B1(new_n1100), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1089), .A2(new_n712), .A3(new_n1090), .A4(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n790), .A2(new_n370), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n635), .B(new_n1115), .C1(new_n678), .C2(new_n679), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n889), .B1(new_n1116), .B2(new_n789), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n843), .A2(new_n844), .B1(new_n850), .B2(new_n848), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n878), .B1(new_n1118), .B2(KEYINPUT38), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n870), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1087), .A2(new_n1088), .B1(new_n870), .B2(new_n890), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n797), .A2(new_n896), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1124), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n890), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1127), .A2(new_n1120), .B1(new_n869), .B2(new_n879), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1114), .B1(new_n1131), .B2(new_n1049), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n905), .A2(G330), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n835), .A2(new_n625), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n889), .B1(new_n704), .B2(new_n791), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1124), .A2(new_n1135), .B1(new_n789), .B2(new_n793), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1116), .A2(new_n789), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n1130), .A3(new_n1125), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1141), .A2(new_n665), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1131), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1132), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(G378));
  INV_X1    g0946(.A(new_n1134), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT115), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n903), .B2(new_n644), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1119), .A2(KEYINPUT40), .A3(new_n899), .A4(new_n900), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(KEYINPUT115), .A4(G330), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1154));
  XNOR2_X1  g0954(.A(new_n394), .B(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n386), .A2(new_n881), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n903), .A2(new_n644), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1157), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(KEYINPUT115), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n893), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n893), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1148), .B(KEYINPUT57), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n893), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT116), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n880), .A2(new_n1169), .A3(new_n892), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n880), .B2(new_n892), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1172), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1168), .A2(new_n1173), .B1(new_n1147), .B2(new_n1141), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1165), .B(new_n665), .C1(new_n1174), .C2(KEYINPUT57), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1157), .A2(new_n727), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G41), .B1(new_n293), .B2(G33), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(G50), .ZN(new_n1178));
  AOI21_X1  g0978(.A(G41), .B1(new_n813), .B2(G124), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n760), .A2(G125), .B1(G137), .B2(new_n822), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n753), .A2(new_n1102), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n766), .A2(G132), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n748), .A2(G150), .B1(new_n780), .B2(G128), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n255), .B(new_n1179), .C1(new_n1184), .C2(KEYINPUT59), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G159), .B2(new_n779), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1178), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n813), .A2(G283), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n760), .A2(G116), .B1(G107), .B2(new_n780), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n779), .A2(G58), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1027), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n267), .B1(new_n360), .B2(new_n822), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G41), .B1(new_n766), .B2(G97), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n992), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT58), .Z(new_n1197));
  AOI21_X1  g0997(.A(new_n807), .B1(new_n1188), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n803), .A2(G50), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1176), .A2(new_n800), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n1201), .B2(new_n711), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1175), .A2(new_n1202), .ZN(G375));
  OAI21_X1  g1003(.A(new_n284), .B1(new_n752), .B2(new_n399), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1032), .B1(new_n742), .B2(new_n762), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT117), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n223), .B2(new_n744), .C1(new_n818), .C2(new_n759), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1204), .B(new_n1207), .C1(G303), .C2(new_n813), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n217), .B2(new_n734), .C1(new_n504), .C2(new_n765), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1191), .B1(new_n221), .B2(new_n747), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n261), .B(new_n1210), .C1(G150), .C2(new_n822), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n1110), .B2(new_n740), .C1(new_n774), .C2(new_n752), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT118), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n760), .A2(G132), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n766), .A2(new_n1102), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n780), .A2(G137), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n807), .B1(new_n1209), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n888), .A2(new_n727), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n803), .A2(G68), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n800), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1139), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1222), .B2(new_n711), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n960), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1225), .B2(new_n1140), .ZN(G381));
  NAND4_X1  g1026(.A1(new_n1081), .A2(new_n984), .A3(new_n1013), .A4(new_n1083), .ZN(new_n1227));
  OR2_X1    g1027(.A1(G393), .A2(G396), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1227), .A2(G384), .A3(G381), .A4(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT119), .ZN(new_n1230));
  INV_X1    g1030(.A(G375), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1145), .A3(new_n1231), .ZN(G407));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1145), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  INV_X1    g1034(.A(KEYINPUT123), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(G387), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(G390), .A2(new_n1236), .A3(KEYINPUT124), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT123), .B1(new_n984), .B2(new_n1013), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1083), .B(new_n1081), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(new_n787), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G387), .B2(new_n1239), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1237), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G390), .A2(G387), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n1227), .A3(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1172), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n960), .B(new_n1148), .C1(new_n1248), .C2(new_n1164), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT120), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1168), .A2(new_n1162), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1200), .B1(new_n1251), .B2(new_n711), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT120), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1201), .A2(new_n1253), .A3(new_n960), .A4(new_n1148), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1145), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT121), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1175), .A2(G378), .A3(new_n1202), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n633), .A2(G213), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1224), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1134), .A2(new_n1139), .A3(KEYINPUT60), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1143), .A2(new_n1265), .A3(new_n665), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1223), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G384), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G384), .A2(new_n1268), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1263), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1262), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1273), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT122), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1271), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(KEYINPUT122), .A3(new_n1269), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1281), .A2(new_n1283), .A3(G2897), .A4(new_n1262), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1262), .A2(G2897), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1272), .A2(KEYINPUT122), .A3(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1278), .B(new_n1279), .C1(new_n1287), .C2(new_n1276), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1247), .B1(new_n1275), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT121), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1261), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1295), .A2(KEYINPUT63), .B1(new_n1273), .B2(new_n1263), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n1262), .B(new_n1272), .C1(new_n1256), .C2(new_n1258), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(KEYINPUT63), .ZN(new_n1300));
  AND4_X1   g1100(.A1(new_n1298), .A2(new_n1276), .A3(KEYINPUT63), .A4(new_n1273), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1297), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1296), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT63), .B1(new_n1263), .B2(new_n1287), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1274), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1246), .A2(new_n1279), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT63), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT125), .B1(new_n1277), .B2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1299), .A2(new_n1298), .A3(KEYINPUT63), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1307), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT126), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1289), .B1(new_n1304), .B2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(new_n1273), .A2(KEYINPUT127), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1246), .B(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G375), .A2(G378), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1233), .B(new_n1316), .C1(KEYINPUT127), .C2(new_n1273), .ZN(new_n1317));
  XOR2_X1   g1117(.A(new_n1315), .B(new_n1317), .Z(G402));
endmodule


