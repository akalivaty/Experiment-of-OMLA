//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n187), .B1(new_n189), .B2(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n191), .A2(new_n188), .A3(KEYINPUT80), .A4(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(new_n194), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n190), .B(new_n192), .C1(new_n195), .C2(new_n191), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G119), .B(G128), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT23), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n200), .A2(KEYINPUT23), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(KEYINPUT23), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n202), .A2(G119), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G110), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n199), .B(KEYINPUT78), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n198), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  OAI22_X1  g025(.A1(new_n206), .A2(G110), .B1(new_n208), .B2(new_n209), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n196), .A2(new_n197), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n189), .A2(new_n194), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n197), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT22), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT72), .B(G953), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT81), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n222), .A3(G221), .A4(G234), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n218), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n218), .A3(new_n223), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(G137), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n221), .A2(new_n218), .A3(new_n223), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n224), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n217), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n211), .A2(new_n227), .A3(new_n216), .A4(new_n230), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(G234), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G902), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n239), .A2(KEYINPUT83), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n236), .A3(new_n233), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT82), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT82), .B(KEYINPUT25), .Z(new_n245));
  OAI211_X1 g059(.A(new_n244), .B(new_n237), .C1(new_n241), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(KEYINPUT83), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n240), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT1), .B1(new_n252), .B2(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n197), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT1), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(G128), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(G146), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n255), .A2(new_n259), .A3(new_n260), .A4(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n250), .A2(new_n263), .A3(new_n260), .A4(G128), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n251), .A2(new_n258), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n228), .A2(G134), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT64), .B1(new_n228), .B2(G134), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n267), .A3(G137), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT11), .B1(new_n267), .B2(G137), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT11), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n228), .A3(G134), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n271), .B1(new_n280), .B2(G131), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n249), .B1(new_n265), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n255), .A2(new_n259), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  OR2_X1    g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n252), .A2(G146), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n197), .A2(G143), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT65), .A2(G131), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n275), .A2(new_n279), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n290), .B1(new_n275), .B2(new_n279), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n284), .B(new_n289), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n272), .A2(new_n274), .B1(new_n276), .B2(new_n278), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n270), .B1(new_n294), .B2(new_n266), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n262), .A2(new_n264), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n203), .B1(new_n253), .B2(KEYINPUT67), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n250), .B1(new_n297), .B2(new_n257), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT68), .B(new_n295), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n282), .A2(new_n293), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT30), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT2), .B(G113), .Z(new_n303));
  XNOR2_X1  g117(.A(G116), .B(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G119), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G116), .ZN(new_n307));
  INV_X1    g121(.A(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n286), .A2(new_n285), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n284), .B(KEYINPUT69), .C1(new_n315), .C2(new_n250), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT69), .B1(new_n289), .B2(new_n284), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n292), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n294), .A2(new_n290), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n258), .A2(new_n251), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n262), .A2(new_n264), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n319), .A2(new_n322), .B1(new_n325), .B2(new_n295), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n314), .B1(new_n326), .B2(KEYINPUT30), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n284), .B1(new_n315), .B2(new_n250), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n331), .B(new_n316), .C1(new_n291), .C2(new_n292), .ZN(new_n332));
  AND4_X1   g146(.A1(new_n314), .A2(new_n328), .A3(KEYINPUT30), .A4(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n302), .B(new_n313), .C1(new_n327), .C2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n313), .B(KEYINPUT71), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n332), .A3(new_n328), .ZN(new_n336));
  INV_X1    g150(.A(G237), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n219), .A2(G210), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G101), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n343), .A2(KEYINPUT74), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n334), .A2(new_n336), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT31), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n328), .A2(KEYINPUT75), .A3(new_n332), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT75), .B1(new_n328), .B2(new_n332), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT28), .B1(new_n349), .B2(new_n335), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n300), .A2(new_n313), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(new_n336), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n342), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT31), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n334), .A2(new_n355), .A3(new_n336), .A4(new_n344), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(G472), .A2(G902), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT76), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT32), .B1(new_n357), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n343), .B1(new_n350), .B2(new_n353), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n334), .A2(new_n336), .A3(new_n342), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n328), .A2(new_n332), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n328), .A2(KEYINPUT75), .A3(new_n332), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n335), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n351), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n304), .B(new_n311), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT71), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n351), .B1(new_n375), .B2(new_n336), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n372), .A2(new_n377), .A3(KEYINPUT29), .A4(new_n343), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT77), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n376), .B1(new_n351), .B2(new_n371), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT77), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT29), .A4(new_n343), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G472), .B1(new_n366), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n248), .B1(new_n362), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G210), .B1(G237), .B2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n265), .A2(new_n193), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n329), .A2(G125), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G224), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G953), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n390), .B(new_n392), .Z(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(KEYINPUT3), .A2(G107), .ZN(new_n396));
  NOR2_X1   g210(.A1(KEYINPUT3), .A2(G107), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n396), .B1(G104), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(G101), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT84), .B(G104), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n398), .B(new_n399), .C1(new_n400), .C2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(G104), .A2(G107), .ZN(new_n402));
  OAI211_X1 g216(.A(G101), .B(new_n402), .C1(new_n400), .C2(G107), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n306), .A3(G116), .ZN(new_n406));
  OAI211_X1 g220(.A(G113), .B(new_n406), .C1(new_n310), .C2(new_n405), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n305), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n411));
  INV_X1    g225(.A(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(G104), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT3), .A2(G107), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n413), .B(new_n414), .C1(new_n400), .C2(new_n397), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n410), .B1(new_n415), .B2(G101), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n373), .B1(new_n416), .B2(new_n401), .ZN(new_n417));
  INV_X1    g231(.A(G104), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT84), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G104), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n397), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n413), .A2(new_n414), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n410), .B(G101), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT86), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n415), .A2(new_n426), .A3(new_n410), .A4(G101), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI221_X4 g242(.A(KEYINPUT89), .B1(new_n404), .B2(new_n409), .C1(new_n417), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT89), .ZN(new_n430));
  OAI21_X1  g244(.A(G101), .B1(new_n422), .B2(new_n423), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n401), .A2(new_n431), .A3(KEYINPUT4), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n313), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n401), .A2(new_n305), .A3(new_n403), .A4(new_n407), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n395), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n434), .A3(new_n394), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT6), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT6), .B(new_n395), .C1(new_n429), .C2(new_n435), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n393), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n401), .A2(new_n403), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n408), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT90), .A3(new_n434), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n394), .B(KEYINPUT8), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n445), .C1(KEYINPUT90), .C2(new_n443), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT7), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n390), .B1(new_n447), .B2(new_n392), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n392), .A2(new_n447), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n388), .A2(new_n389), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n446), .A2(new_n448), .A3(new_n437), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n236), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n387), .B1(new_n441), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n425), .A2(new_n427), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n432), .A2(new_n313), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n434), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT89), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n433), .A2(new_n430), .A3(new_n434), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n394), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n438), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n440), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n393), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n452), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n386), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n453), .A2(new_n465), .A3(KEYINPUT91), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n387), .B(new_n452), .C1(new_n461), .C2(new_n462), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT91), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G214), .B1(G237), .B2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n253), .A2(G128), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n251), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n324), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n404), .A2(new_n477), .A3(KEYINPUT87), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n262), .A2(new_n264), .B1(new_n251), .B2(new_n475), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n442), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n265), .A2(new_n442), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT12), .A3(new_n322), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n478), .A2(new_n481), .B1(new_n265), .B2(new_n442), .ZN(new_n487));
  INV_X1    g301(.A(new_n322), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT10), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n428), .A2(new_n319), .A3(new_n432), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n265), .A2(new_n442), .A3(new_n491), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n322), .B(KEYINPUT88), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n219), .A2(G227), .ZN(new_n498));
  XNOR2_X1  g312(.A(G110), .B(G140), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n490), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n492), .A2(new_n493), .A3(new_n495), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n322), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n500), .B1(new_n503), .B2(new_n497), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n474), .B(new_n236), .C1(new_n501), .C2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT12), .B1(new_n484), .B2(new_n322), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n487), .A2(new_n486), .A3(new_n488), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n497), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n500), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT10), .B1(new_n478), .B2(new_n481), .ZN(new_n510));
  INV_X1    g324(.A(new_n493), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n510), .A2(new_n511), .A3(new_n494), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n509), .B1(new_n512), .B2(new_n496), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n508), .A2(new_n509), .B1(new_n513), .B2(new_n503), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G469), .ZN(new_n515));
  NAND2_X1  g329(.A1(G469), .A2(G902), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n518));
  AND2_X1   g332(.A1(KEYINPUT72), .A2(G953), .ZN(new_n519));
  NOR2_X1   g333(.A1(KEYINPUT72), .A2(G953), .ZN(new_n520));
  OAI211_X1 g334(.A(G214), .B(new_n337), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n252), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n219), .A2(G143), .A3(G214), .A4(new_n337), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n266), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n518), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT18), .A2(G131), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n195), .A2(G146), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n529), .A2(new_n530), .B1(new_n215), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n524), .A2(KEYINPUT92), .A3(KEYINPUT18), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n522), .A2(new_n523), .A3(new_n266), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n196), .A2(new_n197), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n213), .A4(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G113), .B(G122), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT94), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n418), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n534), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n534), .B2(new_n540), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n236), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G475), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT19), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n214), .A2(KEYINPUT93), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n195), .B2(KEYINPUT19), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n550), .B(new_n552), .C1(new_n549), .C2(new_n214), .ZN(new_n553));
  INV_X1    g367(.A(new_n536), .ZN(new_n554));
  OAI221_X1 g368(.A(new_n213), .B1(new_n553), .B2(G146), .C1(new_n524), .C2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n543), .B1(new_n534), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n548), .B1(new_n544), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT20), .B(new_n548), .C1(new_n544), .C2(new_n556), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n547), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(G234), .A2(G237), .ZN(new_n562));
  INV_X1    g376(.A(G953), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(G952), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n219), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(G902), .A3(new_n562), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT21), .B(G898), .Z(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n565), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n252), .A2(G128), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n203), .A2(G143), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT96), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n267), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n572), .A2(new_n573), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT96), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(G134), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G122), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G116), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n308), .A2(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G107), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT14), .B1(new_n583), .B2(G116), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT97), .ZN(new_n589));
  OR3_X1    g403(.A1(new_n583), .A2(KEYINPUT14), .A3(G116), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n591), .B(KEYINPUT14), .C1(new_n583), .C2(G116), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n589), .A2(new_n584), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n587), .B1(new_n593), .B2(G107), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n582), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n586), .B(G107), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n252), .A2(KEYINPUT13), .A3(G128), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n203), .B2(G143), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n572), .A2(KEYINPUT95), .A3(new_n598), .ZN(new_n602));
  AND4_X1   g416(.A1(new_n597), .A2(new_n601), .A3(new_n602), .A4(new_n573), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n596), .B(new_n577), .C1(new_n603), .C2(new_n267), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT9), .B(G234), .Z(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(G217), .A3(new_n563), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n595), .A2(new_n604), .A3(new_n609), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n236), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G478), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n613), .B(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n561), .A2(new_n571), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G221), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n606), .B2(new_n236), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n517), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n385), .A2(new_n473), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(new_n399), .Z(G3));
  NAND2_X1  g437(.A1(new_n357), .A2(new_n359), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(G472), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n357), .A2(new_n236), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(KEYINPUT99), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n357), .A2(new_n629), .A3(new_n236), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n248), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n517), .A2(new_n620), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n612), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n609), .B1(new_n595), .B2(new_n604), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT33), .B1(new_n611), .B2(new_n612), .ZN(new_n639));
  OAI211_X1 g453(.A(G478), .B(new_n236), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT100), .B1(new_n613), .B2(new_n614), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n637), .B1(new_n635), .B2(new_n636), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n611), .A2(KEYINPUT33), .A3(new_n612), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n614), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n642), .B1(new_n645), .B2(new_n236), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT101), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n642), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n640), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n650), .A3(new_n236), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n647), .A2(new_n653), .A3(new_n561), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n453), .A2(new_n465), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n571), .A2(new_n472), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n634), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT34), .B(G104), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  AND4_X1   g474(.A1(new_n616), .A2(new_n547), .A3(new_n559), .A4(new_n560), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n655), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n634), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT35), .B(G107), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  OR3_X1    g480(.A1(new_n217), .A2(new_n231), .A3(KEYINPUT36), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n217), .B1(new_n231), .B2(KEYINPUT36), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n238), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n246), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n246), .A2(KEYINPUT102), .A3(new_n669), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n631), .A2(new_n473), .A3(new_n621), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT37), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(G110), .Z(G12));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n362), .B2(new_n384), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n386), .B1(new_n463), .B2(new_n464), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n471), .B1(new_n680), .B2(new_n467), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n547), .A2(new_n559), .A3(new_n560), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n564), .B1(new_n567), .B2(G900), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n616), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT103), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n472), .B1(new_n453), .B2(new_n465), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n661), .A4(new_n683), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n679), .A2(new_n689), .A3(new_n633), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XNOR2_X1  g505(.A(new_n683), .B(KEYINPUT39), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n633), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n674), .B1(new_n693), .B2(KEYINPUT40), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT32), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n624), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n698));
  INV_X1    g512(.A(new_n336), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n326), .A2(new_n335), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(G902), .B1(new_n701), .B2(new_n342), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n342), .B1(new_n334), .B2(new_n336), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n697), .A2(new_n698), .A3(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n561), .A2(new_n616), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n706), .A2(new_n471), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT38), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n470), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n466), .A2(KEYINPUT38), .A3(new_n469), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n694), .A2(new_n695), .A3(new_n708), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  NAND2_X1  g528(.A1(new_n517), .A2(new_n620), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n681), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n383), .A2(new_n365), .A3(G902), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n697), .B(new_n698), .C1(new_n717), .C2(new_n626), .ZN(new_n718));
  AND4_X1   g532(.A1(new_n561), .A2(new_n647), .A3(new_n653), .A4(new_n683), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n718), .A3(new_n674), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  NOR2_X1   g535(.A1(new_n657), .A2(new_n654), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n503), .A2(new_n497), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n723), .A2(new_n509), .B1(new_n513), .B2(new_n490), .ZN(new_n724));
  OAI21_X1  g538(.A(G469), .B1(new_n724), .B2(G902), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n620), .A3(new_n505), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n718), .A2(new_n722), .A3(new_n632), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT104), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n728), .B(new_n730), .ZN(G15));
  NAND4_X1  g545(.A1(new_n718), .A2(new_n662), .A3(new_n632), .A4(new_n727), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NOR2_X1   g547(.A1(new_n726), .A2(new_n681), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n718), .A2(new_n617), .A3(new_n734), .A4(new_n674), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT105), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n679), .A2(new_n737), .A3(new_n617), .A4(new_n734), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  OAI211_X1 g554(.A(new_n346), .B(new_n356), .C1(new_n343), .C2(new_n380), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(new_n359), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n626), .B1(new_n357), .B2(new_n236), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n742), .A2(new_n743), .A3(new_n248), .ZN(new_n744));
  INV_X1    g558(.A(new_n657), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n707), .A4(new_n727), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NOR3_X1   g561(.A1(new_n678), .A2(new_n742), .A3(new_n743), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n719), .A3(new_n734), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NAND2_X1  g564(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n472), .B1(new_n466), .B2(new_n469), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n718), .A2(new_n632), .A3(new_n633), .A4(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n719), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n752), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n715), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n757), .A2(new_n385), .A3(new_n719), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NOR2_X1   g576(.A1(new_n753), .A2(new_n684), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n267), .ZN(G36));
  NAND2_X1  g578(.A1(new_n508), .A2(new_n509), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n513), .A2(new_n503), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT45), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT107), .B1(new_n767), .B2(new_n474), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n514), .A2(KEYINPUT45), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n770), .B(G469), .C1(new_n514), .C2(KEYINPUT45), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n516), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n516), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n505), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(G472), .A3(new_n630), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n624), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n682), .A2(new_n647), .A3(new_n653), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n682), .A2(new_n647), .A3(new_n653), .A4(KEYINPUT43), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n780), .A2(KEYINPUT44), .A3(new_n674), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n777), .A2(new_n620), .A3(new_n786), .A4(new_n692), .ZN(new_n787));
  INV_X1    g601(.A(new_n630), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n629), .B1(new_n357), .B2(new_n236), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n788), .A2(new_n789), .A3(new_n626), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n785), .B(new_n674), .C1(new_n790), .C2(new_n625), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n752), .B(KEYINPUT108), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT109), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NAND2_X1  g612(.A1(new_n777), .A2(new_n620), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n718), .A2(new_n632), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n777), .A2(new_n802), .A3(new_n620), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n756), .A2(new_n754), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n800), .A2(new_n801), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n807));
  INV_X1    g621(.A(new_n670), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n655), .A2(new_n808), .A3(new_n683), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n715), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n471), .A3(new_n707), .A4(new_n706), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n690), .A2(new_n720), .A3(new_n749), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n715), .B1(new_n685), .B2(new_n688), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n627), .A2(G472), .B1(new_n359), .B2(new_n741), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n674), .A2(new_n816), .A3(new_n719), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n815), .A2(new_n679), .B1(new_n817), .B2(new_n734), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(KEYINPUT52), .A3(new_n720), .A4(new_n811), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n728), .A2(new_n732), .A3(new_n746), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n738), .B2(new_n736), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n718), .A2(new_n633), .A3(new_n674), .A4(new_n752), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n561), .A2(new_n616), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n683), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT111), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  INV_X1    g642(.A(new_n826), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n757), .A2(new_n679), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n763), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n649), .A2(new_n652), .A3(new_n651), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n652), .B1(new_n649), .B2(new_n651), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n661), .B1(new_n834), .B2(new_n561), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n466), .A2(new_n469), .A3(new_n656), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n632), .A3(new_n631), .A4(new_n633), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n748), .A2(new_n633), .A3(new_n719), .A4(new_n752), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n622), .A2(new_n838), .A3(new_n675), .A4(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n823), .A2(new_n831), .A3(new_n840), .A4(new_n761), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n807), .B1(new_n821), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n761), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n728), .A2(new_n732), .A3(new_n746), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n739), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT112), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n807), .B1(new_n814), .B2(new_n819), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n831), .A2(new_n840), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n823), .A2(new_n849), .A3(new_n761), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n842), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT113), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n842), .A2(new_n851), .A3(new_n855), .A4(new_n852), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n843), .A2(new_n845), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n848), .A2(new_n859), .A3(KEYINPUT53), .A4(new_n820), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n842), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n710), .A2(new_n472), .A3(new_n711), .A4(new_n727), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n864), .A2(KEYINPUT115), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n564), .B1(new_n783), .B2(new_n784), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n744), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(KEYINPUT115), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(KEYINPUT50), .A3(new_n867), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n756), .A2(new_n726), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n866), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n874), .B2(new_n866), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n748), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n706), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n879), .A3(new_n632), .A4(new_n565), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n561), .A3(new_n834), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n873), .A2(new_n878), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n867), .A2(new_n794), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n800), .A2(new_n803), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n725), .A2(new_n619), .A3(new_n505), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT114), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n863), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n886), .ZN(new_n890));
  INV_X1    g704(.A(new_n884), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n881), .B1(new_n871), .B2(new_n872), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(KEYINPUT51), .A3(new_n878), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n867), .A2(new_n734), .ZN(new_n895));
  OAI211_X1 g709(.A(G952), .B(new_n563), .C1(new_n880), .C2(new_n654), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n385), .B1(new_n876), .B2(new_n877), .ZN(new_n897));
  OR2_X1    g711(.A1(new_n897), .A2(KEYINPUT48), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(KEYINPUT48), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n889), .A2(new_n894), .A3(new_n895), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n857), .A2(new_n858), .A3(new_n862), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n854), .A2(new_n862), .A3(new_n856), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT117), .B1(new_n904), .B2(new_n901), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT118), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n725), .A2(new_n505), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT49), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n712), .A2(new_n910), .A3(new_n781), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n248), .A2(new_n472), .A3(new_n619), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT110), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n879), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n908), .A2(new_n914), .ZN(G75));
  AOI21_X1  g729(.A(new_n236), .B1(new_n842), .B2(new_n851), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n916), .B2(G210), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n461), .B(KEYINPUT119), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n393), .B(KEYINPUT55), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(KEYINPUT120), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n917), .B(new_n922), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n219), .A2(G952), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G51));
  NAND2_X1  g739(.A1(new_n842), .A2(new_n851), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n853), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n516), .B(KEYINPUT57), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n929), .A2(new_n930), .B1(new_n504), .B2(new_n501), .ZN(new_n931));
  INV_X1    g745(.A(new_n772), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n916), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n924), .B1(new_n931), .B2(new_n933), .ZN(G54));
  INV_X1    g748(.A(new_n924), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n544), .A2(new_n556), .ZN(new_n938));
  OR3_X1    g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n937), .B1(new_n936), .B2(new_n938), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n935), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(G60));
  NAND2_X1  g756(.A1(new_n643), .A2(new_n644), .ZN(new_n943));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT59), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n842), .A2(new_n851), .A3(new_n852), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n852), .B1(new_n842), .B2(new_n851), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n943), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT122), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n928), .A2(new_n950), .A3(new_n943), .A4(new_n945), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n904), .A2(new_n945), .ZN(new_n953));
  INV_X1    g767(.A(new_n943), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n952), .A2(new_n955), .A3(new_n935), .ZN(G63));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT123), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n842), .B2(new_n851), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n667), .A3(new_n668), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n935), .C1(new_n234), .C2(new_n960), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G66));
  OAI21_X1  g778(.A(G953), .B1(new_n570), .B2(new_n391), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n838), .A2(new_n622), .A3(new_n675), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n845), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n967), .B2(new_n566), .ZN(new_n968));
  INV_X1    g782(.A(G898), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n918), .B1(new_n969), .B2(new_n566), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n968), .B(new_n970), .Z(G69));
  AND3_X1   g785(.A1(new_n690), .A2(new_n720), .A3(new_n749), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n713), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT62), .Z(new_n974));
  INV_X1    g788(.A(new_n796), .ZN(new_n975));
  INV_X1    g789(.A(new_n693), .ZN(new_n976));
  INV_X1    g790(.A(new_n835), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n976), .A2(new_n385), .A3(new_n752), .A4(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n974), .A2(new_n975), .A3(new_n805), .A4(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n327), .A2(new_n333), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n301), .B2(new_n300), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(new_n553), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n777), .A2(new_n620), .A3(new_n692), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n385), .A3(new_n686), .A4(new_n707), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n763), .B1(new_n755), .B2(new_n760), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n805), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n972), .B1(new_n787), .B2(new_n795), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT124), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n992), .B(new_n972), .C1(new_n787), .C2(new_n795), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n988), .A2(new_n989), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n993), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n805), .A2(new_n986), .A3(new_n987), .ZN(new_n996));
  OAI21_X1  g810(.A(KEYINPUT125), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(new_n997), .A3(new_n982), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n984), .A2(new_n998), .A3(new_n219), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n219), .B1(new_n982), .B2(G227), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n1000), .B(G900), .C1(G227), .C2(new_n982), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n999), .A2(new_n1001), .ZN(G72));
  NAND3_X1  g816(.A1(new_n994), .A2(new_n997), .A3(new_n967), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n364), .B(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(KEYINPUT127), .A3(new_n935), .ZN(new_n1009));
  INV_X1    g823(.A(new_n967), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n979), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n704), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n861), .A2(new_n364), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n1011), .A2(new_n704), .B1(new_n1013), .B2(new_n1005), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1007), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1015), .B1(new_n1017), .B2(new_n924), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1009), .A2(new_n1014), .A3(new_n1018), .ZN(G57));
endmodule


