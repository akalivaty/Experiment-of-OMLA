//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970;
  AND2_X1   g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n206), .A2(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n210), .A2(KEYINPUT69), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT69), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n208), .B(new_n213), .C1(new_n207), .C2(new_n206), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT27), .B(G183gat), .Z(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT67), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220));
  AOI21_X1  g019(.A(G190gat), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT28), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n216), .A2(new_n223), .A3(G190gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n214), .B(new_n215), .C1(new_n222), .C2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n227));
  OAI211_X1 g026(.A(KEYINPUT23), .B(new_n203), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT24), .A3(new_n215), .ZN(new_n230));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT23), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n205), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n215), .A2(KEYINPUT24), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n228), .A2(new_n230), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n236), .B1(new_n209), .B2(KEYINPUT23), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n242), .A2(new_n230), .A3(new_n234), .A4(new_n233), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT66), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n239), .B1(new_n235), .B2(new_n236), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT66), .B(new_n243), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n202), .B(new_n225), .C1(new_n244), .C2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G197gat), .B(G204gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT22), .ZN(new_n251));
  INV_X1    g050(.A(G211gat), .ZN(new_n252));
  INV_X1    g051(.A(G218gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT76), .ZN(new_n258));
  INV_X1    g057(.A(new_n256), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n255), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT76), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n225), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n202), .A2(KEYINPUT29), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n202), .A3(new_n225), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n225), .B1(new_n244), .B2(new_n248), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(new_n266), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n268), .B1(new_n272), .B2(new_n263), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT37), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(G8gat), .B(G36gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G64gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(G92gat), .Z(new_n278));
  INV_X1    g077(.A(new_n225), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n281), .B2(new_n247), .ZN(new_n282));
  INV_X1    g081(.A(new_n266), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n269), .B(new_n263), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n249), .A2(new_n267), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n284), .B(KEYINPUT37), .C1(new_n285), .C2(new_n263), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT38), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n269), .B1(new_n282), .B2(new_n283), .ZN(new_n290));
  INV_X1    g089(.A(new_n263), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT37), .A3(new_n268), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n275), .A2(KEYINPUT38), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G148gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G141gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT79), .B(G141gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n299), .B2(new_n296), .ZN(new_n300));
  XOR2_X1   g099(.A(G155gat), .B(G162gat), .Z(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT2), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  INV_X1    g107(.A(G141gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G148gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n296), .A2(G141gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(G148gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n313), .A3(KEYINPUT77), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n304), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n315), .A2(new_n316), .A3(new_n301), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n316), .B1(new_n315), .B2(new_n301), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n307), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g119(.A(G127gat), .ZN(new_n321));
  INV_X1    g120(.A(G134gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G127gat), .A2(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G113gat), .ZN(new_n328));
  INV_X1    g127(.A(G113gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G120gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n325), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT70), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n329), .B2(G120gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n327), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n330), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(new_n326), .A3(new_n325), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT71), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n336), .A2(new_n339), .A3(new_n326), .A4(new_n325), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n332), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(new_n307), .C1(new_n317), .C2(new_n318), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n320), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n341), .B(new_n307), .C1(new_n317), .C2(new_n318), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n315), .A2(new_n301), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT78), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n315), .A2(new_n316), .A3(new_n301), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n351), .A2(new_n352), .B1(new_n300), .B2(new_n306), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n345), .A2(new_n346), .A3(new_n349), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n319), .A2(new_n342), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n346), .B1(new_n356), .B2(new_n347), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT5), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G57gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372));
  INV_X1    g171(.A(new_n370), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n362), .A2(new_n365), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n278), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n273), .B2(KEYINPUT38), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n357), .A2(new_n358), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(KEYINPUT5), .A3(new_n359), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n364), .B1(new_n379), .B2(new_n355), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT6), .A4(new_n373), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n362), .A2(new_n365), .A3(KEYINPUT6), .A4(new_n373), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT84), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n295), .A2(new_n375), .A3(new_n377), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n344), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT3), .B1(new_n260), .B2(new_n387), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n388), .A2(new_n291), .B1(new_n319), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT81), .B1(new_n353), .B2(new_n389), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n263), .B1(new_n387), .B2(new_n344), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n353), .A2(new_n389), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n393), .B(new_n392), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n398), .A3(KEYINPUT82), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G22gat), .ZN(new_n400));
  INV_X1    g199(.A(G22gat), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n395), .A2(new_n398), .A3(KEYINPUT82), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n398), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(G78gat), .B(G106gat), .Z(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n400), .A2(new_n406), .A3(new_n409), .A4(new_n402), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n273), .A2(KEYINPUT30), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n292), .A2(new_n416), .A3(new_n268), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n417), .A3(new_n376), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n273), .A2(KEYINPUT30), .A3(new_n278), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n345), .A2(new_n349), .A3(new_n354), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(G225gat), .A3(G233gat), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(KEYINPUT39), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n356), .A2(new_n346), .A3(new_n347), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(KEYINPUT39), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n370), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT40), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n424), .A2(KEYINPUT40), .A3(new_n370), .A4(new_n426), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n421), .A2(new_n429), .A3(new_n374), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n386), .A2(new_n414), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n414), .A2(KEYINPUT83), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n375), .A2(new_n383), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n433), .B(new_n435), .C1(new_n437), .C2(new_n421), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  NAND2_X1  g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n271), .A2(new_n342), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n341), .B(new_n225), .C1(new_n244), .C2(new_n248), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n446), .B2(KEYINPUT33), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT32), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n443), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n282), .A2(new_n341), .ZN(new_n452));
  AOI211_X1 g251(.A(new_n342), .B(new_n279), .C1(new_n281), .C2(new_n247), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  INV_X1    g254(.A(new_n442), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n454), .B(KEYINPUT32), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT75), .B1(new_n450), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT74), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n444), .A2(KEYINPUT73), .A3(new_n443), .A4(new_n445), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT72), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n451), .A2(KEYINPUT73), .B1(KEYINPUT72), .B2(KEYINPUT34), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n452), .A2(new_n453), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n443), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n460), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n462), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT34), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n445), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n465), .B1(new_n472), .B2(new_n451), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(KEYINPUT74), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n454), .A2(KEYINPUT32), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n455), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n442), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n457), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT74), .B1(new_n471), .B2(new_n473), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n464), .A2(new_n468), .A3(new_n460), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT75), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n439), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n474), .A2(new_n469), .A3(new_n457), .A4(new_n478), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n484), .A2(new_n439), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n432), .B(new_n438), .C1(new_n483), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n485), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n413), .B1(new_n385), .B2(new_n375), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n420), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI211_X1 g291(.A(new_n491), .B(new_n413), .C1(new_n475), .C2(new_n482), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n437), .A2(new_n421), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n487), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497));
  INV_X1    g296(.A(G43gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G50gat), .ZN(new_n499));
  INV_X1    g298(.A(G50gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G43gat), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT15), .ZN(new_n502));
  INV_X1    g301(.A(G29gat), .ZN(new_n503));
  INV_X1    g302(.A(G36gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT14), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(G29gat), .A2(G36gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n502), .A2(KEYINPUT87), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT87), .B1(new_n502), .B2(new_n509), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(KEYINPUT88), .A2(G50gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n498), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT15), .B1(new_n515), .B2(new_n501), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n516), .A2(new_n502), .A3(new_n509), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT89), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT87), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT15), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT87), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n515), .A2(new_n501), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n521), .B(new_n520), .C1(new_n525), .C2(KEYINPUT15), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT17), .B1(new_n518), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n532), .A2(G1gat), .ZN(new_n537));
  OAI211_X1 g336(.A(KEYINPUT90), .B(new_n531), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n531), .A2(KEYINPUT90), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n531), .A2(KEYINPUT90), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n539), .A2(new_n535), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n530), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n497), .B1(new_n529), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n512), .A2(new_n517), .A3(KEYINPUT89), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n527), .B1(new_n524), .B2(new_n526), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n544), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(KEYINPUT91), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n518), .A2(new_n528), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n538), .A3(new_n542), .ZN(new_n553));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n545), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT18), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n552), .B(new_n543), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n554), .B(KEYINPUT13), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G169gat), .B(G197gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n570));
  XOR2_X1   g369(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n561), .A3(new_n563), .A4(new_n571), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n572), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(KEYINPUT94), .A3(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n584), .B(KEYINPUT96), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT97), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  XOR2_X1   g390(.A(G57gat), .B(G64gat), .Z(new_n592));
  NAND4_X1  g391(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n543), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n218), .ZN(new_n600));
  AND2_X1   g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n597), .A2(new_n598), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  XOR2_X1   g407(.A(new_n605), .B(new_n608), .Z(new_n609));
  NAND2_X1  g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT7), .ZN(new_n611));
  INV_X1    g410(.A(G99gat), .ZN(new_n612));
  INV_X1    g411(.A(G106gat), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT8), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n611), .B(new_n614), .C1(G85gat), .C2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT98), .Z(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(new_n529), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n530), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n618), .A2(new_n552), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n593), .A4(new_n596), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n597), .B(new_n617), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n637), .A2(new_n634), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n204), .ZN(new_n644));
  INV_X1    g443(.A(G204gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n633), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  NOR4_X1   g447(.A1(new_n640), .A2(KEYINPUT99), .A3(new_n641), .A4(new_n646), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n646), .B1(new_n640), .B2(new_n641), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n609), .A2(new_n632), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n583), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n496), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n436), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n533), .ZN(G1324gat));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n420), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT42), .Z(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n531), .B2(new_n659), .ZN(G1325gat));
  NOR2_X1   g462(.A1(new_n483), .A2(new_n486), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n656), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n656), .A2(G15gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n488), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT100), .Z(G1326gat));
  NAND2_X1  g469(.A1(new_n433), .A2(new_n435), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT101), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n672), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n578), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n576), .A2(KEYINPUT102), .A3(new_n577), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n653), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n609), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n496), .A2(new_n632), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT104), .B1(new_n685), .B2(KEYINPUT44), .ZN(new_n686));
  INV_X1    g485(.A(new_n632), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n493), .A2(new_n494), .B1(new_n491), .B2(new_n490), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n487), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n685), .A2(new_n694), .A3(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT103), .B1(new_n689), .B2(new_n691), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n684), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n436), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n685), .A2(new_n582), .A3(new_n682), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n503), .A3(new_n437), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(G1328gat));
  OAI21_X1  g503(.A(G36gat), .B1(new_n699), .B2(new_n420), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n701), .A2(new_n504), .A3(new_n421), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT46), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(new_n701), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G43gat), .A3(new_n668), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n694), .B1(new_n685), .B2(KEYINPUT44), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n689), .A2(KEYINPUT103), .A3(new_n691), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n690), .A2(new_n496), .A3(new_n691), .A4(new_n632), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n690), .B1(new_n689), .B2(new_n691), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n711), .A2(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n664), .A3(new_n683), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n710), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT106), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n498), .B1(new_n698), .B2(new_n664), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT105), .B(new_n720), .C1(new_n721), .C2(new_n710), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT47), .B1(new_n719), .B2(new_n722), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n513), .A2(new_n514), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n671), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n698), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n671), .A2(new_n727), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT107), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n709), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n726), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n728), .B1(new_n698), .B2(new_n413), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT48), .B1(new_n709), .B2(new_n732), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(KEYINPUT109), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n736), .B(new_n737), .C1(new_n741), .C2(new_n742), .ZN(G1331gat));
  AOI211_X1 g542(.A(new_n609), .B(new_n632), .C1(new_n688), .C2(new_n487), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n679), .A2(new_n681), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n436), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT110), .B(G57gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  NOR2_X1   g548(.A1(new_n746), .A2(new_n420), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n746), .B2(new_n665), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n746), .A2(G71gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(new_n668), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT111), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g558(.A1(new_n746), .A2(new_n671), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(G78gat), .Z(G1335gat));
  NAND3_X1  g560(.A1(new_n715), .A2(new_n609), .A3(new_n745), .ZN(new_n762));
  INV_X1    g561(.A(G85gat), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n762), .A2(new_n763), .A3(new_n436), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n689), .A2(new_n609), .A3(new_n680), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(new_n653), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n437), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n764), .B1(new_n763), .B2(new_n770), .ZN(G1336gat));
  NAND4_X1  g570(.A1(new_n715), .A2(new_n421), .A3(new_n609), .A4(new_n745), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n681), .A2(G92gat), .A3(new_n420), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT112), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT52), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n772), .B2(new_n779), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(G1337gat));
  NOR3_X1   g583(.A1(new_n762), .A2(new_n612), .A3(new_n665), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n488), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n612), .B2(new_n786), .ZN(G1338gat));
  OAI21_X1  g586(.A(G106gat), .B1(new_n762), .B2(new_n671), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n768), .A2(new_n613), .A3(new_n653), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n414), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n789), .A2(KEYINPUT115), .A3(new_n414), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT115), .B1(new_n789), .B2(new_n414), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n715), .A2(new_n413), .A3(new_n609), .A4(new_n745), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G106gat), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n791), .B1(new_n794), .B2(new_n800), .ZN(G1339gat));
  NAND2_X1  g600(.A1(new_n680), .A2(new_n654), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n640), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n636), .A2(new_n639), .A3(new_n635), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT54), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n805), .B(new_n646), .C1(new_n807), .C2(new_n640), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n649), .A2(new_n648), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(KEYINPUT117), .A3(new_n809), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n559), .A2(new_n560), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT118), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n545), .A2(new_n551), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n554), .B1(new_n818), .B2(new_n553), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n569), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n575), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n815), .A2(new_n632), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n679), .A2(new_n815), .B1(new_n653), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n632), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n803), .B1(new_n824), .B2(new_n609), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n436), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n413), .B1(new_n475), .B2(new_n482), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n826), .A2(new_n420), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n329), .A3(new_n679), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n576), .A2(KEYINPUT102), .A3(new_n577), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT102), .B1(new_n576), .B2(new_n577), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n815), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n653), .A2(new_n821), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n632), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n822), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n609), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n802), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n729), .A2(new_n668), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n436), .A2(new_n421), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n582), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n844), .ZN(G1340gat));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n327), .A3(new_n653), .ZN(new_n846));
  OAI21_X1  g645(.A(G120gat), .B1(new_n843), .B2(new_n681), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1341gat));
  INV_X1    g647(.A(new_n609), .ZN(new_n849));
  AOI21_X1  g648(.A(G127gat), .B1(new_n828), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n609), .A2(new_n321), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n842), .B2(new_n851), .ZN(G1342gat));
  NAND3_X1  g651(.A1(new_n828), .A2(new_n322), .A3(new_n632), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT56), .Z(new_n854));
  OAI21_X1  g653(.A(G134gat), .B1(new_n843), .B2(new_n687), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n826), .A2(KEYINPUT120), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n664), .A2(new_n414), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n826), .B2(KEYINPUT120), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT121), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n826), .A2(KEYINPUT120), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n863), .A2(new_n864), .A3(new_n858), .A4(new_n860), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n865), .A3(new_n420), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n582), .A2(G141gat), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n857), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n810), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n580), .A2(new_n581), .A3(new_n870), .A4(new_n811), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n632), .B1(new_n871), .B2(new_n833), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n609), .B1(new_n872), .B2(new_n835), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT119), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n803), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n671), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n825), .A2(KEYINPUT57), .A3(new_n414), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(new_n664), .A3(new_n841), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n298), .B1(new_n883), .B2(new_n583), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n679), .A3(new_n882), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n859), .A2(new_n861), .A3(new_n421), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n885), .A2(new_n299), .B1(new_n886), .B2(new_n867), .ZN(new_n887));
  OAI22_X1  g686(.A1(new_n869), .A2(new_n884), .B1(new_n857), .B2(new_n887), .ZN(G1344gat));
  OAI21_X1  g687(.A(KEYINPUT57), .B1(new_n825), .B2(new_n414), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n654), .A2(new_n582), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n879), .B(new_n729), .C1(new_n874), .C2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n664), .A2(new_n841), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n653), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g696(.A(G148gat), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT59), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n882), .B(new_n653), .C1(new_n879), .C2(new_n878), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n296), .A2(KEYINPUT59), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(KEYINPUT122), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT122), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n866), .A2(G148gat), .A3(new_n681), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1345gat));
  OR2_X1    g705(.A1(new_n866), .A2(new_n609), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n609), .A2(new_n302), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n907), .A2(new_n302), .B1(new_n883), .B2(new_n908), .ZN(G1346gat));
  OAI21_X1  g708(.A(new_n303), .B1(new_n866), .B2(new_n687), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n883), .A2(G162gat), .A3(new_n632), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n437), .A2(new_n420), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n839), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n582), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT124), .B1(new_n825), .B2(new_n437), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n837), .A2(new_n919), .A3(new_n436), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n827), .A2(new_n421), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n679), .A2(new_n203), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n917), .B1(new_n923), .B2(new_n924), .ZN(G1348gat));
  NAND3_X1  g724(.A1(new_n921), .A2(new_n653), .A3(new_n922), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n681), .A2(new_n227), .A3(new_n226), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n926), .A2(new_n204), .B1(new_n915), .B2(new_n927), .ZN(G1349gat));
  NOR2_X1   g727(.A1(new_n609), .A2(new_n216), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n919), .B1(new_n837), .B2(new_n436), .ZN(new_n930));
  AOI211_X1 g729(.A(KEYINPUT124), .B(new_n437), .C1(new_n836), .C2(new_n802), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n922), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n921), .A2(KEYINPUT125), .A3(new_n922), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n218), .B1(new_n915), .B2(new_n849), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT126), .B1(new_n939), .B2(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n934), .B2(new_n935), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n941), .A2(KEYINPUT127), .A3(new_n943), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT127), .B1(new_n941), .B2(new_n943), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n940), .A2(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n916), .B2(new_n687), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT61), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n687), .A2(G190gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n923), .B2(new_n950), .ZN(G1351gat));
  AND3_X1   g750(.A1(new_n921), .A2(new_n421), .A3(new_n860), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n679), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n664), .A2(new_n914), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n892), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G197gat), .B1(new_n956), .B2(new_n582), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n957), .ZN(G1352gat));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n645), .A3(new_n653), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n892), .A2(new_n653), .A3(new_n955), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n960), .B(new_n961), .C1(new_n645), .C2(new_n962), .ZN(G1353gat));
  NAND3_X1  g762(.A1(new_n952), .A2(new_n252), .A3(new_n849), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n892), .A2(new_n849), .A3(new_n955), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  NAND3_X1  g767(.A1(new_n952), .A2(new_n253), .A3(new_n632), .ZN(new_n969));
  OAI21_X1  g768(.A(G218gat), .B1(new_n956), .B2(new_n687), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1355gat));
endmodule


