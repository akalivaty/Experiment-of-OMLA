

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742;

  XNOR2_X1 U369 ( .A(n527), .B(n354), .ZN(n367) );
  BUF_X1 U370 ( .A(G104), .Z(n347) );
  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n532) );
  OR2_X2 U372 ( .A1(n661), .A2(n369), .ZN(n440) );
  OR2_X4 U373 ( .A1(n396), .A2(n459), .ZN(n383) );
  AND2_X4 U374 ( .A1(n348), .A2(n383), .ZN(n709) );
  NAND2_X2 U375 ( .A1(n479), .A2(n478), .ZN(n445) );
  XNOR2_X1 U376 ( .A(G128), .B(G110), .ZN(n467) );
  XNOR2_X1 U377 ( .A(G116), .B(G107), .ZN(n519) );
  INV_X1 U378 ( .A(G953), .ZN(n728) );
  AND2_X2 U379 ( .A1(n377), .A2(n375), .ZN(n374) );
  NOR2_X1 U380 ( .A1(n560), .A2(KEYINPUT44), .ZN(n413) );
  XNOR2_X1 U381 ( .A(n447), .B(KEYINPUT102), .ZN(n401) );
  XNOR2_X1 U382 ( .A(n540), .B(KEYINPUT31), .ZN(n650) );
  NAND2_X1 U383 ( .A1(n408), .A2(n671), .ZN(n540) );
  NOR2_X1 U384 ( .A1(n554), .A2(n350), .ZN(n432) );
  XNOR2_X1 U385 ( .A(KEYINPUT73), .B(G122), .ZN(n458) );
  NAND2_X1 U386 ( .A1(n373), .A2(n699), .ZN(n372) );
  NOR2_X1 U387 ( .A1(n631), .A2(n713), .ZN(n633) );
  NOR2_X1 U388 ( .A1(n626), .A2(n713), .ZN(n627) );
  INV_X1 U389 ( .A(n691), .ZN(n348) );
  XNOR2_X1 U390 ( .A(n413), .B(KEYINPUT71), .ZN(n412) );
  NAND2_X1 U391 ( .A1(n389), .A2(n388), .ZN(n727) );
  NOR2_X1 U392 ( .A1(n432), .A2(n430), .ZN(n429) );
  AND2_X1 U393 ( .A1(n543), .A2(n537), .ZN(n353) );
  OR2_X1 U394 ( .A1(n711), .A2(G902), .ZN(n451) );
  XNOR2_X1 U395 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U396 ( .A(n452), .B(n468), .ZN(n711) );
  XNOR2_X1 U397 ( .A(n469), .B(n472), .ZN(n452) );
  XNOR2_X1 U398 ( .A(n391), .B(n390), .ZN(n531) );
  XNOR2_X1 U399 ( .A(n422), .B(n466), .ZN(n469) );
  XNOR2_X1 U400 ( .A(n467), .B(n465), .ZN(n422) );
  XNOR2_X1 U401 ( .A(n458), .B(KEYINPUT16), .ZN(n443) );
  XOR2_X1 U402 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n465) );
  INV_X1 U403 ( .A(G104), .ZN(n477) );
  AND2_X2 U404 ( .A1(n368), .A2(n619), .ZN(n402) );
  XNOR2_X2 U405 ( .A(n495), .B(n355), .ZN(n427) );
  XNOR2_X2 U406 ( .A(n400), .B(n621), .ZN(n691) );
  OR2_X1 U407 ( .A1(G237), .A2(G902), .ZN(n496) );
  XOR2_X1 U408 ( .A(G137), .B(KEYINPUT4), .Z(n475) );
  NOR2_X1 U409 ( .A1(n727), .A2(n399), .ZN(n398) );
  NOR2_X1 U410 ( .A1(n541), .A2(n680), .ZN(n424) );
  NOR2_X1 U411 ( .A1(n638), .A2(n650), .ZN(n541) );
  XNOR2_X1 U412 ( .A(n727), .B(KEYINPUT75), .ZN(n397) );
  XNOR2_X1 U413 ( .A(n367), .B(KEYINPUT89), .ZN(n723) );
  XNOR2_X1 U414 ( .A(n454), .B(G125), .ZN(n487) );
  INV_X1 U415 ( .A(G146), .ZN(n454) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(KEYINPUT77), .ZN(n456) );
  XNOR2_X1 U417 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n486) );
  XNOR2_X1 U418 ( .A(n617), .B(KEYINPUT83), .ZN(n425) );
  NOR2_X1 U419 ( .A1(n575), .A2(n567), .ZN(n583) );
  INV_X1 U420 ( .A(KEYINPUT92), .ZN(n438) );
  XNOR2_X1 U421 ( .A(n666), .B(n352), .ZN(n568) );
  XNOR2_X1 U422 ( .A(n392), .B(n531), .ZN(n534) );
  XNOR2_X1 U423 ( .A(n393), .B(n530), .ZN(n392) );
  XNOR2_X1 U424 ( .A(n613), .B(n612), .ZN(n618) );
  NOR2_X1 U425 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U426 ( .A1(n431), .A2(n359), .ZN(n430) );
  INV_X1 U427 ( .A(n727), .ZN(n387) );
  INV_X1 U428 ( .A(KEYINPUT69), .ZN(n450) );
  XNOR2_X1 U429 ( .A(n533), .B(n394), .ZN(n393) );
  XNOR2_X1 U430 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n394) );
  XNOR2_X1 U431 ( .A(G137), .B(G119), .ZN(n464) );
  XOR2_X1 U432 ( .A(KEYINPUT68), .B(G131), .Z(n506) );
  NAND2_X1 U433 ( .A1(G234), .A2(G237), .ZN(n497) );
  NOR2_X1 U434 ( .A1(n353), .A2(n649), .ZN(n680) );
  XNOR2_X1 U435 ( .A(G119), .B(G113), .ZN(n390) );
  XNOR2_X1 U436 ( .A(n441), .B(G116), .ZN(n391) );
  INV_X1 U437 ( .A(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U438 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n470) );
  XNOR2_X1 U439 ( .A(n487), .B(n453), .ZN(n724) );
  XNOR2_X1 U440 ( .A(G140), .B(KEYINPUT10), .ZN(n453) );
  XNOR2_X1 U441 ( .A(G113), .B(G122), .ZN(n508) );
  XOR2_X1 U442 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n509) );
  XOR2_X1 U443 ( .A(G146), .B(G140), .Z(n481) );
  XNOR2_X1 U444 ( .A(n490), .B(n491), .ZN(n493) );
  XNOR2_X1 U445 ( .A(n486), .B(n456), .ZN(n455) );
  AND2_X1 U446 ( .A1(n426), .A2(n654), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n419), .B(n448), .ZN(n389) );
  INV_X1 U448 ( .A(KEYINPUT33), .ZN(n439) );
  INV_X1 U449 ( .A(n595), .ZN(n593) );
  NAND2_X1 U450 ( .A1(n395), .A2(n353), .ZN(n595) );
  AND2_X1 U451 ( .A1(n583), .A2(n568), .ZN(n395) );
  INV_X1 U452 ( .A(KEYINPUT101), .ZN(n433) );
  INV_X1 U453 ( .A(KEYINPUT94), .ZN(n435) );
  NOR2_X1 U454 ( .A1(n376), .A2(n713), .ZN(n375) );
  NAND2_X1 U455 ( .A1(n709), .A2(n365), .ZN(n377) );
  NOR2_X1 U456 ( .A1(n423), .A2(G210), .ZN(n376) );
  XNOR2_X1 U457 ( .A(n615), .B(n614), .ZN(n742) );
  AND2_X1 U458 ( .A1(n353), .A2(n618), .ZN(n614) );
  XNOR2_X1 U459 ( .A(n410), .B(KEYINPUT35), .ZN(n737) );
  AND2_X1 U460 ( .A1(n421), .A2(n420), .ZN(n581) );
  INV_X1 U461 ( .A(n580), .ZN(n420) );
  NAND2_X1 U462 ( .A1(n349), .A2(n348), .ZN(n366) );
  OR2_X1 U463 ( .A1(KEYINPUT2), .A2(n692), .ZN(n349) );
  OR2_X1 U464 ( .A1(n599), .A2(n433), .ZN(n350) );
  NOR2_X1 U465 ( .A1(n693), .A2(n361), .ZN(n351) );
  XOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT99), .Z(n352) );
  XNOR2_X1 U467 ( .A(n506), .B(n475), .ZN(n354) );
  AND2_X1 U468 ( .A1(G210), .A2(n496), .ZN(n355) );
  NOR2_X1 U469 ( .A1(n658), .A2(n678), .ZN(n356) );
  XOR2_X1 U470 ( .A(n616), .B(n425), .Z(n357) );
  XNOR2_X1 U471 ( .A(n585), .B(KEYINPUT28), .ZN(n358) );
  AND2_X1 U472 ( .A1(n657), .A2(n666), .ZN(n359) );
  INV_X1 U473 ( .A(n666), .ZN(n584) );
  INV_X1 U474 ( .A(n426), .ZN(n655) );
  XOR2_X1 U475 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n360) );
  OR2_X1 U476 ( .A1(G953), .A2(n656), .ZN(n361) );
  XOR2_X1 U477 ( .A(KEYINPUT1), .B(KEYINPUT65), .Z(n362) );
  XOR2_X1 U478 ( .A(KEYINPUT87), .B(KEYINPUT0), .Z(n363) );
  XOR2_X1 U479 ( .A(G902), .B(KEYINPUT15), .Z(n619) );
  XOR2_X1 U480 ( .A(n629), .B(n628), .Z(n364) );
  AND2_X1 U481 ( .A1(n423), .A2(G210), .ZN(n365) );
  NOR2_X1 U482 ( .A1(G952), .A2(n728), .ZN(n713) );
  NAND2_X1 U483 ( .A1(n366), .A2(n351), .ZN(n694) );
  XNOR2_X1 U484 ( .A(n367), .B(n534), .ZN(n629) );
  AND2_X1 U485 ( .A1(n368), .A2(n387), .ZN(n692) );
  NAND2_X1 U486 ( .A1(n398), .A2(n368), .ZN(n400) );
  AND2_X1 U487 ( .A1(n368), .A2(n728), .ZN(n717) );
  XNOR2_X2 U488 ( .A(n411), .B(KEYINPUT45), .ZN(n368) );
  NOR2_X1 U489 ( .A1(n661), .A2(n662), .ZN(n371) );
  NAND2_X1 U490 ( .A1(n370), .A2(n568), .ZN(n369) );
  INV_X1 U491 ( .A(n662), .ZN(n370) );
  NAND2_X1 U492 ( .A1(n371), .A2(n584), .ZN(n538) );
  NAND2_X1 U493 ( .A1(n374), .A2(n372), .ZN(n418) );
  INV_X1 U494 ( .A(n709), .ZN(n373) );
  XNOR2_X1 U495 ( .A(n529), .B(KEYINPUT22), .ZN(n378) );
  XNOR2_X1 U496 ( .A(n529), .B(KEYINPUT22), .ZN(n554) );
  BUF_X1 U497 ( .A(n638), .Z(n379) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n638) );
  XNOR2_X1 U499 ( .A(n434), .B(n493), .ZN(n380) );
  XNOR2_X1 U500 ( .A(n434), .B(n493), .ZN(n698) );
  NAND2_X1 U501 ( .A1(n599), .A2(n433), .ZN(n431) );
  BUF_X1 U502 ( .A(n427), .Z(n381) );
  NAND2_X1 U503 ( .A1(n383), .A2(n382), .ZN(n630) );
  NOR2_X1 U504 ( .A1(n691), .A2(n386), .ZN(n382) );
  NAND2_X1 U505 ( .A1(n384), .A2(n383), .ZN(n625) );
  NOR2_X1 U506 ( .A1(n691), .A2(n385), .ZN(n384) );
  INV_X1 U507 ( .A(G475), .ZN(n385) );
  INV_X1 U508 ( .A(G472), .ZN(n386) );
  AND2_X2 U509 ( .A1(n402), .A2(n397), .ZN(n396) );
  INV_X1 U510 ( .A(KEYINPUT2), .ZN(n399) );
  NAND2_X1 U511 ( .A1(n557), .A2(n401), .ZN(n560) );
  XNOR2_X1 U512 ( .A(n401), .B(G110), .ZN(G12) );
  NAND2_X1 U513 ( .A1(n405), .A2(n403), .ZN(n409) );
  NAND2_X1 U514 ( .A1(n404), .A2(n408), .ZN(n403) );
  NOR2_X1 U515 ( .A1(n683), .A2(n546), .ZN(n404) );
  NAND2_X1 U516 ( .A1(n406), .A2(n546), .ZN(n405) );
  NAND2_X1 U517 ( .A1(n407), .A2(n408), .ZN(n406) );
  INV_X1 U518 ( .A(n683), .ZN(n407) );
  INV_X1 U519 ( .A(n545), .ZN(n408) );
  NAND2_X1 U520 ( .A1(n409), .A2(n547), .ZN(n410) );
  NAND2_X1 U521 ( .A1(n414), .A2(n412), .ZN(n411) );
  XNOR2_X1 U522 ( .A(n416), .B(n415), .ZN(n414) );
  INV_X1 U523 ( .A(KEYINPUT84), .ZN(n415) );
  NAND2_X1 U524 ( .A1(n559), .A2(n558), .ZN(n416) );
  XNOR2_X1 U525 ( .A(n418), .B(n417), .ZN(G51) );
  INV_X1 U526 ( .A(KEYINPUT56), .ZN(n417) );
  NAND2_X1 U527 ( .A1(n449), .A2(n357), .ZN(n419) );
  XNOR2_X1 U528 ( .A(n573), .B(KEYINPUT30), .ZN(n574) );
  XNOR2_X1 U529 ( .A(n579), .B(KEYINPUT106), .ZN(n421) );
  INV_X1 U530 ( .A(n699), .ZN(n423) );
  NOR2_X2 U531 ( .A1(n657), .A2(n536), .ZN(n634) );
  XNOR2_X1 U532 ( .A(n457), .B(n438), .ZN(n437) );
  NOR2_X2 U533 ( .A1(n424), .A2(n634), .ZN(n542) );
  XNOR2_X2 U534 ( .A(n440), .B(n439), .ZN(n683) );
  XNOR2_X2 U535 ( .A(n586), .B(n362), .ZN(n661) );
  XNOR2_X2 U536 ( .A(n485), .B(n484), .ZN(n586) );
  NAND2_X1 U537 ( .A1(n576), .A2(n577), .ZN(n611) );
  INV_X1 U538 ( .A(n381), .ZN(n578) );
  NAND2_X1 U539 ( .A1(n427), .A2(n675), .ZN(n446) );
  XNOR2_X1 U540 ( .A(n578), .B(KEYINPUT38), .ZN(n676) );
  OR2_X1 U541 ( .A1(n572), .A2(n381), .ZN(n426) );
  NOR2_X1 U542 ( .A1(n378), .A2(n599), .ZN(n556) );
  NAND2_X1 U543 ( .A1(n429), .A2(n428), .ZN(n447) );
  NAND2_X1 U544 ( .A1(n378), .A2(n433), .ZN(n428) );
  NAND2_X1 U545 ( .A1(n434), .A2(n719), .ZN(n720) );
  XNOR2_X2 U546 ( .A(n442), .B(n531), .ZN(n434) );
  NAND2_X1 U547 ( .A1(n437), .A2(n666), .ZN(n436) );
  XNOR2_X2 U548 ( .A(n489), .B(G134), .ZN(n527) );
  XNOR2_X2 U549 ( .A(n535), .B(G472), .ZN(n666) );
  XNOR2_X2 U550 ( .A(n492), .B(n443), .ZN(n442) );
  XNOR2_X2 U551 ( .A(n445), .B(n444), .ZN(n492) );
  XNOR2_X2 U552 ( .A(G101), .B(G110), .ZN(n444) );
  XNOR2_X2 U553 ( .A(n594), .B(n360), .ZN(n582) );
  XNOR2_X2 U554 ( .A(n446), .B(KEYINPUT86), .ZN(n594) );
  INV_X1 U555 ( .A(KEYINPUT48), .ZN(n448) );
  XNOR2_X1 U556 ( .A(n604), .B(n450), .ZN(n449) );
  XNOR2_X2 U557 ( .A(n451), .B(n473), .ZN(n657) );
  XNOR2_X1 U558 ( .A(n455), .B(n487), .ZN(n491) );
  INV_X1 U559 ( .A(n539), .ZN(n545) );
  NAND2_X1 U560 ( .A1(n539), .A2(n577), .ZN(n457) );
  XNOR2_X2 U561 ( .A(n503), .B(n363), .ZN(n539) );
  XNOR2_X1 U562 ( .A(n492), .B(n482), .ZN(n483) );
  AND2_X1 U563 ( .A1(n620), .A2(KEYINPUT2), .ZN(n459) );
  NOR2_X1 U564 ( .A1(n736), .A2(n603), .ZN(n604) );
  INV_X1 U565 ( .A(KEYINPUT90), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U568 ( .A(KEYINPUT70), .B(G469), .ZN(n484) );
  INV_X1 U569 ( .A(KEYINPUT39), .ZN(n612) );
  BUF_X1 U570 ( .A(n582), .Z(n588) );
  XNOR2_X1 U571 ( .A(n630), .B(n364), .ZN(n631) );
  NOR2_X1 U572 ( .A1(n588), .A2(n607), .ZN(n645) );
  XOR2_X1 U573 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n462) );
  INV_X1 U574 ( .A(n619), .ZN(n494) );
  NAND2_X1 U575 ( .A1(n494), .A2(G234), .ZN(n460) );
  XNOR2_X1 U576 ( .A(n460), .B(KEYINPUT20), .ZN(n504) );
  NAND2_X1 U577 ( .A1(n504), .A2(G217), .ZN(n461) );
  XNOR2_X1 U578 ( .A(n462), .B(n461), .ZN(n473) );
  INV_X1 U579 ( .A(n724), .ZN(n468) );
  NAND2_X1 U580 ( .A1(n728), .A2(G234), .ZN(n471) );
  XNOR2_X1 U581 ( .A(n471), .B(n470), .ZN(n521) );
  NAND2_X1 U582 ( .A1(G221), .A2(n521), .ZN(n472) );
  XNOR2_X2 U583 ( .A(G128), .B(KEYINPUT64), .ZN(n474) );
  XNOR2_X2 U584 ( .A(n474), .B(G143), .ZN(n489) );
  INV_X1 U585 ( .A(G107), .ZN(n476) );
  NAND2_X1 U586 ( .A1(G104), .A2(n476), .ZN(n479) );
  NAND2_X1 U587 ( .A1(n477), .A2(G107), .ZN(n478) );
  NAND2_X1 U588 ( .A1(G227), .A2(n728), .ZN(n480) );
  XNOR2_X1 U589 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n723), .B(n483), .ZN(n700) );
  NOR2_X1 U591 ( .A1(n700), .A2(G902), .ZN(n485) );
  INV_X1 U592 ( .A(n661), .ZN(n599) );
  NAND2_X1 U593 ( .A1(G224), .A2(n728), .ZN(n488) );
  NAND2_X1 U594 ( .A1(n698), .A2(n494), .ZN(n495) );
  NAND2_X1 U595 ( .A1(G214), .A2(n496), .ZN(n675) );
  XNOR2_X1 U596 ( .A(n497), .B(KEYINPUT14), .ZN(n498) );
  NAND2_X1 U597 ( .A1(G952), .A2(n498), .ZN(n690) );
  NOR2_X1 U598 ( .A1(G953), .A2(n690), .ZN(n565) );
  NAND2_X1 U599 ( .A1(G902), .A2(n498), .ZN(n499) );
  XOR2_X1 U600 ( .A(KEYINPUT88), .B(n499), .Z(n500) );
  NAND2_X1 U601 ( .A1(G953), .A2(n500), .ZN(n561) );
  NOR2_X1 U602 ( .A1(G898), .A2(n561), .ZN(n501) );
  NOR2_X1 U603 ( .A1(n565), .A2(n501), .ZN(n502) );
  NOR2_X2 U604 ( .A1(n582), .A2(n502), .ZN(n503) );
  NAND2_X1 U605 ( .A1(G221), .A2(n504), .ZN(n505) );
  XNOR2_X1 U606 ( .A(KEYINPUT21), .B(n505), .ZN(n658) );
  XNOR2_X1 U607 ( .A(G143), .B(n506), .ZN(n507) );
  XNOR2_X1 U608 ( .A(n507), .B(n347), .ZN(n511) );
  XNOR2_X1 U609 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U610 ( .A(n511), .B(n510), .ZN(n515) );
  XOR2_X1 U611 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n513) );
  NAND2_X1 U612 ( .A1(G214), .A2(n532), .ZN(n512) );
  XNOR2_X1 U613 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U614 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U615 ( .A(n724), .B(n516), .ZN(n623) );
  NOR2_X1 U616 ( .A1(G902), .A2(n623), .ZN(n518) );
  XNOR2_X1 U617 ( .A(KEYINPUT13), .B(G475), .ZN(n517) );
  XNOR2_X1 U618 ( .A(n518), .B(n517), .ZN(n537) );
  INV_X1 U619 ( .A(n537), .ZN(n544) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(G122), .Z(n520) );
  XNOR2_X1 U621 ( .A(n520), .B(n519), .ZN(n525) );
  XOR2_X1 U622 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n523) );
  NAND2_X1 U623 ( .A1(G217), .A2(n521), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U625 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U626 ( .A(n527), .B(n526), .ZN(n707) );
  NOR2_X1 U627 ( .A1(G902), .A2(n707), .ZN(n528) );
  XNOR2_X1 U628 ( .A(G478), .B(n528), .ZN(n543) );
  NAND2_X1 U629 ( .A1(n544), .A2(n543), .ZN(n678) );
  NAND2_X1 U630 ( .A1(n539), .A2(n356), .ZN(n529) );
  XNOR2_X1 U631 ( .A(G101), .B(G146), .ZN(n530) );
  NAND2_X1 U632 ( .A1(n532), .A2(G210), .ZN(n533) );
  NOR2_X1 U633 ( .A1(G902), .A2(n629), .ZN(n535) );
  INV_X1 U634 ( .A(n568), .ZN(n548) );
  NAND2_X1 U635 ( .A1(n556), .A2(n548), .ZN(n536) );
  NOR2_X1 U636 ( .A1(n537), .A2(n543), .ZN(n649) );
  INV_X1 U637 ( .A(n657), .ZN(n551) );
  INV_X1 U638 ( .A(n658), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n551), .A2(n566), .ZN(n662) );
  NOR2_X1 U640 ( .A1(n662), .A2(n586), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT95), .B(n538), .ZN(n671) );
  XNOR2_X1 U642 ( .A(n542), .B(KEYINPUT100), .ZN(n559) );
  OR2_X1 U643 ( .A1(n544), .A2(n543), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT78), .B(n580), .Z(n547) );
  XOR2_X1 U645 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n546) );
  XNOR2_X1 U646 ( .A(KEYINPUT80), .B(n548), .ZN(n549) );
  NAND2_X1 U647 ( .A1(n549), .A2(n599), .ZN(n550) );
  NOR2_X1 U648 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U649 ( .A(n552), .B(KEYINPUT79), .ZN(n553) );
  NOR2_X1 U650 ( .A1(n378), .A2(n553), .ZN(n555) );
  XNOR2_X1 U651 ( .A(KEYINPUT32), .B(n555), .ZN(n739) );
  NOR2_X1 U652 ( .A1(n737), .A2(n739), .ZN(n557) );
  NAND2_X1 U653 ( .A1(n560), .A2(KEYINPUT44), .ZN(n558) );
  XOR2_X1 U654 ( .A(KEYINPUT103), .B(n561), .Z(n562) );
  NOR2_X1 U655 ( .A1(G900), .A2(n562), .ZN(n563) );
  XNOR2_X1 U656 ( .A(n563), .B(KEYINPUT104), .ZN(n564) );
  NOR2_X1 U657 ( .A1(n565), .A2(n564), .ZN(n575) );
  NAND2_X1 U658 ( .A1(n657), .A2(n566), .ZN(n567) );
  NAND2_X1 U659 ( .A1(n593), .A2(n675), .ZN(n569) );
  NOR2_X1 U660 ( .A1(n599), .A2(n569), .ZN(n570) );
  XOR2_X1 U661 ( .A(KEYINPUT43), .B(n570), .Z(n571) );
  XNOR2_X1 U662 ( .A(n571), .B(KEYINPUT105), .ZN(n572) );
  NAND2_X1 U663 ( .A1(n584), .A2(n675), .ZN(n573) );
  NOR2_X1 U664 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U665 ( .A1(n578), .A2(n611), .ZN(n579) );
  XOR2_X1 U666 ( .A(KEYINPUT107), .B(n581), .Z(n736) );
  INV_X1 U667 ( .A(KEYINPUT74), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n592), .A2(KEYINPUT47), .ZN(n591) );
  AND2_X1 U669 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U670 ( .A(n586), .ZN(n587) );
  NAND2_X1 U671 ( .A1(n358), .A2(n587), .ZN(n607) );
  INV_X1 U672 ( .A(n680), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n645), .A2(n589), .ZN(n590) );
  XNOR2_X1 U674 ( .A(n591), .B(n590), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n592), .A2(KEYINPUT47), .ZN(n600) );
  XNOR2_X1 U676 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n597) );
  NOR2_X1 U677 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U678 ( .A(n597), .B(n596), .Z(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n653) );
  AND2_X1 U680 ( .A1(n600), .A2(n653), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n676), .A2(n675), .ZN(n679) );
  NOR2_X1 U683 ( .A1(n678), .A2(n679), .ZN(n606) );
  XNOR2_X1 U684 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n605) );
  XNOR2_X1 U685 ( .A(n606), .B(n605), .ZN(n674) );
  NOR2_X1 U686 ( .A1(n674), .A2(n607), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n609), .B(n608), .ZN(n740) );
  INV_X1 U689 ( .A(KEYINPUT40), .ZN(n615) );
  INV_X1 U690 ( .A(n676), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n740), .A2(n742), .ZN(n616) );
  INV_X1 U692 ( .A(KEYINPUT46), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n649), .A2(n618), .ZN(n654) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT82), .ZN(n620) );
  INV_X1 U695 ( .A(KEYINPUT76), .ZN(n621) );
  INV_X1 U696 ( .A(KEYINPUT59), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U699 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n628) );
  INV_X1 U700 ( .A(KEYINPUT63), .ZN(n632) );
  XNOR2_X1 U701 ( .A(n633), .B(n632), .ZN(G57) );
  XNOR2_X1 U702 ( .A(G101), .B(n634), .ZN(n635) );
  XNOR2_X1 U703 ( .A(n635), .B(KEYINPUT111), .ZN(G3) );
  NAND2_X1 U704 ( .A1(n379), .A2(n353), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n636), .B(KEYINPUT112), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n347), .B(n637), .ZN(G6) );
  XOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n640) );
  NAND2_X1 U708 ( .A1(n649), .A2(n379), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n642) );
  XOR2_X1 U710 ( .A(G107), .B(KEYINPUT113), .Z(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(n641), .ZN(G9) );
  XOR2_X1 U712 ( .A(G128), .B(KEYINPUT29), .Z(n644) );
  NAND2_X1 U713 ( .A1(n645), .A2(n649), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(G30) );
  NAND2_X1 U715 ( .A1(n645), .A2(n353), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n646), .B(G146), .ZN(G48) );
  NAND2_X1 U717 ( .A1(n650), .A2(n353), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U719 ( .A(G113), .B(n648), .ZN(G15) );
  NAND2_X1 U720 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n651), .B(G116), .ZN(G18) );
  XOR2_X1 U722 ( .A(G125), .B(KEYINPUT37), .Z(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(G27) );
  XNOR2_X1 U724 ( .A(G134), .B(n654), .ZN(G36) );
  XOR2_X1 U725 ( .A(G140), .B(n655), .Z(G42) );
  NOR2_X1 U726 ( .A1(n674), .A2(n683), .ZN(n656) );
  XOR2_X1 U727 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n660) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n669) );
  XOR2_X1 U730 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n664) );
  NAND2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT116), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT51), .B(n672), .Z(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n686) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U744 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n687), .B(KEYINPUT52), .ZN(n688) );
  XNOR2_X1 U746 ( .A(KEYINPUT118), .B(n688), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n693) );
  XOR2_X1 U748 ( .A(KEYINPUT53), .B(n694), .Z(G75) );
  XOR2_X1 U749 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n696) );
  XNOR2_X1 U750 ( .A(KEYINPUT81), .B(KEYINPUT55), .ZN(n695) );
  XNOR2_X1 U751 ( .A(n696), .B(n695), .ZN(n697) );
  XOR2_X1 U752 ( .A(n380), .B(n697), .Z(n699) );
  XOR2_X1 U753 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n702) );
  XNOR2_X1 U754 ( .A(n700), .B(KEYINPUT120), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U756 ( .A1(n709), .A2(G469), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n713), .A2(n705), .ZN(G54) );
  NAND2_X1 U759 ( .A1(G478), .A2(n709), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n713), .A2(n708), .ZN(G63) );
  NAND2_X1 U762 ( .A1(G217), .A2(n709), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U764 ( .A1(n713), .A2(n712), .ZN(G66) );
  NAND2_X1 U765 ( .A1(G953), .A2(G224), .ZN(n714) );
  XNOR2_X1 U766 ( .A(KEYINPUT61), .B(n714), .ZN(n715) );
  NAND2_X1 U767 ( .A1(n715), .A2(G898), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n716), .B(KEYINPUT121), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n722) );
  OR2_X1 U770 ( .A1(G898), .A2(n728), .ZN(n719) );
  XNOR2_X1 U771 ( .A(n720), .B(KEYINPUT122), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(G69) );
  XOR2_X1 U773 ( .A(n723), .B(n724), .Z(n725) );
  XOR2_X1 U774 ( .A(KEYINPUT123), .B(n725), .Z(n730) );
  XOR2_X1 U775 ( .A(KEYINPUT124), .B(n730), .Z(n726) );
  XOR2_X1 U776 ( .A(n727), .B(n726), .Z(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n734) );
  XNOR2_X1 U778 ( .A(G227), .B(n730), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U780 ( .A1(G953), .A2(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U782 ( .A(KEYINPUT125), .B(n735), .Z(G72) );
  XOR2_X1 U783 ( .A(G143), .B(n736), .Z(G45) );
  XOR2_X1 U784 ( .A(n737), .B(G122), .Z(G24) );
  XOR2_X1 U785 ( .A(G119), .B(KEYINPUT126), .Z(n738) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(G21) );
  XOR2_X1 U787 ( .A(G137), .B(n740), .Z(n741) );
  XNOR2_X1 U788 ( .A(KEYINPUT127), .B(n741), .ZN(G39) );
  XNOR2_X1 U789 ( .A(G131), .B(n742), .ZN(G33) );
endmodule

