//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1337, new_n1338,
    new_n1339, new_n1341, new_n1342, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT64), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G1), .B2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n206), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT68), .B(G200), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  INV_X1    g0048(.A(G45), .ZN(new_n249));
  AOI21_X1  g0049(.A(G1), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n252), .A3(G274), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n254), .B1(G226), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G222), .A2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G223), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n212), .A2(G1), .A3(G13), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(G33), .B2(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n266), .C1(G77), .C2(new_n259), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n247), .B1(new_n258), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT69), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n269), .A2(KEYINPUT10), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n258), .A2(new_n267), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G190), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G150), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n206), .A2(G33), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n275), .B1(new_n201), .B2(new_n206), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n264), .A2(new_n265), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G50), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n278), .A2(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n264), .A2(new_n265), .A3(new_n282), .A4(new_n279), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n205), .A2(G20), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(G50), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT9), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n284), .A2(KEYINPUT9), .A3(new_n288), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n271), .A2(new_n273), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n269), .A2(KEYINPUT10), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n294), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n272), .A2(G169), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n272), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n289), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n295), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n276), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(new_n274), .B1(G20), .B2(G77), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT15), .B(G87), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(new_n277), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n306), .A2(new_n280), .B1(new_n202), .B2(new_n283), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n286), .A2(G77), .A3(new_n287), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n254), .B1(G244), .B2(new_n257), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G232), .A2(G1698), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n261), .A2(G238), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n259), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(KEYINPUT67), .A2(G107), .ZN(new_n314));
  NAND2_X1  g0114(.A1(KEYINPUT67), .A2(G107), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n313), .B(new_n266), .C1(new_n259), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n247), .B1(new_n310), .B2(new_n317), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n309), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n309), .B(new_n325), .C1(G179), .C2(new_n318), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n302), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g0130(.A(G226), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n261), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G33), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n231), .A2(G1698), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n330), .A2(new_n332), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G97), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT70), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(new_n339), .A3(new_n266), .ZN(new_n340));
  INV_X1    g0140(.A(G274), .ZN(new_n341));
  INV_X1    g0141(.A(new_n214), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n251), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n257), .A2(G238), .B1(new_n343), .B2(new_n250), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n339), .B1(new_n338), .B2(new_n266), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT13), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n338), .A2(new_n266), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(new_n340), .A4(new_n344), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n347), .A2(G179), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT73), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT73), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n347), .A2(new_n354), .A3(new_n351), .A4(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  INV_X1    g0157(.A(G238), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n253), .B1(new_n358), .B2(new_n256), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n251), .B1(new_n213), .B2(new_n215), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n337), .B2(new_n336), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n359), .B1(new_n361), .B2(new_n339), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n350), .B1(new_n362), .B2(new_n349), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n345), .A2(KEYINPUT13), .A3(new_n346), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n357), .B(G169), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT72), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n347), .A2(new_n351), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n367), .A2(new_n370), .A3(new_n357), .A4(G169), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n356), .A2(new_n366), .A3(new_n369), .A4(new_n371), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n277), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n373));
  INV_X1    g0173(.A(new_n274), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(KEYINPUT71), .B1(new_n281), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n373), .A2(KEYINPUT71), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n280), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT11), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G68), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n205), .B2(G20), .ZN(new_n381));
  OR3_X1    g0181(.A1(new_n282), .A2(KEYINPUT12), .A3(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT12), .B1(new_n282), .B2(G68), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n286), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n377), .B2(new_n378), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n372), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n347), .A2(G190), .A3(new_n351), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n389), .A2(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n367), .A2(G200), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n252), .A2(G232), .A3(new_n255), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n253), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT74), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n333), .A2(KEYINPUT74), .A3(G33), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n330), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n331), .A2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G223), .B2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n396), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  AOI211_X1 g0203(.A(G179), .B(new_n395), .C1(new_n266), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n266), .ZN(new_n405));
  INV_X1    g0205(.A(new_n395), .ZN(new_n406));
  AOI21_X1  g0206(.A(G169), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT76), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n331), .B2(G1698), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n410), .A2(new_n330), .A3(new_n398), .A4(new_n399), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n360), .B1(new_n411), .B2(new_n396), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n324), .B1(new_n412), .B2(new_n395), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT76), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n405), .A2(new_n298), .A3(new_n406), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n276), .B1(new_n205), .B2(G20), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n286), .B1(new_n283), .B2(new_n276), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n280), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n398), .A2(new_n330), .A3(new_n399), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT7), .B1(new_n422), .B2(G20), .ZN(new_n423));
  AND2_X1   g0223(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n424));
  NOR2_X1   g0224(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n400), .A2(new_n206), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(G68), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G58), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n380), .ZN(new_n430));
  NOR2_X1   g0230(.A1(G58), .A2(G68), .ZN(new_n431));
  OAI21_X1  g0231(.A(G20), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G159), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n433), .B2(new_n374), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT16), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n421), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n426), .B1(new_n259), .B2(G20), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n330), .A2(new_n334), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n380), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n435), .B1(new_n441), .B2(new_n434), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n420), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT18), .B1(new_n417), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n427), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT7), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n400), .B2(new_n206), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n445), .A2(new_n447), .A3(new_n380), .ZN(new_n448));
  INV_X1    g0248(.A(new_n436), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n442), .B(new_n280), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G200), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n412), .B2(new_n395), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n405), .A2(new_n319), .A3(new_n406), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(KEYINPUT77), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n395), .B1(new_n403), .B2(new_n266), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT77), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n319), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n450), .A2(new_n454), .A3(new_n419), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n450), .A2(new_n419), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT18), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n408), .A4(new_n416), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n443), .A2(KEYINPUT17), .A3(new_n457), .A4(new_n454), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n444), .A2(new_n460), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n328), .A2(new_n393), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G244), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1698), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n398), .A2(new_n399), .A3(new_n468), .A4(new_n330), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G250), .A2(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(KEYINPUT4), .A2(G244), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(G1698), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n259), .A2(new_n474), .B1(G33), .B2(G283), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n360), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n205), .B(G45), .C1(new_n248), .C2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G41), .ZN(new_n479));
  OAI211_X1 g0279(.A(G257), .B(new_n252), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n252), .A2(G274), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT78), .B1(new_n478), .B2(G41), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT78), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(new_n248), .A3(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n478), .A2(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n249), .A2(G1), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n480), .B1(new_n481), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n476), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n274), .A2(G77), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n491), .A2(new_n492), .A3(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(G97), .B(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n490), .B1(new_n495), .B2(new_n206), .ZN(new_n496));
  INV_X1    g0296(.A(new_n316), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n438), .B2(new_n440), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n280), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n282), .A2(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n329), .A2(G1), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n285), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(G97), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n489), .A2(new_n324), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n471), .A2(new_n475), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n488), .B1(new_n505), .B2(new_n266), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n298), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT80), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n277), .A2(KEYINPUT19), .A3(new_n492), .ZN(new_n510));
  NOR2_X1   g0310(.A1(G87), .A2(G97), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n314), .A2(new_n511), .A3(new_n315), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n337), .A2(new_n206), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n510), .B1(new_n514), .B2(KEYINPUT19), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n398), .A2(new_n399), .A3(new_n206), .A4(new_n330), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n380), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n280), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n305), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n282), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G87), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n285), .A2(new_n522), .A3(new_n501), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n518), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(G250), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n249), .B2(G1), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n205), .A2(new_n341), .A3(G45), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n252), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n467), .A2(G1698), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(G238), .B2(G1698), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n400), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n530), .B1(new_n534), .B2(new_n266), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n247), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n509), .B1(new_n525), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n512), .B2(new_n513), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n539), .A2(new_n510), .B1(new_n380), .B2(new_n516), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n520), .B1(new_n540), .B2(new_n280), .ZN(new_n541));
  INV_X1    g0341(.A(new_n247), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G238), .A2(G1698), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n467), .B2(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n544), .A2(new_n330), .A3(new_n398), .A4(new_n399), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n360), .B1(new_n545), .B2(new_n531), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n546), .B2(new_n530), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n541), .A2(new_n547), .A3(KEYINPUT80), .A4(new_n524), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n534), .A2(new_n266), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n529), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT81), .B1(new_n550), .B2(new_n319), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n535), .A2(new_n552), .A3(G190), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n537), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT79), .B1(new_n489), .B2(new_n319), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n499), .A2(new_n503), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n506), .A2(new_n559), .A3(G190), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n489), .A2(G200), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n502), .A2(new_n519), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n518), .A2(new_n521), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n550), .A2(new_n324), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n535), .A2(new_n298), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AND4_X1   g0367(.A1(new_n508), .A2(new_n555), .A3(new_n562), .A4(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n330), .A2(new_n334), .A3(new_n206), .A4(G87), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT22), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  INV_X1    g0372(.A(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(G20), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n277), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n314), .A2(G20), .A3(new_n315), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT23), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n571), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n516), .A2(new_n570), .A3(new_n522), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT24), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n422), .A2(KEYINPUT22), .A3(new_n206), .A4(G87), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n576), .B1(new_n570), .B2(new_n569), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT24), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n579), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n421), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G13), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(G1), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(G20), .A3(new_n573), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT25), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  AOI22_X1  g0393(.A1(G107), .A2(new_n502), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(G250), .A2(G1698), .ZN(new_n597));
  INV_X1    g0397(.A(G257), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(G1698), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(new_n330), .A3(new_n398), .A4(new_n399), .ZN(new_n600));
  XNOR2_X1  g0400(.A(KEYINPUT84), .B(G294), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G33), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n360), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G264), .B(new_n252), .C1(new_n477), .C2(new_n479), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n481), .B2(new_n487), .ZN(new_n606));
  OAI21_X1  g0406(.A(G169), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n606), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n598), .A2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G250), .B2(G1698), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n400), .A2(new_n610), .B1(new_n329), .B2(new_n601), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n266), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(G179), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n607), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n607), .B2(new_n613), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n596), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n582), .A2(new_n586), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n280), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n451), .B1(new_n604), .B2(new_n606), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n608), .A2(new_n319), .A3(new_n612), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n622), .A3(new_n594), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT86), .B1(new_n617), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n615), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(new_n594), .ZN(new_n627));
  INV_X1    g0427(.A(new_n616), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n623), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n575), .A2(G20), .ZN(new_n635));
  AOI21_X1  g0435(.A(G20), .B1(G33), .B2(G283), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n329), .A2(G97), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n280), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT83), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT20), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n639), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n636), .B2(new_n637), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n280), .A2(new_n645), .A3(new_n635), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT82), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT82), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n280), .A2(new_n645), .A3(new_n648), .A4(new_n635), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(G116), .B1(new_n285), .B2(new_n501), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n282), .A2(new_n575), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n644), .A2(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(G257), .A2(G1698), .ZN(new_n654));
  INV_X1    g0454(.A(G264), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(G1698), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(new_n330), .A3(new_n398), .A4(new_n399), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n439), .A2(G303), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n360), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n252), .B1(new_n477), .B2(new_n479), .ZN(new_n660));
  INV_X1    g0460(.A(G270), .ZN(new_n661));
  OAI22_X1  g0461(.A1(new_n660), .A2(new_n661), .B1(new_n487), .B2(new_n481), .ZN(new_n662));
  OAI21_X1  g0462(.A(G169), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n634), .B1(new_n653), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n639), .A2(new_n641), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT83), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n650), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n651), .A2(new_n652), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(KEYINPUT21), .B(G169), .C1(new_n659), .C2(new_n662), .ZN(new_n671));
  INV_X1    g0471(.A(new_n662), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n655), .A2(G1698), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(G257), .B2(G1698), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n658), .B1(new_n400), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n266), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(G179), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n664), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(G200), .B1(new_n659), .B2(new_n662), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n659), .A2(new_n662), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G190), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n653), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n466), .A2(new_n568), .A3(new_n633), .A4(new_n685), .ZN(G372));
  INV_X1    g0486(.A(new_n300), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n444), .A2(new_n463), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n460), .A2(new_n464), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n326), .B1(new_n390), .B2(new_n391), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n372), .B2(new_n387), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT89), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AOI211_X1 g0494(.A(KEYINPUT89), .B(new_n691), .C1(new_n372), .C2(new_n387), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n689), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n295), .A2(new_n296), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n687), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n489), .A2(new_n324), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n700), .A2(new_n507), .A3(new_n557), .ZN(new_n701));
  XOR2_X1   g0501(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n555), .A2(new_n701), .A3(new_n567), .A4(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT26), .ZN(new_n705));
  NOR4_X1   g0505(.A1(new_n546), .A2(KEYINPUT81), .A3(new_n319), .A4(new_n530), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n552), .B1(new_n535), .B2(G190), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n541), .A2(new_n547), .A3(new_n524), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n567), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n705), .B1(new_n710), .B2(new_n508), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n499), .B(new_n503), .C1(new_n506), .C2(new_n451), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n559), .B1(new_n506), .B2(G190), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n715), .A2(new_n560), .B1(new_n507), .B2(new_n504), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n607), .A2(new_n613), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n587), .B2(new_n595), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n718), .B(new_n679), .C1(KEYINPUT21), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n709), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n565), .A2(new_n566), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n721), .A2(new_n554), .B1(new_n722), .B2(new_n564), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n716), .A2(new_n720), .A3(new_n623), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n567), .B(KEYINPUT87), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n712), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n466), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n699), .A2(new_n727), .ZN(G369));
  NOR3_X1   g0528(.A1(new_n588), .A2(G1), .A3(G20), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT90), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT27), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G213), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G343), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n627), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n625), .A2(new_n631), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n617), .A2(new_n737), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT91), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(KEYINPUT91), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n737), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n653), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n685), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n680), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n746), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n718), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n747), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n680), .A2(new_n737), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n757), .B1(new_n745), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n754), .A2(new_n759), .ZN(G399));
  INV_X1    g0560(.A(new_n209), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G41), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G1), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n512), .A2(G116), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n765), .B1(new_n218), .B2(new_n763), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT29), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n567), .B(KEYINPUT87), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n562), .A2(new_n508), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n520), .B(new_n523), .C1(new_n540), .C2(new_n280), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n771), .B(new_n547), .C1(new_n706), .C2(new_n707), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n623), .A2(new_n772), .A3(new_n567), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n629), .A2(new_n664), .A3(new_n679), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n769), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n555), .A2(new_n701), .A3(new_n567), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(KEYINPUT94), .A3(new_n702), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n723), .A2(KEYINPUT26), .A3(new_n701), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(KEYINPUT94), .B1(new_n777), .B2(new_n702), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n768), .B1(new_n782), .B2(new_n747), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n726), .A2(new_n747), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(KEYINPUT29), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AND4_X1   g0586(.A1(new_n664), .A2(new_n684), .A3(new_n679), .A4(new_n747), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n568), .A2(new_n625), .A3(new_n631), .A4(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n659), .A2(new_n662), .A3(new_n298), .ZN(new_n789));
  INV_X1    g0589(.A(new_n605), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n604), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n789), .A2(new_n506), .A3(new_n535), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT30), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n298), .B1(new_n604), .B2(new_n606), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n682), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT92), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n549), .B2(new_n529), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n506), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n535), .A2(new_n797), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n550), .A2(new_n604), .A3(new_n790), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n802), .A2(KEYINPUT30), .A3(new_n506), .A4(new_n789), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n794), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT31), .B1(new_n804), .B2(new_n737), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT93), .ZN(new_n806));
  AND3_X1   g0606(.A1(new_n804), .A2(KEYINPUT31), .A3(new_n737), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n805), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT93), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n788), .B(new_n806), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G330), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n786), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n767), .B1(new_n813), .B2(G1), .ZN(G364));
  NOR2_X1   g0614(.A1(new_n588), .A2(G20), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n205), .B1(new_n815), .B2(G45), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n762), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(new_n751), .B2(G330), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(G330), .B2(new_n751), .ZN(new_n820));
  INV_X1    g0620(.A(new_n818), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n216), .B1(G20), .B2(new_n324), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n822), .A2(KEYINPUT95), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(KEYINPUT95), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G13), .A2(G33), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G20), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT96), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n761), .A2(new_n439), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(G355), .B1(new_n575), .B2(new_n761), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n761), .A2(new_n422), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(G45), .B2(new_n218), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n245), .A2(new_n249), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n206), .A2(new_n298), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G200), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(G190), .ZN(new_n840));
  INV_X1    g0640(.A(G317), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT33), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n841), .A2(KEYINPUT33), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR4_X1   g0644(.A1(new_n206), .A2(new_n298), .A3(new_n319), .A4(G200), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(G322), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n844), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT100), .ZN(new_n852));
  NOR2_X1   g0652(.A1(G190), .A2(G200), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n838), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n259), .B1(new_n855), .B2(G311), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n319), .A2(G179), .A3(G200), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n206), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n839), .A2(new_n319), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G326), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n856), .B1(new_n601), .B2(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n206), .A2(G179), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n853), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT98), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(KEYINPUT98), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(G329), .ZN(new_n869));
  INV_X1    g0669(.A(G283), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n542), .A2(new_n863), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(G190), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G303), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n319), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n869), .B1(new_n870), .B2(new_n873), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n852), .A2(new_n862), .A3(new_n877), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n878), .A2(KEYINPUT101), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(KEYINPUT101), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n873), .A2(new_n573), .ZN(new_n881));
  INV_X1    g0681(.A(new_n858), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n882), .A2(G97), .B1(new_n855), .B2(G77), .ZN(new_n883));
  INV_X1    g0683(.A(new_n840), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n883), .B1(new_n281), .B2(new_n860), .C1(new_n380), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n849), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n881), .B(new_n885), .C1(G58), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n867), .A2(new_n433), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT32), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n875), .A2(G87), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n259), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT99), .Z(new_n892));
  NAND3_X1  g0692(.A1(new_n887), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n879), .A2(new_n880), .A3(new_n893), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n821), .B(new_n837), .C1(new_n894), .C2(new_n825), .ZN(new_n895));
  INV_X1    g0695(.A(new_n828), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n751), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n820), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(G396));
  INV_X1    g0699(.A(new_n825), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n827), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT102), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n859), .A2(G137), .B1(new_n855), .B2(G159), .ZN(new_n903));
  INV_X1    g0703(.A(G150), .ZN(new_n904));
  INV_X1    g0704(.A(G143), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n903), .B1(new_n904), .B2(new_n884), .C1(new_n849), .C2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT34), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n422), .B1(new_n429), .B2(new_n858), .C1(new_n876), .C2(new_n281), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n872), .A2(G68), .ZN(new_n910));
  INV_X1    g0710(.A(G132), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n867), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n907), .B2(new_n906), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n439), .B1(new_n854), .B2(new_n575), .C1(new_n858), .C2(new_n492), .ZN(new_n915));
  INV_X1    g0715(.A(G294), .ZN(new_n916));
  INV_X1    g0716(.A(G311), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n849), .A2(new_n916), .B1(new_n917), .B2(new_n867), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n872), .A2(G87), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n876), .B2(new_n573), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n870), .A2(new_n884), .B1(new_n860), .B2(new_n874), .ZN(new_n921));
  OR4_X1    g0721(.A1(new_n915), .A2(new_n918), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n818), .B1(G77), .B2(new_n902), .C1(new_n923), .C2(new_n900), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n326), .A2(new_n737), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n309), .A2(new_n737), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n326), .B1(new_n322), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n924), .B1(new_n826), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n327), .A2(new_n747), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n726), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n784), .A2(new_n929), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(KEYINPUT103), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(new_n811), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n818), .B1(new_n936), .B2(new_n811), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n930), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(G384));
  NOR2_X1   g0740(.A1(new_n815), .A2(new_n205), .ZN(new_n941));
  INV_X1    g0741(.A(G330), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n387), .A2(new_n737), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n388), .A2(new_n392), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n392), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n387), .B(new_n737), .C1(new_n372), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n929), .B1(new_n788), .B2(new_n808), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT38), .ZN(new_n951));
  INV_X1    g0751(.A(new_n735), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n408), .B2(new_n416), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n435), .B1(new_n448), .B2(new_n434), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n420), .B1(new_n954), .B2(new_n437), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n458), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT105), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT37), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(new_n956), .B2(KEYINPUT37), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT37), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n960), .B(new_n458), .C1(new_n953), .C2(new_n443), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n958), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n955), .A2(new_n735), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n465), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n951), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n735), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n954), .A2(new_n437), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n419), .ZN(new_n972));
  INV_X1    g0772(.A(new_n457), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n456), .B1(new_n455), .B2(new_n319), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n973), .B1(new_n452), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n970), .A2(new_n972), .B1(new_n443), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT105), .B1(new_n976), .B2(new_n960), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT37), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n978), .A3(new_n961), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(KEYINPUT38), .A3(new_n965), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n967), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT40), .B1(new_n950), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n443), .A2(new_n735), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n465), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n970), .A2(new_n461), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT106), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT37), .A4(new_n458), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n458), .B1(new_n953), .B2(new_n443), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n986), .B1(new_n970), .B2(new_n461), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n960), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(new_n987), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n951), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n980), .A2(new_n992), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT40), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n982), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n788), .A2(new_n808), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n466), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n942), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT107), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT104), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n327), .A2(new_n747), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n769), .B1(new_n774), .B2(new_n720), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n712), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1002), .B1(new_n1005), .B2(new_n925), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n932), .A2(KEYINPUT104), .A3(new_n926), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n981), .A3(new_n947), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT39), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n993), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n967), .A2(KEYINPUT39), .A3(new_n980), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n372), .A2(new_n387), .A3(new_n747), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n688), .A2(new_n735), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1009), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n466), .B1(new_n783), .B2(new_n785), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n699), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1017), .B(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n941), .B1(new_n1001), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n1001), .B2(new_n1020), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n495), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1023), .A2(KEYINPUT35), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(KEYINPUT35), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1024), .A2(G116), .A3(new_n217), .A4(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT36), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n430), .A2(new_n218), .A3(new_n202), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n380), .A2(G50), .ZN(new_n1029));
  OAI211_X1 g0829(.A(G1), .B(new_n588), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1022), .A2(new_n1027), .A3(new_n1030), .ZN(G367));
  AOI22_X1  g0831(.A1(new_n833), .A2(new_n237), .B1(new_n761), .B2(new_n519), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n821), .B1(new_n829), .B2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G68), .A2(new_n882), .B1(new_n859), .B2(G143), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n849), .B2(new_n904), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT111), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n259), .B1(new_n281), .B2(new_n854), .C1(new_n884), .C2(new_n433), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G77), .B2(new_n872), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n868), .A2(G137), .B1(G58), .B2(new_n875), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n872), .A2(G97), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n400), .C1(new_n870), .C2(new_n854), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n849), .A2(new_n874), .B1(new_n841), .B2(new_n867), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n875), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT46), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n876), .B2(new_n575), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n917), .A2(new_n860), .B1(new_n884), .B2(new_n601), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n316), .B2(new_n882), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1042), .A2(new_n1052), .A3(KEYINPUT47), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n825), .ZN(new_n1054));
  AOI21_X1  g0854(.A(KEYINPUT47), .B1(new_n1042), .B2(new_n1052), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1033), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT112), .Z(new_n1057));
  NOR2_X1   g0857(.A1(new_n747), .A2(new_n771), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n710), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n769), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1057), .B1(new_n896), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n716), .B1(new_n558), .B2(new_n747), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n701), .A2(new_n737), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n759), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(KEYINPUT109), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT109), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n759), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT45), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT44), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n759), .B2(new_n1066), .ZN(new_n1074));
  OR3_X1    g0874(.A1(new_n759), .A2(new_n1073), .A3(new_n1066), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1071), .A2(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1068), .A2(new_n1070), .A3(KEYINPUT45), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n754), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1070), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1069), .B1(new_n759), .B2(new_n1066), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1072), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1075), .A2(new_n1074), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1081), .A2(new_n1077), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n753), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n745), .A2(new_n758), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n745), .A2(new_n758), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n752), .B(KEYINPUT110), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n813), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1078), .A2(new_n1084), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n813), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n762), .B(KEYINPUT41), .Z(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n817), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n508), .B1(new_n1064), .B2(new_n629), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n747), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n745), .A2(new_n758), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n1066), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT42), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT42), .B1(new_n1101), .B2(new_n1066), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1062), .A2(KEYINPUT43), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT108), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1102), .B(new_n1103), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT108), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n1107), .A4(new_n1100), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1062), .A2(KEYINPUT43), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1106), .A2(new_n1108), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1109), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n753), .A2(new_n1066), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1063), .B1(new_n1098), .B2(new_n1119), .ZN(G387));
  INV_X1    g0920(.A(new_n1089), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1091), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1121), .A2(new_n1122), .B1(new_n786), .B2(new_n812), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n762), .A3(new_n1092), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n831), .A2(new_n765), .B1(new_n573), .B2(new_n761), .ZN(new_n1125));
  AOI211_X1 g0925(.A(G45), .B(new_n765), .C1(G68), .C2(G77), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT50), .B1(new_n303), .B2(new_n281), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n303), .A2(KEYINPUT50), .A3(new_n281), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n833), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n234), .A2(new_n249), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n821), .B1(new_n830), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n876), .A2(new_n202), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT113), .B(G150), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n868), .B2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n1043), .C1(new_n281), .C2(new_n849), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n859), .A2(G159), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT114), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n422), .B1(new_n380), .B2(new_n854), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n884), .A2(new_n276), .B1(new_n305), .B2(new_n858), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n840), .A2(G311), .B1(new_n855), .B2(G303), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n850), .B2(new_n860), .C1(new_n849), .C2(new_n841), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT48), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n875), .A2(new_n602), .B1(G283), .B2(new_n882), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1150), .A2(KEYINPUT49), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n400), .B1(new_n861), .B2(new_n867), .C1(new_n873), .C2(new_n575), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1150), .B2(KEYINPUT49), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1142), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1133), .B1(new_n1154), .B2(new_n900), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n746), .B2(new_n828), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n817), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1124), .A2(new_n1158), .ZN(G393));
  AOI21_X1  g0959(.A(new_n754), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1083), .A2(new_n753), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1092), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n762), .A3(new_n1094), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1078), .A2(new_n1084), .A3(new_n817), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n829), .B1(new_n492), .B2(new_n209), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n242), .A2(new_n761), .A3(new_n422), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n818), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n849), .A2(new_n917), .B1(new_n841), .B2(new_n860), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n867), .A2(new_n850), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n881), .C1(G283), .C2(new_n875), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n439), .B1(new_n854), .B2(new_n916), .C1(new_n858), .C2(new_n575), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G303), .B2(new_n840), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n849), .A2(new_n433), .B1(new_n904), .B2(new_n860), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT51), .Z(new_n1177));
  OAI221_X1 g0977(.A(new_n919), .B1(new_n905), .B2(new_n867), .C1(new_n876), .C2(new_n380), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n400), .B1(new_n855), .B2(new_n303), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n202), .B2(new_n858), .C1(new_n884), .C2(new_n281), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1175), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1167), .B1(new_n1182), .B2(new_n825), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1066), .B2(new_n896), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1164), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1163), .A2(new_n1185), .ZN(G390));
  NAND3_X1  g0986(.A1(new_n947), .A2(new_n948), .A3(G330), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT104), .B1(new_n932), .B2(new_n926), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1002), .B(new_n925), .C1(new_n726), .C2(new_n931), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n947), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1191), .A2(new_n1013), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n993), .A2(new_n1013), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n782), .A2(new_n747), .A3(new_n928), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n926), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n947), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1188), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n777), .A2(new_n702), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT94), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n779), .A3(new_n778), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n737), .B1(new_n1201), .B2(new_n776), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n925), .B1(new_n1202), .B2(new_n928), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n947), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n993), .B(new_n1013), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n929), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n810), .A2(new_n947), .A3(G330), .A4(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1014), .B1(new_n1008), .B2(new_n947), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT39), .B1(new_n980), .B2(new_n992), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n979), .A2(KEYINPUT38), .A3(new_n965), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT38), .B1(new_n979), .B2(new_n965), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1209), .B1(new_n1212), .B2(KEYINPUT39), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1205), .B(new_n1207), .C1(new_n1208), .C2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1197), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n810), .A2(G330), .A3(new_n1206), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1204), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1187), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1008), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n948), .A2(G330), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1203), .B(new_n1207), .C1(new_n947), .C2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n466), .A2(G330), .A3(new_n996), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n699), .A2(new_n1018), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1224), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1197), .A3(new_n1214), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n762), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1197), .A2(new_n1214), .A3(new_n817), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n860), .A2(new_n870), .B1(new_n854), .B2(new_n492), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n316), .B2(new_n840), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT117), .Z(new_n1234));
  OAI22_X1  g1034(.A1(new_n849), .A2(new_n575), .B1(new_n202), .B2(new_n858), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT118), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n868), .A2(G294), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n439), .A2(new_n1237), .A3(new_n890), .A4(new_n910), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1234), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(KEYINPUT54), .B(G143), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n259), .B1(new_n854), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G128), .ZN(new_n1242));
  INV_X1    g1042(.A(G137), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1242), .A2(new_n860), .B1(new_n884), .B2(new_n1243), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1241), .B(new_n1244), .C1(G159), .C2(new_n882), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n886), .A2(G132), .B1(G125), .B2(new_n868), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n875), .A2(new_n1135), .ZN(new_n1247));
  XOR2_X1   g1047(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1248));
  XNOR2_X1  g1048(.A(new_n1247), .B(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n872), .A2(G50), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1245), .A2(new_n1246), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n900), .B1(new_n1239), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n902), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n821), .B(new_n1252), .C1(new_n276), .C2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1213), .B2(new_n827), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1230), .A2(new_n1231), .A3(new_n1255), .ZN(G378));
  NAND2_X1  g1056(.A1(new_n1229), .A2(new_n1225), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1009), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n980), .A2(new_n992), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT40), .ZN(new_n1260));
  OAI21_X1  g1060(.A(G330), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n952), .A2(new_n289), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n301), .B(new_n1262), .Z(new_n1263));
  XNOR2_X1  g1063(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1263), .B(new_n1265), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n982), .A2(new_n1261), .A3(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1263), .B(new_n1264), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT40), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1212), .B2(new_n949), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n942), .B1(new_n994), .B2(new_n993), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1268), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1258), .B1(new_n1267), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT122), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1266), .B1(new_n982), .B2(new_n1261), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1270), .A2(new_n1271), .A3(new_n1268), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1017), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1275), .A2(new_n1017), .A3(new_n1276), .A4(KEYINPUT122), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1257), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT57), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n763), .B1(new_n1283), .B2(new_n1257), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1278), .A2(new_n817), .A3(new_n1279), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n873), .A2(new_n429), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n886), .B2(G107), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n870), .B2(new_n867), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n882), .A2(G68), .B1(new_n855), .B2(new_n519), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n1290), .B1(new_n492), .B2(new_n884), .C1(new_n575), .C2(new_n860), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n422), .A2(G41), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NOR4_X1   g1093(.A1(new_n1289), .A2(new_n1134), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1294), .B(KEYINPUT119), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT58), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(G33), .A2(G41), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1292), .A2(G50), .A3(new_n1298), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n858), .A2(new_n904), .B1(new_n854), .B2(new_n1243), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n884), .A2(new_n911), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1300), .B(new_n1301), .C1(G125), .C2(new_n859), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1302), .B1(new_n1242), .B2(new_n849), .C1(new_n876), .C2(new_n1240), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1303), .A2(KEYINPUT59), .ZN(new_n1304));
  INV_X1    g1104(.A(G124), .ZN(new_n1305));
  OAI221_X1 g1105(.A(new_n1298), .B1(new_n1305), .B2(new_n867), .C1(new_n873), .C2(new_n433), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1303), .B2(KEYINPUT59), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1299), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n825), .B1(new_n1297), .B2(new_n1309), .ZN(new_n1310));
  XOR2_X1   g1110(.A(new_n1310), .B(KEYINPUT120), .Z(new_n1311));
  OAI21_X1  g1111(.A(new_n818), .B1(new_n901), .B2(G50), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(KEYINPUT121), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1311), .B(new_n1313), .C1(new_n1266), .C2(new_n827), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1286), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1285), .A2(new_n1315), .ZN(G375));
  NAND2_X1  g1116(.A1(new_n1222), .A2(new_n817), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n400), .B(new_n1287), .C1(G150), .C2(new_n855), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n886), .A2(G137), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n868), .A2(G128), .B1(G159), .B2(new_n875), .ZN(new_n1320));
  OAI22_X1  g1120(.A1(new_n884), .A2(new_n1240), .B1(new_n281), .B2(new_n858), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(G132), .B2(new_n859), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  OAI221_X1 g1123(.A(new_n439), .B1(new_n858), .B2(new_n305), .C1(new_n497), .C2(new_n854), .ZN(new_n1324));
  OAI22_X1  g1124(.A1(new_n202), .A2(new_n873), .B1(new_n876), .B2(new_n492), .ZN(new_n1325));
  OAI22_X1  g1125(.A1(new_n849), .A2(new_n870), .B1(new_n874), .B2(new_n867), .ZN(new_n1326));
  OAI22_X1  g1126(.A1(new_n575), .A2(new_n884), .B1(new_n860), .B2(new_n916), .ZN(new_n1327));
  OR4_X1    g1127(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n900), .B1(new_n1323), .B2(new_n1328), .ZN(new_n1329));
  AOI211_X1 g1129(.A(new_n821), .B(new_n1329), .C1(new_n380), .C2(new_n1253), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1330), .B1(new_n947), .B2(new_n827), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1317), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1219), .A2(new_n1224), .A3(new_n1221), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1226), .A2(new_n1097), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(G381));
  NAND3_X1  g1136(.A1(new_n1124), .A2(new_n1158), .A3(new_n898), .ZN(new_n1337));
  OR2_X1    g1137(.A1(new_n1337), .A2(G384), .ZN(new_n1338));
  OR3_X1    g1138(.A1(new_n1338), .A2(G378), .A3(G381), .ZN(new_n1339));
  OR4_X1    g1139(.A1(G387), .A2(new_n1339), .A3(G390), .A4(G375), .ZN(G407));
  INV_X1    g1140(.A(G378), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n736), .ZN(new_n1342));
  OAI211_X1 g1142(.A(G407), .B(G213), .C1(G375), .C2(new_n1342), .ZN(G409));
  NAND2_X1  g1143(.A1(G393), .A2(G396), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1337), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1163), .A2(new_n1345), .A3(new_n1185), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1163), .B2(new_n1185), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(G387), .A2(new_n1346), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1345), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(G390), .A2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1163), .A2(new_n1345), .A3(new_n1185), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1096), .B1(new_n1094), .B2(new_n813), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1118), .B(new_n1117), .C1(new_n1352), .C2(new_n817), .ZN(new_n1353));
  AOI22_X1  g1153(.A1(new_n1350), .A2(new_n1351), .B1(new_n1353), .B2(new_n1063), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1348), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1285), .A2(G378), .A3(new_n1315), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1277), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1017), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1358));
  OAI21_X1  g1158(.A(KEYINPUT123), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT123), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1273), .A2(new_n1360), .A3(new_n1277), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1359), .A2(new_n817), .A3(new_n1361), .ZN(new_n1362));
  OAI211_X1 g1162(.A(new_n1362), .B(new_n1314), .C1(new_n1280), .C2(new_n1096), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(new_n1341), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1356), .A2(new_n1364), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n733), .A2(G343), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1365), .A2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT125), .ZN(new_n1369));
  XNOR2_X1  g1169(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1334), .B1(new_n1228), .B2(new_n1371), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1219), .A2(new_n1224), .A3(KEYINPUT60), .A4(new_n1221), .ZN(new_n1373));
  AND2_X1   g1173(.A1(new_n1373), .A2(new_n762), .ZN(new_n1374));
  AOI211_X1 g1174(.A(new_n939), .B(new_n1332), .C1(new_n1372), .C2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1372), .ZN(new_n1376));
  AOI21_X1  g1176(.A(G384), .B1(new_n1376), .B2(new_n1333), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1369), .B1(new_n1375), .B2(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1373), .A2(new_n762), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1226), .A2(new_n1370), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1379), .B1(new_n1380), .B2(new_n1334), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n939), .B1(new_n1381), .B2(new_n1332), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1376), .A2(G384), .A3(new_n1333), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1382), .A2(KEYINPUT125), .A3(new_n1383), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1366), .A2(G2897), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1378), .A2(new_n1384), .A3(new_n1385), .ZN(new_n1386));
  OAI211_X1 g1186(.A(G2897), .B(new_n1366), .C1(new_n1375), .C2(new_n1377), .ZN(new_n1387));
  AND2_X1   g1187(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(KEYINPUT61), .B1(new_n1368), .B2(new_n1388), .ZN(new_n1389));
  AOI21_X1  g1189(.A(new_n1366), .B1(new_n1356), .B2(new_n1364), .ZN(new_n1390));
  AND2_X1   g1190(.A1(new_n1378), .A2(new_n1384), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1390), .A2(new_n1391), .ZN(new_n1392));
  XOR2_X1   g1192(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1393));
  NAND2_X1  g1193(.A1(new_n1392), .A2(new_n1393), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1390), .A2(KEYINPUT63), .A3(new_n1391), .ZN(new_n1395));
  NAND4_X1  g1195(.A1(new_n1355), .A2(new_n1389), .A3(new_n1394), .A4(new_n1395), .ZN(new_n1396));
  INV_X1    g1196(.A(KEYINPUT62), .ZN(new_n1397));
  AND3_X1   g1197(.A1(new_n1390), .A2(new_n1397), .A3(new_n1391), .ZN(new_n1398));
  INV_X1    g1198(.A(KEYINPUT61), .ZN(new_n1399));
  NAND2_X1  g1199(.A1(new_n1386), .A2(new_n1387), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1399), .B1(new_n1390), .B2(new_n1400), .ZN(new_n1401));
  AOI21_X1  g1201(.A(new_n1397), .B1(new_n1390), .B2(new_n1391), .ZN(new_n1402));
  NOR3_X1   g1202(.A1(new_n1398), .A2(new_n1401), .A3(new_n1402), .ZN(new_n1403));
  OAI21_X1  g1203(.A(new_n1396), .B1(new_n1403), .B2(new_n1355), .ZN(G405));
  INV_X1    g1204(.A(KEYINPUT127), .ZN(new_n1405));
  INV_X1    g1205(.A(new_n1356), .ZN(new_n1406));
  AOI21_X1  g1206(.A(G378), .B1(new_n1285), .B2(new_n1315), .ZN(new_n1407));
  OAI211_X1 g1207(.A(new_n1405), .B(new_n1391), .C1(new_n1406), .C2(new_n1407), .ZN(new_n1408));
  NOR2_X1   g1208(.A1(new_n1375), .A2(new_n1377), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(G375), .A2(new_n1341), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1410), .A2(new_n1356), .ZN(new_n1411));
  OAI21_X1  g1211(.A(new_n1408), .B1(new_n1409), .B2(new_n1411), .ZN(new_n1412));
  AOI21_X1  g1212(.A(new_n1405), .B1(new_n1411), .B2(new_n1391), .ZN(new_n1413));
  OAI22_X1  g1213(.A1(new_n1412), .A2(new_n1413), .B1(new_n1348), .B2(new_n1354), .ZN(new_n1414));
  NAND2_X1  g1214(.A1(new_n1411), .A2(new_n1391), .ZN(new_n1415));
  NAND2_X1  g1215(.A1(new_n1415), .A2(KEYINPUT127), .ZN(new_n1416));
  OR2_X1    g1216(.A1(new_n1411), .A2(new_n1409), .ZN(new_n1417));
  NAND4_X1  g1217(.A1(new_n1355), .A2(new_n1416), .A3(new_n1417), .A4(new_n1408), .ZN(new_n1418));
  NAND2_X1  g1218(.A1(new_n1414), .A2(new_n1418), .ZN(G402));
endmodule


