//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  AND2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT22), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n207), .B2(KEYINPUT29), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n211), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n212), .A2(KEYINPUT81), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n212), .A2(KEYINPUT81), .ZN(new_n219));
  OAI21_X1  g018(.A(G155gat), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n220), .B2(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n215), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n211), .A2(new_n216), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(KEYINPUT2), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT85), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n208), .A2(new_n230), .A3(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n207), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT81), .B(G162gat), .Z(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(G155gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n202), .B(new_n224), .C1(new_n237), .C2(new_n217), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G228gat), .ZN(new_n240));
  INV_X1    g039(.A(G233gat), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(KEYINPUT86), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n228), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n244), .A2(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT86), .B1(new_n232), .B2(new_n242), .ZN(new_n247));
  OAI21_X1  g046(.A(G22gat), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  INV_X1    g048(.A(G22gat), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n243), .A4(new_n245), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT31), .B(G50gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n248), .A2(new_n251), .A3(KEYINPUT87), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G113gat), .A2(G120gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G113gat), .A2(G120gat), .ZN(new_n263));
  OR3_X1    g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT1), .ZN(new_n264));
  NOR2_X1   g063(.A1(G127gat), .A2(G134gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT72), .B(G127gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G134gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271));
  NAND2_X1  g070(.A1(G127gat), .A2(G134gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(G127gat), .A2(G134gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT74), .B1(new_n274), .B2(new_n265), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT1), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n263), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT73), .A3(new_n261), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n262), .B2(new_n263), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n276), .A2(KEYINPUT75), .A3(new_n281), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n270), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n288));
  INV_X1    g087(.A(G169gat), .ZN(new_n289));
  INV_X1    g088(.A(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(KEYINPUT23), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT67), .B(KEYINPUT24), .ZN(new_n297));
  AND2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT68), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT24), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(new_n298), .B2(KEYINPUT24), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n299), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n296), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n299), .A2(new_n307), .A3(KEYINPUT69), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n289), .A2(KEYINPUT23), .ZN(new_n314));
  AND2_X1   g113(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n294), .B1(KEYINPUT23), .B2(new_n287), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT66), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT66), .ZN(new_n320));
  INV_X1    g119(.A(new_n316), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n292), .B(new_n320), .C1(new_n323), .C2(new_n314), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n298), .A2(KEYINPUT24), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n300), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n325), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n319), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n312), .A2(new_n313), .B1(new_n293), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n291), .A2(KEYINPUT71), .A3(KEYINPUT26), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n333), .B(new_n287), .C1(new_n291), .C2(KEYINPUT26), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT71), .B1(new_n291), .B2(KEYINPUT26), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT27), .B(G183gat), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n336), .A2(new_n341), .A3(new_n306), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n286), .B1(new_n332), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n298), .B1(new_n301), .B2(new_n303), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n309), .B1(new_n344), .B2(new_n305), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n297), .A2(KEYINPUT68), .A3(new_n298), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n311), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n296), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n313), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n293), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n276), .A2(KEYINPUT75), .A3(new_n281), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT75), .B1(new_n276), .B2(new_n281), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n269), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n341), .A3(new_n306), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n343), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G227gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n241), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n361), .A2(KEYINPUT34), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(KEYINPUT34), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n359), .A3(new_n356), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n343), .A2(new_n356), .A3(KEYINPUT76), .A4(new_n359), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT33), .B1(new_n369), .B2(new_n370), .ZN(new_n372));
  XOR2_X1   g171(.A(G15gat), .B(G43gat), .Z(new_n373));
  XNOR2_X1  g172(.A(G71gat), .B(G99gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n371), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  AOI221_X4 g176(.A(new_n366), .B1(KEYINPUT33), .B2(new_n375), .C1(new_n369), .C2(new_n370), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n365), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n372), .A2(new_n376), .ZN(new_n380));
  INV_X1    g179(.A(new_n371), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n378), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n364), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n252), .A2(new_n253), .A3(new_n257), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n260), .A2(new_n379), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT0), .ZN(new_n388));
  XNOR2_X1  g187(.A(G57gat), .B(G85gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n354), .A2(new_n227), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n226), .B(new_n269), .C1(new_n352), .C2(new_n353), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n392), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n394), .A2(new_n400), .A3(KEYINPUT4), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n394), .B2(KEYINPUT4), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(new_n221), .B2(new_n225), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n238), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n286), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n405), .A2(new_n238), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT82), .B1(new_n409), .B2(new_n354), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n396), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT84), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT83), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n400), .A3(KEYINPUT4), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n407), .B1(new_n286), .B2(new_n406), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(new_n354), .A3(KEYINPUT82), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n397), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n399), .B1(new_n412), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n419), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n426), .A2(KEYINPUT5), .A3(new_n397), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n391), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n421), .B1(new_n417), .B2(new_n420), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n398), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n427), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n390), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT6), .B(new_n391), .C1(new_n423), .C2(new_n427), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT78), .B1(new_n332), .B2(new_n342), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n351), .A2(new_n439), .A3(new_n355), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G226gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n241), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT29), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n351), .A2(new_n443), .A3(new_n355), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n207), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n443), .A3(new_n440), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n351), .A2(new_n355), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n444), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n207), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT79), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n448), .A2(new_n453), .A3(new_n207), .A4(new_n450), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n447), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456));
  XOR2_X1   g255(.A(G8gat), .B(G36gat), .Z(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT80), .ZN(new_n458));
  XOR2_X1   g257(.A(G64gat), .B(G92gat), .Z(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n452), .A2(new_n454), .ZN(new_n463));
  INV_X1    g262(.A(new_n447), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT30), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n455), .A2(new_n461), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n437), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT35), .B1(new_n386), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n384), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT77), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n379), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n382), .A2(new_n383), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT77), .A3(new_n365), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n260), .A2(new_n385), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n437), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n470), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n463), .A2(new_n486), .A3(new_n464), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n461), .A2(KEYINPUT38), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n448), .A2(new_n233), .A3(new_n450), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n489), .A2(KEYINPUT37), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n445), .A2(new_n446), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n207), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n487), .A2(new_n493), .B1(new_n455), .B2(new_n461), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n435), .A2(new_n494), .A3(new_n436), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n487), .A2(new_n460), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n455), .A2(new_n486), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT38), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n500), .B(KEYINPUT38), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n396), .B1(new_n424), .B2(new_n425), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n395), .A2(new_n397), .ZN(new_n505));
  OR3_X1    g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n504), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n390), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n506), .A2(KEYINPUT40), .A3(new_n390), .A4(new_n507), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n510), .A2(new_n428), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n480), .A2(new_n482), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n502), .A2(new_n513), .A3(new_n477), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n379), .A2(new_n384), .A3(KEYINPUT36), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n476), .B2(KEYINPUT36), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n260), .A2(new_n385), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n469), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n485), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n485), .B(KEYINPUT90), .C1(new_n515), .C2(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT12), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  INV_X1    g331(.A(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n535), .A2(new_n536), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n537), .A2(new_n538), .B1(KEYINPUT15), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n537), .B1(KEYINPUT15), .B2(new_n539), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT17), .ZN(new_n543));
  XOR2_X1   g342(.A(G15gat), .B(G22gat), .Z(new_n544));
  INV_X1    g343(.A(G1gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(G8gat), .B1(new_n546), .B2(KEYINPUT94), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n545), .A2(KEYINPUT93), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(KEYINPUT93), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n546), .B1(new_n551), .B2(new_n544), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n547), .B(new_n552), .ZN(new_n553));
  MUX2_X1   g352(.A(new_n542), .B(new_n543), .S(new_n553), .Z(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(KEYINPUT18), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n553), .B(new_n542), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n555), .B(KEYINPUT13), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n531), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n559), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT18), .B1(new_n554), .B2(new_n555), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n562), .B(new_n565), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n525), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT100), .ZN(new_n571));
  NOR2_X1   g370(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G99gat), .B(G106gat), .Z(new_n574));
  INV_X1    g373(.A(G99gat), .ZN(new_n575));
  INV_X1    g374(.A(G106gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT8), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT101), .B(G85gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(G92gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT102), .ZN(new_n580));
  OR3_X1    g379(.A1(new_n573), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n574), .B1(new_n573), .B2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n583), .A2(new_n542), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT41), .ZN(new_n585));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n583), .ZN(new_n587));
  OAI221_X1 g386(.A(new_n584), .B1(new_n585), .B2(new_n586), .C1(new_n543), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n585), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n590), .A2(new_n592), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT103), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OR3_X1    g396(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n593), .B2(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G57gat), .B(G64gat), .Z(new_n601));
  AND2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(KEYINPUT9), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT9), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(KEYINPUT96), .ZN(new_n605));
  NOR2_X1   g404(.A1(G71gat), .A2(G78gat), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n605), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n603), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT97), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n608), .B(KEYINPUT98), .Z(new_n618));
  OAI21_X1  g417(.A(new_n553), .B1(new_n618), .B2(new_n609), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n617), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G230gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n241), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n583), .A2(new_n618), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT105), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n608), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n608), .A2(new_n631), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n583), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n583), .A2(new_n633), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n627), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n627), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n645), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n600), .A2(new_n625), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT106), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n651), .A2(KEYINPUT106), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n568), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n437), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n545), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n654), .A2(new_n483), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(KEYINPUT42), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n657), .B(KEYINPUT107), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(G8gat), .ZN(new_n662));
  OAI221_X1 g461(.A(new_n659), .B1(KEYINPUT42), .B2(new_n658), .C1(new_n660), .C2(new_n662), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n654), .B2(new_n517), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT77), .B1(new_n474), .B2(new_n365), .ZN(new_n665));
  AOI211_X1 g464(.A(new_n472), .B(new_n364), .C1(new_n382), .C2(new_n383), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n384), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(G15gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n664), .B1(new_n654), .B2(new_n668), .ZN(G1326gat));
  OR3_X1    g468(.A1(new_n654), .A2(KEYINPUT108), .A3(new_n477), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT108), .B1(new_n654), .B2(new_n477), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT43), .B(G22gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  INV_X1    g473(.A(new_n625), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n650), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n600), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n568), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(G29gat), .A3(new_n437), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT45), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(new_n600), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n514), .A2(KEYINPUT109), .A3(new_n517), .A4(new_n519), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n485), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n686), .A2(new_n516), .B1(new_n469), .B2(new_n518), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT109), .B1(new_n687), .B2(new_n514), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n682), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n600), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n523), .A2(new_n524), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR4_X1   g493(.A1(new_n694), .A2(new_n437), .A3(new_n567), .A4(new_n676), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n680), .B(new_n681), .C1(new_n533), .C2(new_n695), .ZN(G1328gat));
  NAND2_X1  g495(.A1(new_n484), .A2(new_n534), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n678), .A2(KEYINPUT46), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT110), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT46), .B1(new_n678), .B2(new_n697), .ZN(new_n700));
  NOR4_X1   g499(.A1(new_n694), .A2(new_n483), .A3(new_n567), .A4(new_n676), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n699), .B(new_n700), .C1(new_n534), .C2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(new_n694), .ZN(new_n703));
  INV_X1    g502(.A(new_n517), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n676), .A2(new_n567), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n703), .A2(G43gat), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n678), .A2(new_n667), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(G43gat), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g508(.A1(new_n691), .A2(new_n518), .A3(new_n693), .A4(new_n705), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G50gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n477), .A2(G50gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n568), .A2(new_n677), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(KEYINPUT48), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(KEYINPUT111), .A3(G50gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n713), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT111), .B1(new_n710), .B2(G50gat), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT112), .B(new_n715), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n711), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n716), .A3(new_n713), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT112), .B1(new_n723), .B2(new_n715), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n714), .B1(new_n720), .B2(new_n724), .ZN(G1331gat));
  OR2_X1    g524(.A1(new_n684), .A2(new_n688), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n682), .A2(new_n675), .A3(new_n566), .A4(new_n650), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n437), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n484), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  AND2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n733), .B2(new_n732), .ZN(G1333gat));
  NAND2_X1  g535(.A1(new_n728), .A2(new_n704), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n667), .A2(G71gat), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n737), .A2(G71gat), .B1(new_n728), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g539(.A1(new_n728), .A2(new_n518), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT114), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT113), .B(G78gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1335gat));
  NOR2_X1   g543(.A1(new_n625), .A2(new_n566), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n694), .A2(new_n650), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(new_n729), .ZN(new_n748));
  INV_X1    g547(.A(new_n578), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n682), .B(new_n745), .C1(new_n684), .C2(new_n688), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n649), .A2(new_n729), .A3(new_n749), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n748), .A2(new_n749), .B1(new_n754), .B2(new_n755), .ZN(G1336gat));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n752), .A2(KEYINPUT115), .A3(new_n753), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n650), .A2(G92gat), .A3(new_n483), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n750), .A2(new_n760), .A3(new_n751), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n650), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n691), .A2(new_n484), .A3(new_n693), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G92gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n757), .B1(new_n766), .B2(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  AOI211_X1 g567(.A(KEYINPUT116), .B(new_n768), .C1(new_n762), .C2(new_n765), .ZN(new_n769));
  INV_X1    g568(.A(new_n765), .ZN(new_n770));
  INV_X1    g569(.A(new_n759), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n754), .B2(new_n771), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n767), .A2(new_n769), .B1(new_n770), .B2(new_n772), .ZN(G1337gat));
  AND2_X1   g572(.A1(new_n747), .A2(new_n704), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n649), .A2(new_n575), .A3(new_n476), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n774), .A2(new_n575), .B1(new_n754), .B2(new_n775), .ZN(G1338gat));
  AOI21_X1  g575(.A(new_n576), .B1(new_n747), .B2(new_n518), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n649), .A2(new_n576), .A3(new_n518), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT117), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n758), .A2(new_n761), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT53), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n754), .B2(new_n778), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n777), .B2(new_n783), .ZN(G1339gat));
  NAND3_X1  g583(.A1(new_n630), .A2(new_n636), .A3(new_n627), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n638), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n646), .B1(new_n637), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n788), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n791), .A2(new_n566), .A3(new_n647), .A4(new_n792), .ZN(new_n793));
  OAI22_X1  g592(.A1(new_n554), .A2(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n565), .A2(new_n531), .B1(new_n530), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n649), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n793), .A2(new_n796), .A3(KEYINPUT118), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n682), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n598), .A2(new_n599), .A3(new_n795), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n791), .A2(new_n647), .A3(new_n792), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n675), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n651), .A2(new_n566), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n667), .A2(new_n518), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n484), .A2(new_n437), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(G113gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n812), .A2(new_n813), .A3(new_n567), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n809), .A2(new_n811), .ZN(new_n815));
  INV_X1    g614(.A(new_n386), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n566), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n814), .B1(new_n819), .B2(new_n813), .ZN(G1340gat));
  INV_X1    g619(.A(G120gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n812), .A2(new_n821), .A3(new_n650), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n649), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n821), .ZN(G1341gat));
  OAI21_X1  g623(.A(new_n267), .B1(new_n812), .B2(new_n675), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n675), .A2(new_n267), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT119), .ZN(G1342gat));
  OAI21_X1  g627(.A(G134gat), .B1(new_n812), .B2(new_n600), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n809), .A2(new_n682), .A3(new_n811), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n386), .A2(G134gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n830), .A2(KEYINPUT120), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT120), .B1(new_n830), .B2(new_n832), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n833), .A2(KEYINPUT56), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n829), .B1(new_n835), .B2(new_n836), .ZN(G1343gat));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  INV_X1    g637(.A(new_n800), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT118), .B1(new_n793), .B2(new_n796), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n600), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n625), .B1(new_n841), .B2(new_n804), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n838), .B(new_n518), .C1(new_n842), .C2(new_n807), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n811), .A2(new_n517), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n797), .A2(new_n600), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n625), .B1(new_n845), .B2(new_n804), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n518), .B1(new_n846), .B2(new_n807), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(KEYINPUT57), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G141gat), .B1(new_n849), .B2(new_n567), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n704), .A2(new_n477), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n815), .A2(new_n209), .A3(new_n566), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n855), .A3(KEYINPUT58), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n850), .B(new_n852), .C1(new_n854), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n210), .A2(KEYINPUT59), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n815), .A2(new_n851), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n862), .B2(new_n649), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n849), .A2(new_n650), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n653), .A2(new_n567), .A3(new_n652), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n838), .B(new_n518), .C1(new_n865), .C2(new_n846), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n477), .B1(new_n806), .B2(new_n808), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n649), .B(new_n866), .C1(new_n867), .C2(new_n838), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n844), .B(KEYINPUT122), .Z(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT59), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n864), .A2(KEYINPUT59), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n863), .B1(G148gat), .B2(new_n871), .ZN(G1345gat));
  OAI21_X1  g671(.A(G155gat), .B1(new_n849), .B2(new_n675), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n625), .A2(new_n214), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n861), .B2(new_n874), .ZN(G1346gat));
  INV_X1    g674(.A(new_n236), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n851), .A2(new_n876), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n830), .A2(KEYINPUT123), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n236), .B1(new_n849), .B2(new_n600), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT123), .B1(new_n830), .B2(new_n877), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n483), .A2(new_n729), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT124), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n809), .A2(new_n810), .A3(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(new_n289), .A3(new_n567), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n809), .A2(new_n882), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n816), .A3(new_n566), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n289), .B2(new_n888), .ZN(G1348gat));
  AOI211_X1 g688(.A(new_n650), .B(new_n885), .C1(new_n321), .C2(new_n322), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n816), .A3(new_n649), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n290), .B2(new_n891), .ZN(G1349gat));
  OAI21_X1  g691(.A(G183gat), .B1(new_n885), .B2(new_n675), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n887), .A2(new_n816), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n625), .A2(new_n337), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g696(.A1(new_n885), .A2(new_n600), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(G190gat), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n898), .B2(G190gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n682), .A2(new_n338), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n901), .A2(new_n902), .B1(new_n894), .B2(new_n903), .ZN(G1351gat));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n851), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n567), .A2(G197gat), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n905), .A2(KEYINPUT125), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n883), .A2(new_n704), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n866), .B(new_n909), .C1(new_n867), .C2(new_n838), .ZN(new_n910));
  OAI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n567), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT125), .B1(new_n905), .B2(new_n907), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(G1352gat));
  INV_X1    g712(.A(new_n909), .ZN(new_n914));
  OAI21_X1  g713(.A(G204gat), .B1(new_n868), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n650), .A2(G204gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n905), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(KEYINPUT62), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n905), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n915), .B1(new_n918), .B2(new_n920), .ZN(G1353gat));
  NOR2_X1   g720(.A1(new_n675), .A2(G211gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n887), .A2(new_n851), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT126), .ZN(new_n924));
  OAI21_X1  g723(.A(G211gat), .B1(new_n910), .B2(new_n675), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT63), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(G211gat), .C1(new_n910), .C2(new_n675), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(G1354gat));
  OAI21_X1  g728(.A(G218gat), .B1(new_n910), .B2(new_n600), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n600), .A2(G218gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n887), .A2(new_n851), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(KEYINPUT127), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1355gat));
endmodule


