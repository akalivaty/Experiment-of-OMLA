//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n449), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT67), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n475), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n463), .A2(new_n469), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G62), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n504), .A2(G651), .B1(new_n510), .B2(G88), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  AND2_X1   g087(.A1(G50), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT68), .B(new_n513), .C1(new_n517), .C2(new_n505), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n511), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n522), .B1(new_n512), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n506), .A2(KEYINPUT70), .A3(new_n507), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NOR3_X1   g103(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT69), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n530), .B1(new_n508), .B2(new_n509), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n510), .A2(G89), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n528), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n532), .A2(G64), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n510), .A2(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n526), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(new_n532), .A2(G56), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n539), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n551), .B1(new_n550), .B2(new_n549), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT72), .B(G81), .Z(new_n553));
  AOI22_X1  g128(.A1(new_n527), .A2(G43), .B1(new_n510), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  OAI21_X1  g136(.A(new_n523), .B1(new_n517), .B2(new_n505), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n525), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(KEYINPUT73), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n563), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n502), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n510), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  NAND4_X1  g147(.A1(new_n525), .A2(new_n562), .A3(G49), .A4(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT74), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n524), .A2(new_n575), .A3(G49), .A4(new_n525), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n578), .B1(new_n529), .B2(new_n531), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(G87), .B2(new_n510), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G288));
  INV_X1    g156(.A(G73), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT75), .B1(new_n582), .B2(new_n522), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n584), .A2(G73), .A3(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n583), .B(new_n585), .C1(new_n502), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(G48), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n502), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(new_n512), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n539), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n527), .A2(G47), .B1(G85), .B2(new_n510), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(new_n508), .A2(new_n509), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n598), .A2(new_n512), .A3(G92), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n527), .A2(G54), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n598), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n539), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT76), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(G868), .B2(new_n611), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(G868), .B2(new_n611), .ZN(G280));
  INV_X1    g188(.A(new_n604), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n555), .A2(new_n605), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n604), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n605), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g195(.A1(new_n463), .A2(new_n469), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n473), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n475), .A2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n481), .A2(G123), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n460), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(G156));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2084), .B(G2090), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT77), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT79), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n653), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n651), .B(new_n660), .C1(new_n655), .C2(new_n657), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT80), .B(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n668), .A2(new_n671), .A3(new_n675), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT32), .ZN(new_n686));
  INV_X1    g261(.A(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(G16), .A2(G22), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G166), .B2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G23), .B(G288), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(KEYINPUT33), .B(G1976), .Z(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n688), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n696), .A2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G24), .ZN(new_n702));
  INV_X1    g277(.A(G290), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n475), .A2(G131), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT81), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n481), .A2(G119), .ZN(new_n709));
  NOR2_X1   g284(.A1(G95), .A2(G2105), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT82), .ZN(new_n711));
  OAI21_X1  g286(.A(G2104), .B1(new_n460), .B2(G107), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n708), .B(new_n709), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G25), .B(new_n713), .S(G29), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n706), .A2(KEYINPUT84), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n699), .A2(new_n700), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT30), .B(G28), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  OR2_X1    g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  NAND2_X1  g299(.A1(KEYINPUT31), .A2(G11), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n632), .B2(new_n723), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n701), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n701), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n727), .B1(new_n729), .B2(G1966), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G1966), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n701), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n701), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n731), .B1(G1961), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT91), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n556), .B2(G16), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G1341), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G1341), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n701), .A2(G20), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT23), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G299), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n739), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n723), .A2(G32), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n481), .A2(G129), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT90), .Z(new_n747));
  AND2_X1   g322(.A1(new_n473), .A2(G105), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT26), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n748), .B(new_n750), .C1(G141), .C2(new_n475), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n745), .B1(new_n753), .B2(new_n723), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(G164), .A2(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G27), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G2078), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n723), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n723), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT29), .B(G2090), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n756), .A2(new_n760), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n723), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n475), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n481), .A2(G128), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n460), .A2(G116), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n769), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NOR2_X1   g350(.A1(G4), .A2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT85), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n604), .B2(new_n701), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT86), .B(G1348), .Z(new_n779));
  OAI221_X1 g354(.A(new_n775), .B1(new_n778), .B2(new_n779), .C1(new_n754), .C2(new_n755), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n766), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(G160), .A2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(G29), .B1(new_n783), .B2(KEYINPUT24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(KEYINPUT24), .B2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(G2084), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n733), .A2(G1961), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n788), .B(new_n789), .C1(new_n779), .C2(new_n778), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(KEYINPUT89), .A3(G2084), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n723), .A2(G33), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n621), .A2(G127), .ZN(new_n793));
  NAND2_X1  g368(.A1(G115), .A2(G2104), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n460), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n796));
  NAND3_X1  g371(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G139), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n476), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n792), .B1(new_n801), .B2(new_n723), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT88), .B(G2072), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(KEYINPUT89), .B1(new_n787), .B2(G2084), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n781), .A2(new_n790), .A3(new_n791), .A4(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n735), .A2(new_n744), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n720), .A2(new_n721), .A3(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  NAND2_X1  g385(.A1(new_n532), .A2(G67), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n539), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n510), .A2(G93), .ZN(new_n814));
  INV_X1    g389(.A(G55), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n526), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT92), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n555), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n556), .A2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n614), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  INV_X1    g403(.A(new_n817), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n831), .ZN(G145));
  NOR2_X1   g407(.A1(new_n801), .A2(KEYINPUT93), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n475), .A2(G142), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n481), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n460), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n833), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(G164), .B(new_n773), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n752), .A2(new_n840), .B1(new_n801), .B2(KEYINPUT93), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n752), .B2(new_n840), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n839), .B(new_n842), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n713), .B(new_n623), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n844), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(G160), .B(new_n632), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  AOI21_X1  g425(.A(G37), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n848), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT95), .B(KEYINPUT40), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(G395));
  NAND2_X1  g429(.A1(new_n829), .A2(new_n605), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n856));
  XNOR2_X1  g431(.A(G290), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G288), .ZN(new_n858));
  XNOR2_X1  g433(.A(G303), .B(G305), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT98), .B(KEYINPUT42), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n822), .B(new_n618), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n604), .B1(new_n611), .B2(KEYINPUT96), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n865));
  NAND2_X1  g440(.A1(G299), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n864), .B(new_n866), .Z(new_n867));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n864), .B(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT41), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n863), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n870), .B2(new_n863), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n862), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n855), .B1(new_n875), .B2(new_n605), .ZN(G295));
  OAI21_X1  g451(.A(new_n855), .B1(new_n875), .B2(new_n605), .ZN(G331));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  XNOR2_X1  g453(.A(G171), .B(G286), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n820), .B2(new_n821), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n820), .A2(new_n821), .A3(new_n879), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n867), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n872), .ZN(new_n884));
  INV_X1    g459(.A(new_n882), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(new_n880), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n860), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n881), .A2(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n870), .A2(KEYINPUT99), .A3(KEYINPUT41), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n890), .B(new_n891), .C1(new_n872), .C2(KEYINPUT99), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n860), .B1(new_n892), .B2(new_n883), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n889), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n882), .A2(new_n881), .B1(new_n869), .B2(new_n871), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n885), .A2(new_n870), .A3(new_n880), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n898), .B2(new_n860), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n887), .A2(new_n888), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT43), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT44), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT43), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n894), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(G397));
  NAND2_X1  g482(.A1(new_n495), .A2(new_n497), .ZN(new_n908));
  INV_X1    g483(.A(new_n492), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G1384), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT105), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(G164), .B2(G1384), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT100), .B(G40), .Z(new_n918));
  NOR4_X1   g493(.A1(new_n472), .A2(new_n478), .A3(G2084), .A4(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT112), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1966), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT45), .B1(new_n912), .B2(new_n914), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n910), .A2(KEYINPUT45), .A3(new_n911), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n472), .A2(new_n478), .A3(new_n918), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n916), .A2(KEYINPUT112), .A3(new_n917), .A4(new_n919), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n922), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(G8), .ZN(new_n931));
  NAND2_X1  g506(.A1(G286), .A2(G8), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT120), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(G8), .B(new_n935), .C1(new_n930), .C2(G286), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n932), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n930), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT121), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT121), .ZN(new_n943));
  INV_X1    g518(.A(new_n941), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n943), .B(new_n944), .C1(new_n937), .C2(new_n938), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT62), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n938), .ZN(new_n947));
  AOI211_X1 g522(.A(new_n940), .B(new_n935), .C1(new_n930), .C2(G8), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n943), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT62), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n939), .A2(KEYINPUT121), .A3(new_n941), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n912), .A2(new_n926), .A3(new_n914), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n577), .A2(new_n580), .A3(G1976), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(G8), .A3(new_n956), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n957), .A2(KEYINPUT52), .ZN(new_n958));
  INV_X1    g533(.A(G1976), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(G288), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(new_n955), .A3(G8), .A4(new_n956), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT49), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n588), .A2(new_n592), .A3(new_n687), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n687), .B1(new_n588), .B2(new_n592), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G305), .A2(G1981), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n588), .A2(new_n592), .A3(new_n687), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(KEYINPUT49), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n955), .A2(new_n965), .A3(new_n968), .A4(G8), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n954), .B1(new_n958), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n957), .A2(KEYINPUT52), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(KEYINPUT111), .A3(new_n961), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G2090), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n916), .A2(new_n975), .A3(new_n926), .A4(new_n917), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(G164), .B2(G1384), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n925), .A2(new_n926), .A3(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n976), .A2(KEYINPUT107), .B1(new_n691), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n916), .A2(new_n917), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(new_n975), .A4(new_n926), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n511), .B2(new_n519), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n987), .B2(KEYINPUT55), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n598), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n598), .A2(new_n512), .ZN(new_n990));
  INV_X1    g565(.A(G88), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n989), .A2(new_n539), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT68), .B1(new_n512), .B2(new_n513), .ZN(new_n993));
  INV_X1    g568(.A(new_n518), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT109), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n988), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT55), .B(G8), .C1(new_n992), .C2(new_n995), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT108), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n987), .A2(new_n1002), .A3(KEYINPUT55), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n999), .A2(new_n1004), .A3(KEYINPUT110), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT110), .B1(new_n999), .B2(new_n1004), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n984), .A2(new_n1007), .A3(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n915), .B1(new_n912), .B2(new_n914), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n910), .A2(new_n1010), .A3(new_n911), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n926), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1009), .A2(new_n1012), .A3(G2090), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n979), .A2(new_n691), .ZN(new_n1014));
  OAI21_X1  g589(.A(G8), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n999), .A2(new_n1004), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AND4_X1   g593(.A1(KEYINPUT126), .A2(new_n974), .A3(new_n1008), .A4(new_n1018), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n971), .A2(new_n973), .B1(new_n1017), .B2(new_n1015), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT126), .B1(new_n1020), .B2(new_n1008), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n916), .A2(new_n926), .A3(new_n917), .ZN(new_n1022));
  INV_X1    g597(.A(G1961), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n979), .B2(G2078), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n924), .A2(G2078), .A3(new_n927), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G171), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1019), .A2(new_n1021), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n946), .A2(new_n953), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n759), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n472), .A2(new_n478), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n925), .A2(new_n1038), .A3(new_n978), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT125), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1041), .B2(G171), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n1032), .B2(G171), .ZN(new_n1043));
  AND4_X1   g618(.A1(G301), .A2(new_n1040), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1032), .B2(G171), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1047), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n950), .A2(new_n952), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n925), .A2(new_n926), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT56), .B(G2072), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(KEYINPUT115), .A3(new_n978), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1956), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n925), .A2(new_n926), .A3(new_n978), .A4(new_n1052), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n566), .B2(new_n570), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1063), .A2(new_n1053), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT61), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n955), .ZN(new_n1071));
  INV_X1    g646(.A(G2067), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1022), .A2(new_n779), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1073), .B2(new_n604), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1067), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT116), .B1(new_n1073), .B2(new_n604), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1067), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1066), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1022), .A2(new_n779), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(KEYINPUT60), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT118), .A3(new_n604), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1073), .A2(KEYINPUT60), .ZN(new_n1086));
  XOR2_X1   g661(.A(new_n604), .B(KEYINPUT118), .Z(new_n1087));
  NAND3_X1  g662(.A1(new_n1073), .A2(KEYINPUT60), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT58), .B(G1341), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1071), .A2(new_n1090), .B1(G1996), .B2(new_n979), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n556), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT59), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1065), .B1(new_n604), .B2(new_n1073), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1089), .A2(new_n1093), .B1(new_n1067), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1050), .B1(new_n1081), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1067), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1069), .A2(new_n1068), .B1(new_n1074), .B2(new_n1067), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT61), .B1(new_n1077), .B2(new_n1067), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1065), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1102), .A3(KEYINPUT119), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1048), .A2(new_n1049), .A3(new_n1096), .A4(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n931), .A2(G286), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1105), .A2(KEYINPUT63), .A3(new_n1008), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT113), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n979), .A2(new_n691), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n1111));
  OAI21_X1  g686(.A(G8), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1017), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n958), .A2(new_n970), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n986), .B1(new_n980), .B2(new_n983), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1107), .B(new_n1114), .C1(new_n1116), .C2(new_n1016), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1106), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT114), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1106), .B(new_n1121), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1020), .A2(new_n1008), .A3(new_n1105), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1120), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n969), .A2(new_n959), .A3(new_n577), .A4(new_n580), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n986), .B(new_n1071), .C1(new_n1127), .C2(new_n967), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1008), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1114), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1035), .A2(new_n1104), .A3(new_n1126), .A4(new_n1130), .ZN(new_n1131));
  NOR4_X1   g706(.A1(new_n978), .A2(new_n472), .A3(new_n478), .A4(new_n918), .ZN(new_n1132));
  INV_X1    g707(.A(G1996), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT101), .Z(new_n1135));
  XNOR2_X1  g710(.A(new_n1132), .B(KEYINPUT102), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n773), .B(new_n1072), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n753), .B2(new_n1133), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1135), .A2(new_n753), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n713), .B(new_n715), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT103), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1136), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n703), .A2(new_n705), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G290), .A2(G1986), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1132), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT104), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1131), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n715), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n713), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1139), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n773), .A2(G2067), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1136), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1154), .A2(KEYINPUT127), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1137), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1136), .B1(new_n752), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT46), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1135), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1135), .A2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1161), .A2(KEYINPUT47), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(KEYINPUT47), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1145), .A2(new_n1132), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT48), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1162), .A2(new_n1163), .B1(new_n1143), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1154), .A2(KEYINPUT127), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1155), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1149), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g744(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1171));
  OAI211_X1 g745(.A(new_n852), .B(new_n1171), .C1(new_n904), .C2(new_n905), .ZN(G225));
  INV_X1    g746(.A(G225), .ZN(G308));
endmodule


