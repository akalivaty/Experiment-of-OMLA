//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919;
  XOR2_X1   g000(.A(KEYINPUT74), .B(KEYINPUT32), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G134), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI22_X1  g007(.A1(new_n193), .A2(G137), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n195), .A2(new_n196), .A3(new_n191), .A4(G134), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n189), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(new_n192), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G131), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n189), .A3(G131), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(KEYINPUT0), .B2(G128), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT0), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT64), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n211), .A2(new_n212), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT0), .A3(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n205), .A2(new_n206), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n205), .A2(new_n225), .A3(new_n206), .A4(new_n222), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n198), .A2(new_n199), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n191), .A2(G134), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n193), .A2(G137), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT68), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n210), .B1(new_n233), .B2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(G128), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT69), .B1(new_n211), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n219), .A2(new_n237), .A3(new_n233), .A4(G128), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n208), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n227), .A2(new_n243), .A3(new_n230), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n232), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n224), .A2(new_n226), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT30), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G116), .B(G119), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n251), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n227), .A2(new_n230), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n242), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n223), .A2(new_n256), .A3(KEYINPUT30), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n248), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n254), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n223), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT70), .B(G237), .Z(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n258), .A2(new_n260), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT31), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n258), .A2(new_n275), .A3(new_n260), .A4(new_n272), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n260), .B(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n246), .A2(new_n254), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n274), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G472), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  AND4_X1   g097(.A1(KEYINPUT73), .A2(new_n281), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n279), .B1(new_n273), .B2(KEYINPUT31), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n285), .B2(new_n276), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT73), .B1(new_n286), .B2(new_n282), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n188), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT75), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT32), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n258), .A2(new_n260), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(new_n272), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n277), .A2(new_n272), .A3(new_n278), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(KEYINPUT29), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n223), .A2(new_n256), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n254), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n277), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n272), .A2(KEYINPUT29), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n283), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G472), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n292), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n290), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n286), .A2(KEYINPUT73), .A3(new_n282), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n188), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n289), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  XNOR2_X1  g127(.A(G125), .B(G140), .ZN(new_n314));
  MUX2_X1   g128(.A(new_n313), .B(new_n314), .S(KEYINPUT16), .Z(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(G146), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n216), .A2(G119), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n321));
  INV_X1    g135(.A(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G128), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n318), .B2(new_n317), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n321), .B(new_n323), .C1(new_n325), .C2(new_n320), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(G110), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n318), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n316), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n315), .A2(new_n207), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n314), .A2(new_n207), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n329), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n326), .B2(G110), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n332), .B(new_n333), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n335), .A2(new_n336), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT79), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT22), .B(G137), .Z(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n331), .B(new_n343), .C1(new_n337), .C2(new_n338), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n283), .A3(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n347), .B(KEYINPUT25), .Z(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n283), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(new_n350), .B2(new_n347), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G214), .B1(G237), .B2(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G952), .ZN(new_n356));
  AOI211_X1 g170(.A(G953), .B(new_n356), .C1(G234), .C2(G237), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n283), .B(new_n266), .C1(G234), .C2(G237), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT21), .B(G898), .Z(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n221), .A2(G125), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT89), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n221), .A2(new_n364), .A3(G125), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n363), .B(new_n365), .C1(G125), .C2(new_n242), .ZN(new_n366));
  INV_X1    g180(.A(G224), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G953), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n366), .B(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n370), .A2(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n370), .A2(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT80), .A4(G104), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n372), .A2(new_n373), .A3(new_n374), .A4(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(KEYINPUT82), .A3(G104), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n376), .B2(G104), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n371), .A2(G107), .ZN(new_n382));
  OAI211_X1 g196(.A(G101), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT84), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n322), .A3(G116), .ZN(new_n387));
  OAI211_X1 g201(.A(G113), .B(new_n387), .C1(new_n250), .C2(new_n386), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n252), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G101), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT4), .A3(new_n378), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT81), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n391), .A2(new_n394), .A3(KEYINPUT4), .A4(new_n378), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n391), .A2(KEYINPUT4), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n393), .A2(new_n254), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(G110), .B(G122), .Z(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n389), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n389), .B2(new_n397), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n404), .A2(KEYINPUT88), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT88), .B1(new_n404), .B2(new_n405), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n369), .B(new_n403), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n399), .B(KEYINPUT8), .Z(new_n409));
  INV_X1    g223(.A(new_n389), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n388), .A2(new_n252), .B1(new_n378), .B2(new_n383), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n368), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n366), .B1(KEYINPUT7), .B2(new_n413), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n412), .B(new_n402), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n283), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G210), .B1(G237), .B2(G902), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n408), .A2(new_n416), .A3(new_n283), .A4(new_n418), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n355), .B(new_n361), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G128), .B(G143), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n193), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n209), .A2(G128), .ZN(new_n426));
  OAI21_X1  g240(.A(G134), .B1(new_n426), .B2(KEYINPUT13), .ZN(new_n427));
  XNOR2_X1  g241(.A(G116), .B(G122), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n430), .A2(G107), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(G107), .ZN(new_n432));
  OAI221_X1 g246(.A(new_n424), .B1(new_n425), .B2(new_n427), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n423), .B(new_n193), .ZN(new_n434));
  INV_X1    g248(.A(G116), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT14), .A3(G122), .ZN(new_n436));
  INV_X1    g250(.A(new_n428), .ZN(new_n437));
  OAI211_X1 g251(.A(G107), .B(new_n436), .C1(new_n437), .C2(KEYINPUT14), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n434), .B(new_n438), .C1(new_n430), .C2(G107), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT9), .B(G234), .Z(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(new_n349), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n433), .A2(new_n439), .A3(new_n443), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT15), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G478), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n449), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G475), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n267), .A2(G214), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n209), .ZN(new_n456));
  AND4_X1   g270(.A1(G143), .A2(new_n261), .A3(G214), .A4(new_n266), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT17), .A3(G131), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(new_n199), .A3(new_n458), .ZN(new_n461));
  AOI21_X1  g275(.A(G143), .B1(new_n267), .B2(G214), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n462), .B2(new_n457), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n316), .B(new_n460), .C1(new_n464), .C2(KEYINPUT17), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n314), .B(new_n207), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT18), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(new_n199), .ZN(new_n468));
  OAI221_X1 g282(.A(new_n466), .B1(new_n463), .B2(new_n467), .C1(new_n459), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G113), .B(G122), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n371), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n469), .A3(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n454), .B1(new_n476), .B2(new_n283), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n464), .A2(KEYINPUT90), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n314), .B(KEYINPUT19), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n207), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n480), .A2(KEYINPUT91), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(KEYINPUT91), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(new_n332), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n461), .A2(new_n484), .A3(new_n463), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n486), .A2(new_n469), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n475), .B1(new_n487), .B2(new_n472), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n454), .A4(new_n283), .ZN(new_n490));
  INV_X1    g304(.A(new_n475), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n472), .B1(new_n486), .B2(new_n469), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n454), .B(new_n283), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT20), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n477), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n422), .A2(new_n453), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n384), .B1(new_n239), .B2(new_n241), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n385), .B2(new_n242), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n205), .A2(new_n206), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(KEYINPUT85), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT12), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n499), .A2(KEYINPUT85), .A3(new_n504), .A4(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT83), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n497), .B2(KEYINPUT10), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT10), .ZN(new_n509));
  AOI211_X1 g323(.A(new_n240), .B(new_n234), .C1(new_n236), .C2(new_n238), .ZN(new_n510));
  OAI211_X1 g324(.A(KEYINPUT83), .B(new_n509), .C1(new_n510), .C2(new_n384), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n393), .A2(new_n222), .A3(new_n395), .A4(new_n396), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n385), .A2(KEYINPUT10), .A3(new_n242), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n512), .A2(new_n500), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n266), .A2(G227), .ZN(new_n516));
  XNOR2_X1  g330(.A(G110), .B(G140), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n506), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n501), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n515), .ZN(new_n523));
  INV_X1    g337(.A(new_n518), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT87), .B(G469), .Z(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G469), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n519), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n515), .A2(KEYINPUT86), .A3(new_n518), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n515), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n524), .B1(new_n506), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(G902), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n528), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G221), .B1(new_n442), .B2(G902), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n496), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n311), .A2(new_n353), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n374), .ZN(G3));
  OR2_X1    g356(.A1(new_n286), .A2(new_n282), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n308), .A2(new_n422), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n538), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n352), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n537), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n447), .A2(G478), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n445), .A2(new_n446), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT33), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT33), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n549), .B1(new_n556), .B2(G478), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n495), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n548), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT34), .B(G104), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(G6));
  INV_X1    g376(.A(new_n495), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(new_n453), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n548), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G107), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(G9));
  NOR2_X1   g382(.A1(new_n350), .A2(G902), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n345), .A2(new_n346), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT94), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n343), .A2(KEYINPUT36), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n345), .A2(new_n574), .A3(new_n346), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n573), .B1(new_n571), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n569), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n351), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n308), .A2(new_n543), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n308), .A2(KEYINPUT95), .A3(new_n543), .A4(new_n579), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n540), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT37), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(G110), .Z(G12));
  INV_X1    g400(.A(new_n539), .ZN(new_n587));
  INV_X1    g401(.A(G900), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n357), .B1(new_n358), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n495), .A2(new_n452), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n355), .B1(new_n420), .B2(new_n421), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(KEYINPUT96), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  INV_X1    g409(.A(new_n593), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n595), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n311), .A2(new_n587), .A3(new_n579), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G128), .ZN(G30));
  NAND2_X1  g414(.A1(new_n420), .A2(new_n421), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n601), .B(KEYINPUT97), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT38), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n495), .A2(new_n453), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n603), .A2(new_n354), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n579), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n309), .B1(new_n308), .B2(new_n188), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT75), .B(new_n187), .C1(new_n306), .C2(new_n307), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n272), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n293), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n260), .A3(new_n298), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n283), .ZN(new_n613));
  OAI21_X1  g427(.A(G472), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n609), .A2(new_n292), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n589), .B(KEYINPUT98), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT39), .Z(new_n617));
  NAND2_X1  g431(.A1(new_n587), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n605), .A2(new_n606), .A3(new_n615), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G143), .ZN(G45));
  AOI21_X1  g436(.A(new_n606), .B1(new_n609), .B2(new_n304), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n495), .A2(new_n557), .A3(new_n589), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n593), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(KEYINPUT100), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n623), .A2(new_n587), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G146), .ZN(G48));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n526), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G469), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n526), .A2(new_n631), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n538), .B(new_n528), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n311), .A2(new_n353), .A3(new_n422), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n559), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT41), .B(G113), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G15));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n565), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n435), .ZN(G18));
  OAI21_X1  g456(.A(KEYINPUT102), .B1(new_n635), .B2(new_n596), .ZN(new_n643));
  INV_X1    g457(.A(new_n528), .ZN(new_n644));
  INV_X1    g458(.A(new_n634), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n529), .B1(new_n526), .B2(new_n631), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n538), .A4(new_n593), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n643), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n563), .A2(new_n361), .A3(new_n452), .ZN(new_n651));
  AND4_X1   g465(.A1(new_n311), .A2(new_n650), .A3(new_n579), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n322), .ZN(G21));
  NAND2_X1  g467(.A1(new_n299), .A2(new_n610), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n274), .A2(new_n276), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n282), .A3(new_n283), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n543), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n352), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n636), .A3(new_n422), .A4(new_n604), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G122), .ZN(G24));
  NOR2_X1   g474(.A1(new_n606), .A2(new_n657), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n650), .A2(new_n624), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT103), .B(G125), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G27));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n533), .A2(new_n535), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n283), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n665), .B1(new_n667), .B2(G469), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n533), .A2(new_n535), .A3(new_n665), .A4(new_n283), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n529), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n528), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n601), .A2(new_n355), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n671), .A2(new_n538), .A3(new_n624), .A4(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n311), .A3(new_n353), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n291), .A2(KEYINPUT32), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n353), .B1(new_n303), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n677), .B2(new_n673), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n199), .ZN(G33));
  INV_X1    g494(.A(new_n670), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n536), .B2(new_n529), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n644), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n672), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n546), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n311), .A2(new_n353), .A3(new_n685), .A4(new_n592), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G134), .ZN(G36));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n557), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n690), .B1(new_n691), .B2(new_n495), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n495), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n688), .B2(new_n689), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n692), .B1(new_n694), .B2(new_n690), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n308), .A2(new_n543), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n695), .A2(new_n696), .A3(new_n606), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n672), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n666), .B(KEYINPUT45), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(KEYINPUT46), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n528), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n704), .A2(new_n538), .A3(new_n617), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n697), .A2(KEYINPUT44), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n698), .A2(new_n707), .A3(new_n672), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n700), .A2(new_n705), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G137), .ZN(G39));
  INV_X1    g524(.A(new_n311), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n624), .A2(new_n352), .A3(new_n672), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n704), .A2(KEYINPUT47), .A3(new_n538), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT47), .B1(new_n704), .B2(new_n538), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G140), .ZN(G42));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n603), .B1(new_n717), .B2(KEYINPUT49), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(KEYINPUT49), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n647), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n615), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n547), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n693), .B(new_n722), .C1(new_n647), .C2(new_n719), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n718), .A2(new_n354), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n452), .B(KEYINPUT108), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n725), .A2(new_n495), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n691), .A2(new_n495), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n545), .A2(new_n537), .A3(new_n547), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n584), .A2(new_n729), .A3(new_n659), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n652), .A2(new_n730), .A3(new_n541), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n685), .A2(new_n624), .A3(new_n661), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n678), .A2(new_n686), .A3(new_n675), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n725), .A2(new_n495), .A3(new_n590), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n684), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n726), .A2(KEYINPUT109), .A3(new_n590), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n736), .A2(KEYINPUT110), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT110), .B1(new_n736), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n587), .A3(new_n623), .ZN(new_n741));
  INV_X1    g555(.A(new_n637), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n558), .B2(new_n564), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n731), .A2(new_n733), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n311), .A2(new_n587), .A3(new_n579), .A4(new_n628), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n599), .B(new_n662), .C1(new_n746), .C2(new_n626), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n604), .A2(new_n593), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n748), .A2(new_n683), .A3(new_n546), .A4(new_n589), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n615), .A2(new_n606), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT111), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n744), .B1(new_n745), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(KEYINPUT111), .B(KEYINPUT52), .C1(new_n747), .C2(new_n750), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT53), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n747), .B2(new_n750), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n599), .A2(new_n662), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n615), .A2(new_n606), .A3(new_n749), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n629), .A3(new_n745), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n744), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT54), .B1(new_n754), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n357), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n635), .A2(new_n684), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n353), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n615), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n558), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n695), .A2(new_n763), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(new_n658), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n650), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(G952), .A3(new_n262), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n760), .B1(new_n759), .B2(new_n744), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n776));
  INV_X1    g590(.A(new_n744), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n751), .A2(new_n745), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT53), .A4(new_n753), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT112), .B(new_n760), .C1(new_n759), .C2(new_n744), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n775), .A2(new_n776), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n768), .A2(new_n764), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n677), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(KEYINPUT48), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(KEYINPUT48), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n782), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n762), .A2(new_n772), .A3(new_n781), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n647), .A2(new_n546), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n713), .A2(new_n714), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n791), .B2(KEYINPUT113), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(KEYINPUT113), .B2(new_n791), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n672), .A3(new_n769), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n768), .A2(new_n636), .A3(new_n658), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n354), .A3(new_n603), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT50), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n768), .A2(new_n661), .A3(new_n764), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(KEYINPUT50), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n766), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n563), .A3(new_n691), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT51), .B1(new_n794), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n713), .A2(new_n714), .A3(new_n790), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n769), .A2(new_n672), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n801), .A2(new_n808), .A3(new_n803), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n788), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(G952), .A2(G953), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n724), .B1(new_n810), .B2(new_n811), .ZN(G75));
  NAND3_X1  g626(.A1(new_n775), .A2(new_n779), .A3(new_n780), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(G210), .A3(G902), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n403), .B1(new_n406), .B2(new_n407), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(new_n369), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT55), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n814), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n814), .B2(new_n815), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n266), .A2(G952), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT115), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(G51));
  NAND2_X1  g637(.A1(new_n813), .A2(KEYINPUT54), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n781), .ZN(new_n825));
  NAND2_X1  g639(.A1(G469), .A2(G902), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT57), .Z(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n520), .A2(new_n525), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n813), .A2(G469), .A3(G902), .A4(new_n701), .ZN(new_n832));
  INV_X1    g646(.A(new_n827), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n824), .B2(new_n781), .ZN(new_n834));
  INV_X1    g648(.A(new_n830), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT116), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n821), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(G54));
  NAND4_X1  g653(.A1(new_n813), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n840));
  INV_X1    g654(.A(new_n488), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(new_n821), .ZN(G60));
  NAND2_X1  g658(.A1(new_n554), .A2(new_n555), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n825), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(G478), .A2(G902), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT59), .Z(new_n848));
  NOR2_X1   g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n762), .B2(new_n781), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n845), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n851), .A3(new_n822), .ZN(G63));
  NAND2_X1  g666(.A1(G217), .A2(G902), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT60), .Z(new_n854));
  NAND2_X1  g668(.A1(new_n813), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n822), .B1(new_n855), .B2(new_n570), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n813), .B(new_n854), .C1(new_n576), .C2(new_n577), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT61), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n858), .B(new_n860), .ZN(G66));
  OAI21_X1  g675(.A(G953), .B1(new_n360), .B2(new_n367), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n731), .A2(new_n743), .ZN(new_n863));
  INV_X1    g677(.A(new_n266), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT118), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n816), .B1(G898), .B2(new_n266), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(G69));
  NAND2_X1  g682(.A1(new_n248), .A2(new_n257), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n479), .ZN(new_n870));
  INV_X1    g684(.A(new_n715), .ZN(new_n871));
  INV_X1    g685(.A(new_n747), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n621), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n621), .A2(KEYINPUT62), .A3(new_n872), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n728), .A2(KEYINPUT119), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n618), .A3(new_n684), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n728), .A2(KEYINPUT119), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n311), .A3(new_n353), .A4(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n709), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT120), .B(new_n870), .C1(new_n883), .C2(new_n864), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n864), .B1(new_n877), .B2(new_n882), .ZN(new_n886));
  INV_X1    g700(.A(new_n870), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(KEYINPUT121), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(G227), .A2(G900), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n864), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n700), .A2(new_n706), .A3(new_n708), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n677), .B2(new_n748), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n679), .B1(new_n893), .B2(new_n705), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n715), .A2(new_n686), .A3(new_n872), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n266), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n896), .B(new_n887), .C1(new_n588), .C2(new_n266), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n897), .A2(new_n884), .A3(new_n888), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n891), .B(new_n898), .ZN(G72));
  INV_X1    g713(.A(new_n293), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n863), .A3(new_n895), .ZN(new_n901));
  XNOR2_X1  g715(.A(KEYINPUT122), .B(KEYINPUT63), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT123), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n282), .A2(new_n283), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT124), .Z(new_n906));
  AOI211_X1 g720(.A(new_n900), .B(new_n272), .C1(new_n901), .C2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n906), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n883), .B2(new_n863), .ZN(new_n909));
  INV_X1    g723(.A(new_n611), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n838), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n754), .A2(new_n761), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n273), .A2(KEYINPUT125), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n294), .B(new_n913), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n905), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT126), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT127), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(KEYINPUT127), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n907), .B(new_n911), .C1(new_n918), .C2(new_n919), .ZN(G57));
endmodule


