//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202));
  XNOR2_X1  g001(.A(G99gat), .B(G106gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT7), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT7), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(G85gat), .A3(G92gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT8), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT96), .B(G85gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G92gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n204), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n206), .A2(new_n208), .B1(KEYINPUT8), .B2(new_n210), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n216), .B(new_n203), .C1(G92gat), .C2(new_n213), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  OR2_X1    g018(.A1(G71gat), .A2(G78gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT9), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(G71gat), .A2(G78gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(KEYINPUT9), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT95), .ZN(new_n227));
  NOR3_X1   g026(.A1(new_n226), .A2(new_n227), .A3(new_n221), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n229));
  XOR2_X1   g028(.A(G57gat), .B(G64gat), .Z(new_n230));
  AOI21_X1  g029(.A(KEYINPUT95), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n223), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n218), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT10), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n227), .B1(new_n226), .B2(new_n221), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT95), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n237), .A2(new_n215), .A3(new_n223), .A4(new_n217), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n218), .ZN(new_n240));
  INV_X1    g039(.A(new_n232), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT10), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G230gat), .A2(G233gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT99), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n202), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  AOI211_X1 g046(.A(KEYINPUT101), .B(new_n245), .C1(new_n239), .C2(new_n242), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n233), .B2(new_n238), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G120gat), .B(G148gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(G176gat), .B(G204gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT102), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n243), .A2(new_n246), .ZN(new_n256));
  INV_X1    g055(.A(new_n249), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT100), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n247), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n202), .A3(new_n246), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT102), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n253), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n255), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT103), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n255), .A2(new_n260), .A3(new_n265), .A4(KEYINPUT103), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n241), .A2(KEYINPUT21), .ZN(new_n274));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275));
  INV_X1    g074(.A(G1gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT16), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n275), .A2(G1gat), .ZN(new_n279));
  OAI21_X1  g078(.A(G8gat), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n277), .ZN(new_n281));
  INV_X1    g080(.A(G8gat), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n281), .B(new_n282), .C1(G1gat), .C2(new_n275), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G183gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n237), .A2(KEYINPUT21), .A3(new_n223), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n274), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  INV_X1    g090(.A(new_n274), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G231gat), .A2(G233gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n290), .B2(new_n293), .ZN(new_n298));
  XNOR2_X1  g097(.A(G127gat), .B(G155gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(G211gat), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n300), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n290), .A2(new_n293), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n294), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n304), .B2(new_n296), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n273), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G43gat), .B(G50gat), .Z(new_n307));
  INV_X1    g106(.A(KEYINPUT15), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G43gat), .B(G50gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT14), .ZN(new_n312));
  INV_X1    g111(.A(G29gat), .ZN(new_n313));
  INV_X1    g112(.A(G36gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n315), .A2(new_n316), .B1(G29gat), .B2(G36gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  NAND2_X1  g118(.A1(G29gat), .A2(G36gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(KEYINPUT15), .A3(new_n310), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT17), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n322), .A3(KEYINPUT17), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n218), .ZN(new_n327));
  NAND3_X1  g126(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n240), .A2(new_n323), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G190gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(new_n331), .ZN(new_n334));
  XNOR2_X1  g133(.A(G134gat), .B(G162gat), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n333), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT97), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n339), .A2(KEYINPUT97), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(new_n334), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n337), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT98), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT98), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n345), .A3(new_n337), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n340), .A2(new_n341), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n300), .B1(new_n297), .B2(new_n298), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n304), .A2(new_n302), .A3(new_n296), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n272), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n306), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n271), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT104), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n271), .A2(KEYINPUT104), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G78gat), .B(G106gat), .Z(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G148gat), .ZN(new_n364));
  INV_X1    g163(.A(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G141gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT78), .B1(new_n363), .B2(G148gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  XNOR2_X1  g169(.A(G141gat), .B(G148gat), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n370), .B(KEYINPUT79), .C1(new_n371), .C2(new_n362), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT2), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n369), .A2(new_n372), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n371), .A2(KEYINPUT2), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n381), .A2(new_n375), .A3(new_n377), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G197gat), .B(G204gat), .ZN(new_n386));
  INV_X1    g185(.A(G211gat), .ZN(new_n387));
  INV_X1    g186(.A(G218gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n386), .B1(KEYINPUT22), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G211gat), .B(G218gat), .Z(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n369), .A2(new_n372), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397));
  INV_X1    g196(.A(new_n382), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT82), .B1(new_n380), .B2(new_n382), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT3), .B1(new_n392), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G228gat), .ZN(new_n405));
  INV_X1    g204(.A(G233gat), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n393), .A2(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  OAI221_X1 g207(.A(new_n408), .B1(new_n383), .B2(new_n403), .C1(new_n385), .C2(new_n392), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n360), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(KEYINPUT85), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G22gat), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n407), .A2(KEYINPUT85), .A3(new_n415), .A4(new_n409), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n410), .A2(new_n411), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n414), .A2(new_n416), .B1(new_n418), .B2(new_n359), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G120gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT69), .ZN(new_n422));
  INV_X1    g221(.A(G113gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(G113gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT70), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT1), .ZN(new_n430));
  XNOR2_X1  g229(.A(G127gat), .B(G134gat), .ZN(new_n431));
  AND2_X1   g230(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n433));
  OAI21_X1  g232(.A(G120gat), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT70), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n427), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n429), .A2(new_n430), .A3(new_n431), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n431), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT68), .ZN(new_n439));
  XNOR2_X1  g238(.A(G113gat), .B(G120gat), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n438), .B(new_n439), .C1(KEYINPUT1), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n423), .A2(G120gat), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT1), .B1(new_n427), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT68), .B1(new_n443), .B2(new_n431), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n437), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT71), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n437), .A2(new_n445), .A3(KEYINPUT71), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT25), .ZN(new_n451));
  AND3_X1   g250(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(G183gat), .A2(G190gat), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G169gat), .ZN(new_n456));
  INV_X1    g255(.A(G176gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT23), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(G169gat), .B2(G176gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(G169gat), .A2(G176gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n451), .B1(new_n455), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT64), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT64), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(new_n451), .C1(new_n455), .C2(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n453), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n285), .A2(KEYINPUT65), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G183gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G190gat), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AOI211_X1 g274(.A(KEYINPUT66), .B(G190gat), .C1(new_n470), .C2(new_n472), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT67), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n451), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n468), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT65), .B(G183gat), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT66), .B1(new_n481), .B2(G190gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n473), .A2(new_n469), .A3(new_n474), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n462), .B1(new_n484), .B2(KEYINPUT67), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n467), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(KEYINPUT27), .ZN(new_n487));
  OR2_X1    g286(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n488));
  AOI211_X1 g287(.A(KEYINPUT28), .B(G190gat), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G183gat), .Z(new_n490));
  OAI21_X1  g289(.A(KEYINPUT28), .B1(new_n490), .B2(G190gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(G183gat), .A2(G190gat), .ZN(new_n492));
  OR3_X1    g291(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n461), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n450), .B1(new_n486), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n285), .A2(new_n474), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(new_n461), .A3(new_n460), .A4(new_n458), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n465), .B1(new_n504), .B2(new_n451), .ZN(new_n505));
  INV_X1    g304(.A(new_n466), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT67), .B(new_n468), .C1(new_n475), .C2(new_n476), .ZN(new_n508));
  INV_X1    g307(.A(new_n462), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT25), .B1(new_n484), .B2(KEYINPUT67), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n497), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n448), .A3(new_n449), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT32), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT72), .B(G71gat), .ZN(new_n521));
  INV_X1    g320(.A(G99gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G43gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  NAND3_X1  g324(.A1(new_n518), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n525), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n517), .B(KEYINPUT32), .C1(new_n519), .C2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n498), .A2(new_n514), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n515), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n531), .B2(KEYINPUT73), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n516), .B1(new_n498), .B2(new_n514), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT73), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT34), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n526), .B(new_n528), .C1(new_n532), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(KEYINPUT73), .A3(new_n529), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT34), .B1(new_n533), .B2(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n528), .A4(new_n526), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n528), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT75), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AND4_X1   g348(.A1(new_n420), .A2(new_n543), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551));
  INV_X1    g350(.A(G226gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n406), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n479), .A2(new_n485), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n497), .B1(new_n555), .B2(new_n507), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n556), .B2(KEYINPUT29), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n556), .B2(new_n554), .ZN(new_n559));
  INV_X1    g358(.A(new_n392), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n512), .A2(new_n513), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT76), .A3(new_n553), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n557), .A2(new_n559), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n553), .B1(new_n561), .B2(new_n402), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n556), .A2(new_n554), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n392), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G8gat), .B(G36gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G64gat), .B(G92gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n563), .A2(new_n566), .A3(KEYINPUT77), .A4(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT35), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n563), .A2(new_n566), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n577));
  INV_X1    g376(.A(new_n569), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n574), .B(new_n575), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n383), .B(new_n446), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT5), .ZN(new_n584));
  NAND2_X1  g383(.A1(G225gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n396), .A2(new_n384), .A3(new_n398), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT3), .B1(new_n380), .B2(new_n382), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n446), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n450), .A2(new_n401), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT4), .ZN(new_n595));
  INV_X1    g394(.A(new_n446), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n596), .B2(new_n383), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n591), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n587), .B1(new_n599), .B2(KEYINPUT5), .ZN(new_n600));
  INV_X1    g399(.A(new_n586), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n590), .A2(KEYINPUT5), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n450), .A2(new_n401), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n596), .A2(new_n383), .A3(new_n595), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n603), .A2(new_n592), .B1(KEYINPUT83), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT83), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n596), .A2(new_n383), .A3(new_n606), .A4(new_n595), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n602), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT87), .B1(new_n600), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n610));
  XNOR2_X1  g409(.A(G57gat), .B(G85gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G1gat), .B(G29gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(KEYINPUT5), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n448), .A2(new_n449), .B1(new_n399), .B2(new_n400), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n597), .B1(new_n616), .B2(new_n593), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n617), .B2(new_n591), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n604), .A2(KEYINPUT83), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(new_n607), .C1(new_n616), .C2(new_n593), .ZN(new_n620));
  INV_X1    g419(.A(new_n602), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT87), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n587), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n614), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n618), .A2(new_n622), .A3(new_n587), .ZN(new_n626));
  INV_X1    g425(.A(new_n614), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT6), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n600), .A2(new_n608), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n614), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT89), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n618), .A2(new_n622), .A3(new_n614), .A4(new_n587), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT6), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n582), .B1(new_n629), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n550), .A2(new_n551), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n628), .B(new_n633), .ZN(new_n639));
  INV_X1    g438(.A(new_n581), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n640), .A2(new_n579), .B1(new_n572), .B2(new_n573), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n543), .A2(new_n420), .A3(new_n546), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT35), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n625), .A2(new_n628), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n631), .A2(new_n635), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n641), .B(new_n575), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n543), .A2(new_n420), .A3(new_n547), .A4(new_n549), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT90), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n638), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n543), .B2(new_n546), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n543), .A2(new_n547), .A3(new_n549), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n651), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n574), .B1(new_n580), .B2(new_n581), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n583), .A2(new_n601), .ZN(new_n656));
  OAI211_X1 g455(.A(KEYINPUT39), .B(new_n656), .C1(new_n599), .C2(new_n601), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n658), .B(new_n586), .C1(new_n617), .C2(new_n591), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n659), .A2(KEYINPUT86), .A3(new_n627), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT86), .B1(new_n659), .B2(new_n627), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n657), .B(KEYINPUT40), .C1(new_n660), .C2(new_n661), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n655), .A2(new_n664), .A3(new_n625), .A4(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT76), .B1(new_n561), .B2(new_n553), .ZN(new_n667));
  AOI211_X1 g466(.A(new_n558), .B(new_n554), .C1(new_n512), .C2(new_n513), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n669), .A2(KEYINPUT88), .A3(new_n392), .A4(new_n557), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n557), .A2(new_n559), .A3(new_n392), .A4(new_n562), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT88), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n560), .B1(new_n564), .B2(new_n565), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT37), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT37), .ZN(new_n677));
  AOI211_X1 g476(.A(KEYINPUT38), .B(new_n578), .C1(new_n576), .C2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n576), .A2(new_n677), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n563), .A2(new_n566), .A3(KEYINPUT37), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n569), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT38), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n636), .A2(new_n679), .A3(new_n683), .A4(new_n629), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n576), .A2(new_n578), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n666), .B(new_n420), .C1(new_n684), .C2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n420), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n642), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n654), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n650), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n325), .A2(new_n284), .A3(new_n326), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n280), .A2(new_n283), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n323), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT93), .ZN(new_n696));
  NAND2_X1  g495(.A1(G229gat), .A2(G233gat), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT18), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n693), .B(new_n323), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n697), .B(KEYINPUT13), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n692), .A2(new_n694), .A3(new_n697), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT18), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT93), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n698), .A2(new_n701), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n707));
  XNOR2_X1  g506(.A(G169gat), .B(G197gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(G113gat), .B(G141gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT92), .B(KEYINPUT12), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n706), .A2(new_n713), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n691), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT94), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n691), .A2(KEYINPUT94), .A3(new_n717), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n356), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n639), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT105), .B(G1gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1324gat));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n727));
  INV_X1    g526(.A(new_n356), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT94), .B1(new_n691), .B2(new_n717), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n719), .B(new_n716), .C1(new_n650), .C2(new_n690), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n655), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT16), .B(G8gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(G8gat), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n731), .A2(new_n727), .A3(new_n732), .ZN(new_n737));
  OAI211_X1 g536(.A(KEYINPUT106), .B(new_n727), .C1(new_n731), .C2(new_n732), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n735), .A2(new_n736), .A3(new_n737), .A4(new_n738), .ZN(G1325gat));
  AOI21_X1  g538(.A(G15gat), .B1(new_n722), .B2(new_n653), .ZN(new_n740));
  INV_X1    g539(.A(new_n654), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(G15gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n722), .B2(new_n742), .ZN(G1326gat));
  NAND2_X1  g542(.A1(new_n722), .A2(new_n688), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT43), .B(G22gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1327gat));
  NAND2_X1  g545(.A1(new_n720), .A2(new_n721), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n306), .A2(new_n350), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n270), .A2(new_n748), .A3(new_n347), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT107), .Z(new_n750));
  NAND3_X1  g549(.A1(new_n747), .A2(new_n723), .A3(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(KEYINPUT45), .A3(G29gat), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n347), .B1(new_n650), .B2(new_n690), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n306), .A2(KEYINPUT109), .A3(new_n350), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT109), .B1(new_n306), .B2(new_n350), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n270), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n714), .B2(new_n715), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n706), .A2(new_n713), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n706), .A2(new_n713), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(KEYINPUT108), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n756), .A2(new_n723), .A3(new_n760), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n753), .B1(new_n768), .B2(G29gat), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n751), .A2(G29gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n752), .B1(new_n769), .B2(new_n770), .ZN(G1328gat));
  OAI211_X1 g570(.A(new_n314), .B(new_n750), .C1(new_n729), .C2(new_n730), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n641), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n756), .A2(new_n655), .A3(new_n760), .A4(new_n767), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(G36gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n747), .A2(new_n314), .A3(new_n655), .A4(new_n750), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT110), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(G1329gat));
  INV_X1    g580(.A(new_n347), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n691), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n755), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n782), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n784), .A2(new_n760), .A3(new_n785), .A4(new_n767), .ZN(new_n786));
  OAI21_X1  g585(.A(G43gat), .B1(new_n786), .B2(new_n654), .ZN(new_n787));
  INV_X1    g586(.A(G43gat), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n747), .A2(new_n788), .A3(new_n653), .A4(new_n750), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT47), .B1(new_n789), .B2(KEYINPUT111), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n787), .B(new_n789), .C1(KEYINPUT111), .C2(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(G1330gat));
  OAI21_X1  g593(.A(G50gat), .B1(new_n786), .B2(new_n420), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n420), .A2(G50gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n747), .A2(new_n750), .A3(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n796), .B1(new_n795), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(G1331gat));
  AND2_X1   g600(.A1(new_n691), .A2(new_n351), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n271), .A2(new_n767), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n723), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n802), .A2(new_n655), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n808), .A2(KEYINPUT112), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(KEYINPUT112), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n812));
  INV_X1    g611(.A(G64gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n809), .A2(new_n812), .A3(new_n813), .A4(new_n810), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1333gat));
  INV_X1    g616(.A(G71gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n804), .A2(new_n818), .A3(new_n653), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n803), .ZN(new_n820));
  OAI21_X1  g619(.A(G71gat), .B1(new_n820), .B2(new_n654), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n822), .B(new_n823), .ZN(G1334gat));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n688), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g625(.A1(new_n767), .A2(new_n748), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n691), .A2(new_n782), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT51), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n754), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n723), .A3(new_n270), .ZN(new_n833));
  INV_X1    g632(.A(new_n213), .ZN(new_n834));
  INV_X1    g633(.A(new_n756), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n827), .A2(new_n270), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n639), .A2(new_n834), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n833), .A2(new_n834), .B1(new_n837), .B2(new_n838), .ZN(G1336gat));
  INV_X1    g638(.A(new_n836), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n784), .A2(new_n655), .A3(new_n785), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G92gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n641), .A2(G92gat), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n829), .A2(new_n270), .A3(new_n831), .A4(new_n843), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  OR2_X1    g644(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g645(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n847));
  AND4_X1   g646(.A1(new_n846), .A2(new_n842), .A3(new_n847), .A4(new_n844), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n845), .A2(new_n848), .ZN(G1337gat));
  NOR3_X1   g648(.A1(new_n835), .A2(new_n654), .A3(new_n836), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n522), .A3(new_n270), .ZN(new_n851));
  INV_X1    g650(.A(new_n653), .ZN(new_n852));
  OAI22_X1  g651(.A1(new_n850), .A2(new_n522), .B1(new_n851), .B2(new_n852), .ZN(G1338gat));
  INV_X1    g652(.A(G106gat), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n829), .A2(new_n854), .A3(new_n270), .A4(new_n831), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n856), .B2(new_n688), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n756), .A2(new_n858), .A3(new_n688), .A4(new_n840), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n784), .A2(new_n688), .A3(new_n785), .A4(new_n840), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n861), .A3(G106gat), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n860), .A2(G106gat), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n855), .A2(new_n420), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT53), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n863), .A2(new_n866), .ZN(G1339gat));
  OR2_X1    g666(.A1(new_n695), .A2(new_n697), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(KEYINPUT116), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(KEYINPUT116), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n699), .A2(new_n700), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n763), .B1(new_n872), .B2(new_n711), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n268), .B2(new_n269), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n875), .B1(new_n247), .B2(new_n248), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n239), .A2(new_n242), .A3(new_n245), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n256), .A2(KEYINPUT54), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n878), .A3(new_n253), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT55), .A4(new_n253), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n260), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n766), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n347), .B1(new_n874), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n873), .ZN(new_n886));
  INV_X1    g685(.A(new_n883), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n782), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n759), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n351), .A2(new_n268), .A3(new_n269), .A4(new_n766), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n271), .A2(KEYINPUT115), .A3(new_n351), .A4(new_n766), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n543), .A2(new_n546), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n897), .A2(new_n723), .A3(new_n420), .A4(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT117), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(new_n641), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n901), .B(new_n767), .C1(new_n433), .C2(new_n432), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n639), .B1(new_n891), .B2(new_n896), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n641), .A3(new_n550), .ZN(new_n904));
  OAI21_X1  g703(.A(G113gat), .B1(new_n904), .B2(new_n716), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(G1340gat));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n421), .A3(new_n270), .ZN(new_n907));
  OAI21_X1  g706(.A(G120gat), .B1(new_n904), .B2(new_n271), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1341gat));
  INV_X1    g708(.A(G127gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n904), .A2(new_n910), .A3(new_n890), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n901), .A2(new_n748), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n910), .ZN(G1342gat));
  INV_X1    g712(.A(G134gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n655), .A2(new_n347), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n917));
  OAI21_X1  g716(.A(G134gat), .B1(new_n904), .B2(new_n347), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n900), .A2(new_n919), .A3(new_n914), .A4(new_n915), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(G1343gat));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n654), .A2(new_n688), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT120), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n897), .A2(new_n924), .A3(new_n723), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n923), .A2(KEYINPUT120), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n926), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n928), .A2(KEYINPUT121), .A3(new_n903), .A4(new_n924), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n927), .A2(new_n641), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n716), .A2(G141gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n270), .A2(new_n886), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n883), .A2(new_n716), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT119), .B1(new_n874), .B2(new_n936), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n347), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n748), .B1(new_n940), .B2(new_n888), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n894), .A2(new_n895), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n688), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT57), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n759), .B1(new_n885), .B2(new_n888), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n688), .B1(new_n945), .B2(new_n942), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n946), .A2(KEYINPUT57), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n654), .A2(new_n723), .A3(new_n641), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT118), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n944), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G141gat), .B1(new_n950), .B2(new_n716), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n933), .A3(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n931), .ZN(new_n953));
  NOR4_X1   g752(.A1(new_n925), .A2(new_n926), .A3(new_n655), .A4(new_n953), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n950), .A2(new_n766), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(G141gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n956), .B2(new_n933), .ZN(G1344gat));
  NOR2_X1   g756(.A1(new_n365), .A2(KEYINPUT59), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n950), .B2(new_n271), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT123), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n420), .A2(KEYINPUT57), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n354), .A2(new_n716), .A3(new_n355), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n941), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n946), .A2(KEYINPUT57), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n270), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G148gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT59), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n968), .B(new_n958), .C1(new_n950), .C2(new_n271), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n960), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n930), .A2(new_n971), .A3(new_n365), .A4(new_n270), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n927), .A2(new_n365), .A3(new_n641), .A4(new_n929), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT122), .B1(new_n973), .B2(new_n271), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n970), .A2(new_n975), .ZN(G1345gat));
  NOR3_X1   g775(.A1(new_n950), .A2(new_n373), .A3(new_n890), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n930), .A2(new_n748), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(new_n373), .ZN(G1346gat));
  OAI21_X1  g778(.A(G162gat), .B1(new_n950), .B2(new_n347), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n927), .A2(new_n374), .A3(new_n915), .A4(new_n929), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1347gat));
  AOI21_X1  g781(.A(new_n723), .B1(new_n891), .B2(new_n896), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n983), .A2(new_n655), .A3(new_n550), .ZN(new_n984));
  OAI21_X1  g783(.A(G169gat), .B1(new_n984), .B2(new_n716), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n897), .A2(new_n639), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT124), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n643), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(new_n655), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n767), .A2(new_n456), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n985), .B1(new_n991), .B2(new_n992), .ZN(G1348gat));
  NOR3_X1   g792(.A1(new_n984), .A2(new_n457), .A3(new_n271), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n990), .A2(new_n655), .A3(new_n270), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n994), .B1(new_n995), .B2(new_n457), .ZN(G1349gat));
  INV_X1    g795(.A(new_n490), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n990), .A2(new_n997), .A3(new_n655), .A4(new_n748), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n481), .B1(new_n984), .B2(new_n890), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(KEYINPUT60), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT60), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n998), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(G1350gat));
  OAI21_X1  g803(.A(G190gat), .B1(new_n984), .B2(new_n347), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT61), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n990), .A2(new_n474), .A3(new_n655), .A4(new_n782), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(G1351gat));
  AND2_X1   g810(.A1(new_n963), .A2(new_n964), .ZN(new_n1012));
  NOR3_X1   g811(.A1(new_n741), .A2(new_n723), .A3(new_n641), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1014), .A2(new_n717), .ZN(new_n1015));
  XOR2_X1   g814(.A(KEYINPUT126), .B(G197gat), .Z(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n923), .B1(new_n987), .B2(new_n989), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(new_n655), .ZN(new_n1019));
  OR2_X1    g818(.A1(new_n766), .A2(new_n1016), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(G1352gat));
  INV_X1    g820(.A(G204gat), .ZN(new_n1022));
  NAND4_X1  g821(.A1(new_n1018), .A2(new_n1022), .A3(new_n655), .A4(new_n270), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1025));
  AND3_X1   g824(.A1(new_n1012), .A2(new_n270), .A3(new_n1013), .ZN(new_n1026));
  OAI211_X1 g825(.A(new_n1024), .B(new_n1025), .C1(new_n1022), .C2(new_n1026), .ZN(G1353gat));
  NAND4_X1  g826(.A1(new_n1018), .A2(new_n387), .A3(new_n655), .A4(new_n748), .ZN(new_n1028));
  NAND4_X1  g827(.A1(new_n963), .A2(new_n748), .A3(new_n964), .A4(new_n1013), .ZN(new_n1029));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1030));
  XNOR2_X1  g829(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  AOI21_X1  g830(.A(KEYINPUT63), .B1(new_n1031), .B2(G211gat), .ZN(new_n1032));
  NAND4_X1  g831(.A1(new_n1012), .A2(new_n1030), .A3(new_n748), .A4(new_n1013), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1034));
  AND4_X1   g833(.A1(KEYINPUT63), .A2(new_n1033), .A3(G211gat), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1028), .B1(new_n1032), .B2(new_n1035), .ZN(G1354gat));
  AND2_X1   g835(.A1(new_n1014), .A2(new_n782), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n782), .A2(new_n388), .ZN(new_n1038));
  OAI22_X1  g837(.A1(new_n1037), .A2(new_n388), .B1(new_n1019), .B2(new_n1038), .ZN(G1355gat));
endmodule


