//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT66), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT28), .B1(new_n203), .B2(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT26), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n207), .A2(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n206), .B2(KEYINPUT26), .ZN(new_n211));
  OR3_X1    g010(.A1(new_n206), .A2(new_n210), .A3(KEYINPUT26), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n202), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n204), .A2(new_n213), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(KEYINPUT24), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n205), .B1(KEYINPUT23), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  OR3_X1    g025(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n219), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT25), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n225), .A2(KEYINPUT25), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n218), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G113gat), .A2(G120gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g033(.A1(G113gat), .A2(G120gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G134gat), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n237), .A2(G127gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(G127gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(G113gat), .B2(G120gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n235), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n238), .A2(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n236), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n231), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT64), .ZN(new_n248));
  OR3_X1    g047(.A1(new_n246), .A2(KEYINPUT34), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT34), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n246), .A2(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT33), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G15gat), .B(G43gat), .Z(new_n255));
  XNOR2_X1  g054(.A(G71gat), .B(G99gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n251), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n257), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(new_n250), .A3(new_n249), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n252), .A2(KEYINPUT32), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n258), .B2(new_n260), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT35), .ZN(new_n265));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G64gat), .B(G92gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n270), .B1(new_n218), .B2(new_n230), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n218), .A2(new_n270), .A3(new_n230), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT70), .B(KEYINPUT29), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n277));
  INV_X1    g076(.A(G197gat), .ZN(new_n278));
  INV_X1    g077(.A(G204gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n231), .A2(KEYINPUT71), .ZN(new_n286));
  INV_X1    g085(.A(new_n273), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n218), .A2(new_n288), .A3(new_n230), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n276), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n274), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n287), .B1(new_n292), .B2(new_n271), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n287), .A2(KEYINPUT29), .ZN(new_n294));
  INV_X1    g093(.A(new_n289), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n288), .B1(new_n218), .B2(new_n230), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n285), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n269), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n273), .B1(new_n272), .B2(new_n274), .ZN(new_n300));
  INV_X1    g099(.A(new_n294), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(new_n286), .B2(new_n289), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n284), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n276), .A2(new_n285), .A3(new_n290), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n268), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(KEYINPUT30), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n303), .A2(new_n304), .A3(new_n307), .A4(new_n268), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n285), .A2(KEYINPUT29), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314));
  INV_X1    g113(.A(G155gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(KEYINPUT74), .A2(G155gat), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT75), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(G155gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n315), .A2(G162gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(G141gat), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G148gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n323), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n330));
  AND2_X1   g129(.A1(KEYINPUT74), .A2(G155gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(KEYINPUT74), .A2(G155gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n330), .B(KEYINPUT2), .C1(new_n333), .C2(new_n313), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n320), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n323), .B1(new_n336), .B2(KEYINPUT2), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n323), .B(KEYINPUT72), .C1(new_n336), .C2(KEYINPUT2), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n311), .A2(new_n312), .B1(new_n335), .B2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n335), .A2(new_n312), .A3(new_n339), .A4(new_n340), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n284), .B1(new_n344), .B2(new_n275), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n284), .A2(KEYINPUT81), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n282), .A2(KEYINPUT81), .A3(new_n283), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n275), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n312), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n320), .A2(new_n334), .A3(new_n329), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(new_n341), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n347), .ZN(new_n354));
  OAI22_X1  g153(.A1(new_n346), .A2(new_n347), .B1(new_n354), .B2(new_n345), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(G22gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT82), .ZN(new_n358));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT31), .B(G50gat), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n359), .B(new_n360), .Z(new_n361));
  OAI21_X1  g160(.A(new_n357), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n264), .A2(new_n265), .A3(new_n310), .A4(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT3), .B1(new_n352), .B2(new_n341), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n344), .A3(new_n245), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT76), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n335), .A2(new_n339), .A3(new_n340), .A4(new_n244), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n342), .A2(KEYINPUT4), .A3(new_n335), .A4(new_n244), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n368), .A2(new_n371), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n377));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT0), .ZN(new_n379));
  XNOR2_X1  g178(.A(G57gat), .B(G85gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n374), .A2(new_n375), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(KEYINPUT77), .A3(new_n371), .A4(new_n368), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n244), .B1(new_n342), .B2(new_n335), .ZN(new_n388));
  INV_X1    g187(.A(new_n372), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n370), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT5), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n382), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  AOI211_X1 g192(.A(KEYINPUT78), .B(new_n391), .C1(new_n384), .C2(new_n386), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n377), .B(new_n381), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT6), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n377), .B1(new_n393), .B2(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n381), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT85), .B(new_n377), .C1(new_n393), .C2(new_n394), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n395), .A2(KEYINPUT79), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n398), .A2(new_n404), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n402), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n404), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n391), .B1(new_n384), .B2(new_n386), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(new_n382), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n412), .A2(new_n397), .A3(new_n377), .A4(new_n381), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT86), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n366), .B1(new_n409), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n413), .A2(new_n406), .A3(new_n414), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n408), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n310), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT80), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(KEYINPUT80), .A3(new_n310), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n264), .A2(new_n365), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n417), .B1(new_n427), .B2(KEYINPUT35), .ZN(new_n428));
  INV_X1    g227(.A(new_n365), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT80), .B1(new_n420), .B2(new_n310), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n422), .B(new_n309), .C1(new_n419), .C2(new_n408), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n264), .A2(KEYINPUT36), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n264), .A2(KEYINPUT36), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT37), .B1(new_n291), .B2(new_n298), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n268), .B1(new_n303), .B2(new_n304), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n269), .A2(KEYINPUT37), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n438), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n442), .A2(KEYINPUT88), .A3(KEYINPUT38), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n285), .B1(new_n300), .B2(new_n302), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n276), .A2(new_n284), .A3(new_n290), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT37), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT87), .A4(KEYINPUT37), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT38), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n439), .B2(new_n441), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n305), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT88), .B1(new_n442), .B2(KEYINPUT38), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n443), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n416), .A2(new_n455), .A3(new_n408), .A4(new_n407), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n371), .B1(new_n385), .B2(new_n368), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n402), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n388), .A2(new_n389), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT39), .B1(new_n460), .B2(new_n370), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT40), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n310), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n429), .B1(new_n466), .B2(new_n404), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n436), .A2(new_n437), .B1(new_n456), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n432), .A2(KEYINPUT83), .A3(new_n435), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n428), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G43gat), .B(G50gat), .Z(new_n471));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G29gat), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n474), .A2(KEYINPUT14), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G36gat), .ZN(new_n476));
  INV_X1    g275(.A(G36gat), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n474), .B2(KEYINPUT14), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(new_n475), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n472), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT89), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n473), .A2(new_n479), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT17), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT90), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n488), .A2(G1gat), .ZN(new_n489));
  INV_X1    g288(.A(G8gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT16), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n488), .B1(new_n491), .B2(G1gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT92), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n489), .B1(new_n495), .B2(new_n492), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n492), .A2(new_n495), .ZN(new_n497));
  OAI21_X1  g296(.A(G8gat), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n484), .A2(new_n485), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n484), .B2(new_n499), .ZN(new_n504));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT93), .Z(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(KEYINPUT18), .A3(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n507), .B(KEYINPUT94), .Z(new_n508));
  AOI21_X1  g307(.A(KEYINPUT18), .B1(new_n504), .B2(new_n506), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n506), .B(new_n510), .ZN(new_n511));
  OR3_X1    g310(.A1(new_n499), .A2(KEYINPUT96), .A3(new_n484), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n499), .A2(new_n484), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT96), .B1(new_n499), .B2(new_n484), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n509), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G197gat), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT11), .B(G169gat), .Z(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n521), .B(KEYINPUT12), .Z(new_n522));
  NAND2_X1  g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n522), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n524), .A3(new_n516), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n470), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531));
  INV_X1    g330(.A(G85gat), .ZN(new_n532));
  INV_X1    g331(.A(G92gat), .ZN(new_n533));
  AOI22_X1  g332(.A1(KEYINPUT8), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT101), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G99gat), .B(G106gat), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n535), .B(KEYINPUT101), .ZN(new_n540));
  INV_X1    g339(.A(new_n538), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n543), .A2(new_n484), .B1(KEYINPUT41), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n543), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT102), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(KEYINPUT102), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n501), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n545), .B1(new_n549), .B2(new_n487), .ZN(new_n550));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n553));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n552), .B(new_n555), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(KEYINPUT98), .Z(new_n559));
  XOR2_X1   g358(.A(G57gat), .B(G64gat), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(G71gat), .B2(G78gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n562), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n560), .A2(new_n567), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n568), .A2(new_n559), .A3(new_n564), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G127gat), .ZN(new_n576));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n500), .B1(new_n572), .B2(new_n571), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT100), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n315), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n580), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n578), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n543), .B(new_n571), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n543), .A2(KEYINPUT10), .A3(new_n566), .A4(new_n570), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G230gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT103), .Z(new_n592));
  AND2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n586), .A2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G120gat), .B(G148gat), .Z(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT104), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n595), .A2(new_n598), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n557), .A2(new_n585), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT105), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n528), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n420), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n309), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT16), .B(G8gat), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT42), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(G8gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT106), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(G1325gat));
  XOR2_X1   g414(.A(new_n435), .B(KEYINPUT107), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(G15gat), .B1(new_n604), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n264), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n619), .A2(G15gat), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n604), .B2(new_n620), .ZN(G1326gat));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n365), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT43), .B(G22gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(G1327gat));
  OAI21_X1  g423(.A(new_n600), .B1(new_n595), .B2(new_n598), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n625), .A2(new_n585), .A3(new_n557), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT108), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n528), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n474), .A3(new_n606), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT45), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n600), .A2(new_n601), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n526), .A2(new_n584), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT44), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n456), .A2(new_n467), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n634), .A2(new_n432), .A3(new_n435), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n633), .B(new_n556), .C1(new_n635), .C2(new_n428), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT109), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n425), .A2(new_n309), .ZN(new_n638));
  INV_X1    g437(.A(new_n416), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n407), .A2(new_n408), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n638), .B(new_n265), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n430), .A2(new_n431), .A3(new_n425), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(new_n265), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n634), .A2(new_n432), .A3(new_n435), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n557), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT109), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n633), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n637), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT44), .B1(new_n470), .B2(new_n557), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n632), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(new_n606), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n630), .B1(new_n474), .B2(new_n651), .ZN(G1328gat));
  NAND4_X1  g451(.A1(new_n528), .A2(new_n477), .A3(new_n309), .A4(new_n627), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT46), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n477), .B1(new_n650), .B2(new_n309), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT110), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1329gat));
  INV_X1    g457(.A(new_n650), .ZN(new_n659));
  OAI21_X1  g458(.A(G43gat), .B1(new_n659), .B2(new_n617), .ZN(new_n660));
  INV_X1    g459(.A(G43gat), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n628), .A2(new_n661), .A3(new_n264), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n435), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n661), .B1(new_n650), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(KEYINPUT47), .ZN(new_n666));
  OAI22_X1  g465(.A1(new_n663), .A2(KEYINPUT47), .B1(new_n665), .B2(new_n666), .ZN(G1330gat));
  INV_X1    g466(.A(G50gat), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(new_n650), .B2(new_n429), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT111), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n528), .A2(new_n668), .A3(new_n429), .A4(new_n627), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n669), .B2(new_n670), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(KEYINPUT48), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(KEYINPUT112), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT112), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n669), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n674), .A2(KEYINPUT48), .B1(new_n677), .B2(new_n679), .ZN(G1331gat));
  NAND2_X1  g479(.A1(new_n643), .A2(new_n644), .ZN(new_n681));
  NOR4_X1   g480(.A1(new_n526), .A2(new_n631), .A3(new_n584), .A4(new_n556), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n606), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g485(.A1(new_n683), .A2(new_n310), .ZN(new_n687));
  NOR2_X1   g486(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n688));
  AND2_X1   g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n687), .B2(new_n688), .ZN(G1333gat));
  NAND3_X1  g490(.A1(new_n684), .A2(G71gat), .A3(new_n616), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n683), .A2(new_n619), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(G71gat), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g494(.A1(new_n684), .A2(new_n429), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G78gat), .ZN(G1335gat));
  INV_X1    g496(.A(KEYINPUT113), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n526), .A2(new_n585), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n625), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n648), .B2(new_n649), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n702), .B2(new_n420), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(KEYINPUT113), .A3(new_n606), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(G85gat), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n645), .A2(new_n699), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT51), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n645), .A2(KEYINPUT51), .A3(new_n699), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n631), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n532), .A3(new_n606), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n705), .A2(new_n711), .ZN(G1336gat));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n533), .A3(new_n309), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n702), .A2(new_n310), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n533), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g515(.A(G99gat), .B1(new_n702), .B2(new_n617), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n708), .A2(new_n709), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n631), .A2(new_n619), .A3(G99gat), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT114), .Z(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(G1338gat));
  NOR2_X1   g521(.A1(new_n636), .A2(KEYINPUT109), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n646), .B1(new_n645), .B2(new_n633), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n365), .B1(new_n423), .B2(new_n424), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n437), .B1(new_n725), .B2(new_n664), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n469), .A3(new_n634), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n557), .B1(new_n727), .B2(new_n643), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n723), .A2(new_n724), .B1(new_n728), .B2(new_n633), .ZN(new_n729));
  INV_X1    g528(.A(new_n700), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n429), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G106gat), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT53), .B1(new_n732), .B2(KEYINPUT115), .ZN(new_n733));
  INV_X1    g532(.A(G106gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n701), .B2(new_n429), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n365), .A2(G106gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n710), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT116), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n732), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n733), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n365), .B(new_n700), .C1(new_n648), .C2(new_n649), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT115), .B1(new_n744), .B2(new_n734), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n739), .A2(new_n741), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n742), .A2(new_n746), .ZN(G1339gat));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n598), .B1(new_n593), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n590), .A2(new_n592), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n590), .A2(new_n592), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(KEYINPUT54), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n752), .A3(KEYINPUT55), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(KEYINPUT117), .Z(new_n754));
  AND2_X1   g553(.A1(new_n749), .A2(new_n752), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT55), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n600), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n504), .A2(new_n506), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n515), .A2(new_n511), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n521), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n525), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n758), .A2(new_n556), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n758), .A2(new_n526), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT118), .B1(new_n631), .B2(new_n762), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n768), .A3(new_n625), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n765), .B1(new_n770), .B2(new_n557), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n771), .A2(new_n585), .B1(new_n526), .B2(new_n602), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(new_n606), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n638), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n526), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n625), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n585), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g579(.A1(new_n773), .A2(new_n638), .A3(new_n556), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT56), .B1(new_n781), .B2(G134gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n781), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(G134gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT119), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(G1343gat));
  NOR3_X1   g587(.A1(new_n616), .A2(new_n309), .A3(new_n365), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n527), .A2(G141gat), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n606), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n772), .A2(new_n794), .A3(new_n429), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n602), .A2(new_n526), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n758), .A2(new_n526), .B1(new_n763), .B2(new_n625), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n764), .B1(new_n797), .B2(new_n556), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n584), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT57), .B1(new_n799), .B2(new_n365), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n664), .A2(new_n420), .A3(new_n309), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n795), .A2(new_n526), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n793), .B1(new_n802), .B2(G141gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT124), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n802), .A2(new_n805), .A3(G141gat), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n802), .B2(G141gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n791), .B(KEYINPUT122), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(G1344gat));
  AND2_X1   g610(.A1(new_n773), .A2(new_n789), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n324), .A2(new_n325), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n625), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n794), .B1(new_n772), .B2(new_n429), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n584), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n603), .A2(new_n527), .ZN(new_n818));
  AOI211_X1 g617(.A(KEYINPUT57), .B(new_n365), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n625), .A3(new_n801), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n815), .B1(new_n821), .B2(G148gat), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n795), .A2(new_n800), .A3(new_n801), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT59), .B(new_n813), .C1(new_n823), .C2(new_n625), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n814), .B1(new_n822), .B2(new_n824), .ZN(G1345gat));
  NAND3_X1  g624(.A1(new_n812), .A2(new_n333), .A3(new_n585), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n823), .A2(new_n585), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n333), .ZN(G1346gat));
  AOI21_X1  g627(.A(G162gat), .B1(new_n812), .B2(new_n556), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n557), .A2(new_n313), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n823), .B2(new_n830), .ZN(G1347gat));
  NOR3_X1   g630(.A1(new_n606), .A2(new_n425), .A3(new_n310), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n772), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(G169gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n834), .A3(new_n527), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n833), .B(KEYINPUT125), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n526), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n837), .B2(new_n834), .ZN(G1348gat));
  INV_X1    g637(.A(G176gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n839), .A3(new_n625), .ZN(new_n840));
  OAI21_X1  g639(.A(G176gat), .B1(new_n833), .B2(new_n631), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1349gat));
  NOR2_X1   g641(.A1(new_n833), .A2(new_n584), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(G183gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n203), .B2(new_n843), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g645(.A(KEYINPUT126), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n848));
  OAI221_X1 g647(.A(G190gat), .B1(new_n847), .B2(new_n848), .C1(new_n833), .C2(new_n557), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n215), .A3(new_n556), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1351gat));
  NAND2_X1  g652(.A1(new_n772), .A2(new_n429), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n617), .A2(new_n420), .A3(new_n309), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(G197gat), .B1(new_n856), .B2(new_n526), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n816), .A2(new_n819), .A3(new_n855), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n527), .A2(new_n278), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(G1352gat));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n279), .A3(new_n625), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT62), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(KEYINPUT62), .ZN(new_n863));
  NOR4_X1   g662(.A1(new_n816), .A2(new_n819), .A3(new_n631), .A4(new_n855), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n279), .ZN(G1353gat));
  INV_X1    g664(.A(G211gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n856), .A2(new_n866), .A3(new_n585), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n858), .A2(new_n585), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT63), .B1(new_n868), .B2(G211gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(G1354gat));
  INV_X1    g670(.A(G218gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n872), .A3(new_n556), .ZN(new_n873));
  NOR4_X1   g672(.A1(new_n816), .A2(new_n819), .A3(new_n557), .A4(new_n855), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n872), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT127), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1355gat));
endmodule


