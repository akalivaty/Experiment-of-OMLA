

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U322 ( .A(n424), .B(n364), .ZN(n469) );
  INV_X1 U323 ( .A(KEYINPUT81), .ZN(n364) );
  XOR2_X1 U324 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n290) );
  XNOR2_X1 U325 ( .A(n444), .B(KEYINPUT120), .ZN(n445) );
  XNOR2_X1 U326 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U327 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n448) );
  XNOR2_X1 U328 ( .A(n363), .B(n362), .ZN(n424) );
  XNOR2_X1 U329 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U330 ( .A(n308), .B(n307), .Z(n532) );
  XOR2_X1 U331 ( .A(KEYINPUT94), .B(n466), .Z(n516) );
  XNOR2_X1 U332 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U333 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT0), .B(G127GAT), .Z(n337) );
  XOR2_X1 U335 ( .A(G134GAT), .B(G99GAT), .Z(n292) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G190GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(n337), .B(n293), .Z(n295) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U341 ( .A(n296), .B(G120GAT), .Z(n300) );
  XOR2_X1 U342 ( .A(G183GAT), .B(KEYINPUT17), .Z(n298) );
  XNOR2_X1 U343 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n443) );
  XNOR2_X1 U345 ( .A(G113GAT), .B(n443), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n308) );
  XOR2_X1 U347 ( .A(G176GAT), .B(G71GAT), .Z(n302) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G15GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U350 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U353 ( .A(n306), .B(n305), .Z(n307) );
  INV_X1 U354 ( .A(n532), .ZN(n456) );
  XOR2_X1 U355 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n310) );
  XNOR2_X1 U356 ( .A(G218GAT), .B(G106GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U358 ( .A(n311), .B(KEYINPUT22), .Z(n313) );
  XOR2_X1 U359 ( .A(KEYINPUT74), .B(G78GAT), .Z(n410) );
  XNOR2_X1 U360 ( .A(G22GAT), .B(n410), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n330) );
  XOR2_X1 U362 ( .A(KEYINPUT92), .B(KEYINPUT86), .Z(n315) );
  NAND2_X1 U363 ( .A1(G228GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n351) );
  XOR2_X1 U366 ( .A(n316), .B(n351), .Z(n328) );
  XOR2_X1 U367 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n318) );
  XNOR2_X1 U368 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U370 ( .A(n319), .B(G211GAT), .Z(n321) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n438) );
  XOR2_X1 U373 ( .A(KEYINPUT91), .B(KEYINPUT2), .Z(n323) );
  XNOR2_X1 U374 ( .A(KEYINPUT90), .B(KEYINPUT3), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U376 ( .A(n324), .B(G155GAT), .Z(n326) );
  XNOR2_X1 U377 ( .A(G141GAT), .B(G148GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n342) );
  XNOR2_X1 U379 ( .A(n438), .B(n342), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n460) );
  XOR2_X1 U382 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n336) );
  XOR2_X1 U383 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n332) );
  XNOR2_X1 U384 ( .A(G162GAT), .B(KEYINPUT5), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n334) );
  XNOR2_X1 U386 ( .A(G29GAT), .B(G134GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n333), .B(G85GAT), .ZN(n359) );
  XNOR2_X1 U388 ( .A(n334), .B(n359), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G57GAT), .Z(n409) );
  XOR2_X1 U391 ( .A(n337), .B(n409), .Z(n339) );
  NAND2_X1 U392 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n344) );
  XOR2_X1 U395 ( .A(G113GAT), .B(G1GAT), .Z(n397) );
  XNOR2_X1 U396 ( .A(n397), .B(n342), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n466) );
  XOR2_X1 U398 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n346) );
  XNOR2_X1 U399 ( .A(KEYINPUT65), .B(KEYINPUT9), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U401 ( .A(G99GAT), .B(G106GAT), .Z(n404) );
  XOR2_X1 U402 ( .A(n347), .B(n404), .Z(n353) );
  INV_X1 U403 ( .A(KEYINPUT7), .ZN(n350) );
  XNOR2_X1 U404 ( .A(KEYINPUT8), .B(G43GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n290), .B(n348), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n388) );
  XNOR2_X1 U407 ( .A(n388), .B(n351), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n363) );
  XOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT80), .Z(n355) );
  NAND2_X1 U410 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U412 ( .A(n356), .B(KEYINPUT79), .Z(n361) );
  XOR2_X1 U413 ( .A(G92GAT), .B(G218GAT), .Z(n358) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(G190GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n433) );
  XNOR2_X1 U416 ( .A(n359), .B(n433), .ZN(n360) );
  XOR2_X1 U417 ( .A(n361), .B(n360), .Z(n362) );
  INV_X1 U418 ( .A(n469), .ZN(n543) );
  XNOR2_X1 U419 ( .A(n543), .B(KEYINPUT99), .ZN(n366) );
  INV_X1 U420 ( .A(KEYINPUT36), .ZN(n365) );
  XNOR2_X1 U421 ( .A(n366), .B(n365), .ZN(n486) );
  XOR2_X1 U422 ( .A(G78GAT), .B(G211GAT), .Z(n368) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(G127GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n381) );
  XOR2_X1 U425 ( .A(G71GAT), .B(KEYINPUT13), .Z(n401) );
  XOR2_X1 U426 ( .A(KEYINPUT14), .B(n401), .Z(n370) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U429 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n372) );
  XNOR2_X1 U430 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U432 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U433 ( .A(G15GAT), .B(G22GAT), .Z(n386) );
  XOR2_X1 U434 ( .A(G64GAT), .B(G57GAT), .Z(n376) );
  XNOR2_X1 U435 ( .A(G1GAT), .B(G155GAT), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n386), .B(n377), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n578) );
  NAND2_X1 U440 ( .A1(n486), .A2(n578), .ZN(n383) );
  XOR2_X1 U441 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n422) );
  XOR2_X1 U443 ( .A(G197GAT), .B(G29GAT), .Z(n385) );
  XNOR2_X1 U444 ( .A(G36GAT), .B(G50GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U446 ( .A(n387), .B(n386), .Z(n390) );
  XOR2_X1 U447 ( .A(G169GAT), .B(G8GAT), .Z(n439) );
  XNOR2_X1 U448 ( .A(n388), .B(n439), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U450 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n392) );
  NAND2_X1 U451 ( .A1(G229GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U453 ( .A(n394), .B(n393), .Z(n400) );
  XOR2_X1 U454 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n396) );
  XNOR2_X1 U455 ( .A(G141GAT), .B(KEYINPUT30), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U458 ( .A(n400), .B(n399), .Z(n572) );
  XOR2_X1 U459 ( .A(G176GAT), .B(G64GAT), .Z(n436) );
  XOR2_X1 U460 ( .A(n436), .B(n401), .Z(n403) );
  XNOR2_X1 U461 ( .A(G85GAT), .B(G92GAT), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n408) );
  XOR2_X1 U463 ( .A(n404), .B(KEYINPUT32), .Z(n406) );
  NAND2_X1 U464 ( .A1(G230GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U466 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n420) );
  XOR2_X1 U469 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n414) );
  XNOR2_X1 U470 ( .A(G204GAT), .B(G148GAT), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U472 ( .A(KEYINPUT77), .B(KEYINPUT75), .Z(n416) );
  XNOR2_X1 U473 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U475 ( .A(n418), .B(n417), .Z(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n575) );
  NOR2_X1 U477 ( .A1(n572), .A2(n575), .ZN(n421) );
  AND2_X1 U478 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n423), .B(KEYINPUT113), .ZN(n430) );
  INV_X1 U480 ( .A(n578), .ZN(n484) );
  NAND2_X1 U481 ( .A1(n424), .A2(n484), .ZN(n427) );
  XOR2_X1 U482 ( .A(KEYINPUT41), .B(n575), .Z(n559) );
  AND2_X1 U483 ( .A1(n572), .A2(n559), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n425), .B(KEYINPUT46), .ZN(n426) );
  NOR2_X1 U485 ( .A1(n427), .A2(n426), .ZN(n428) );
  XNOR2_X1 U486 ( .A(KEYINPUT47), .B(n428), .ZN(n429) );
  NAND2_X1 U487 ( .A1(n430), .A2(n429), .ZN(n432) );
  XNOR2_X1 U488 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n529) );
  XOR2_X1 U490 ( .A(KEYINPUT95), .B(n433), .Z(n435) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U496 ( .A(n443), .B(n442), .Z(n518) );
  AND2_X1 U497 ( .A1(n529), .A2(n518), .ZN(n446) );
  INV_X1 U498 ( .A(KEYINPUT54), .ZN(n444) );
  NOR2_X1 U499 ( .A1(n516), .A2(n447), .ZN(n569) );
  NAND2_X1 U500 ( .A1(n460), .A2(n569), .ZN(n449) );
  NOR2_X1 U501 ( .A1(n456), .A2(n450), .ZN(n564) );
  NAND2_X1 U502 ( .A1(n564), .A2(n543), .ZN(n454) );
  XOR2_X1 U503 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n452) );
  INV_X1 U504 ( .A(G190GAT), .ZN(n451) );
  XNOR2_X1 U505 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U506 ( .A(n518), .B(KEYINPUT27), .ZN(n462) );
  NAND2_X1 U507 ( .A1(n516), .A2(n462), .ZN(n530) );
  XNOR2_X1 U508 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(n460), .ZN(n534) );
  NOR2_X1 U510 ( .A1(n530), .A2(n534), .ZN(n457) );
  NAND2_X1 U511 ( .A1(n457), .A2(n456), .ZN(n468) );
  NAND2_X1 U512 ( .A1(n532), .A2(n518), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n460), .A2(n458), .ZN(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n459), .Z(n464) );
  NOR2_X1 U515 ( .A1(n460), .A2(n532), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT26), .ZN(n570) );
  NAND2_X1 U517 ( .A1(n570), .A2(n462), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n468), .A2(n467), .ZN(n483) );
  NAND2_X1 U521 ( .A1(n469), .A2(n578), .ZN(n470) );
  XOR2_X1 U522 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  AND2_X1 U523 ( .A1(n483), .A2(n471), .ZN(n504) );
  INV_X1 U524 ( .A(n572), .ZN(n502) );
  NOR2_X1 U525 ( .A1(n575), .A2(n502), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n472), .B(KEYINPUT78), .ZN(n489) );
  NAND2_X1 U527 ( .A1(n504), .A2(n489), .ZN(n473) );
  XOR2_X1 U528 ( .A(KEYINPUT96), .B(n473), .Z(n481) );
  NAND2_X1 U529 ( .A1(n516), .A2(n481), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n481), .A2(n518), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n478) );
  NAND2_X1 U534 ( .A1(n532), .A2(n481), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n480) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT97), .Z(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U538 ( .A1(n481), .A2(n534), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NAND2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT100), .B(n485), .Z(n487) );
  NAND2_X1 U543 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U544 ( .A(n488), .B(KEYINPUT37), .ZN(n515) );
  NAND2_X1 U545 ( .A1(n489), .A2(n515), .ZN(n490) );
  XNOR2_X1 U546 ( .A(n490), .B(KEYINPUT101), .ZN(n491) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(n491), .ZN(n499) );
  NAND2_X1 U548 ( .A1(n516), .A2(n499), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U550 ( .A1(n499), .A2(n518), .ZN(n494) );
  XNOR2_X1 U551 ( .A(n494), .B(KEYINPUT102), .ZN(n495) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U554 ( .A1(n532), .A2(n499), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n499), .A2(n534), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n500), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  NAND2_X1 U560 ( .A1(n559), .A2(n502), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n503), .B(KEYINPUT105), .ZN(n514) );
  AND2_X1 U562 ( .A1(n514), .A2(n504), .ZN(n511) );
  NAND2_X1 U563 ( .A1(n516), .A2(n511), .ZN(n505) );
  XNOR2_X1 U564 ( .A(KEYINPUT42), .B(n505), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U566 ( .A1(n511), .A2(n518), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n507), .B(KEYINPUT106), .ZN(n508) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  XOR2_X1 U569 ( .A(G71GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U570 ( .A1(n511), .A2(n532), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U573 ( .A1(n511), .A2(n534), .ZN(n512) );
  XNOR2_X1 U574 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  AND2_X1 U575 ( .A1(n515), .A2(n514), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n524), .A2(n516), .ZN(n517) );
  XNOR2_X1 U577 ( .A(n517), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n524), .A2(n518), .ZN(n519) );
  XNOR2_X1 U579 ( .A(n519), .B(KEYINPUT108), .ZN(n520) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n522) );
  NAND2_X1 U582 ( .A1(n524), .A2(n532), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n528) );
  XOR2_X1 U586 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n526) );
  NAND2_X1 U587 ( .A1(n524), .A2(n534), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n528), .B(n527), .ZN(G1339GAT) );
  INV_X1 U590 ( .A(n529), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n547) );
  NAND2_X1 U592 ( .A1(n532), .A2(n547), .ZN(n533) );
  NOR2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n544) );
  NAND2_X1 U594 ( .A1(n572), .A2(n544), .ZN(n535) );
  XNOR2_X1 U595 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U597 ( .A1(n544), .A2(n559), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U599 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n542) );
  XOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U602 ( .A1(n544), .A2(n578), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n547), .A2(n570), .ZN(n548) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(n548), .Z(n555) );
  NAND2_X1 U610 ( .A1(n572), .A2(n555), .ZN(n549) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U613 ( .A1(n555), .A2(n559), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n555), .A2(n578), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT119), .Z(n557) );
  INV_X1 U619 ( .A(n424), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n572), .A2(n564), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n564), .A2(n559), .ZN(n561) );
  XOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .Z(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n563) );
  XNOR2_X1 U627 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT123), .Z(n566) );
  NAND2_X1 U630 ( .A1(n564), .A2(n578), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT126), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(n568), .Z(n574) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT125), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U640 ( .A1(n580), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n578), .A2(n580), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n486), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

