//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT88), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(G110), .B(G122), .Z(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G107), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n192), .A2(new_n195), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT4), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT77), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n192), .A2(new_n195), .A3(new_n197), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(G101), .A3(new_n200), .ZN(new_n205));
  XNOR2_X1  g019(.A(G116), .B(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n207));
  INV_X1    g021(.A(G113), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G113), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n211), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n206), .B2(KEYINPUT68), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n204), .A2(new_n205), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n191), .A2(G107), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n194), .A2(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n198), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n198), .B2(new_n218), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(new_n206), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G116), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n224), .A2(new_n226), .A3(KEYINPUT5), .ZN(new_n227));
  OAI21_X1  g041(.A(G113), .B1(new_n224), .B2(KEYINPUT5), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n222), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n220), .A2(new_n221), .A3(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n190), .B1(new_n215), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n190), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n198), .A2(new_n218), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT80), .ZN(new_n234));
  INV_X1    g048(.A(new_n228), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n206), .A2(KEYINPUT5), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n235), .A2(new_n236), .B1(new_n206), .B2(new_n213), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n198), .A2(new_n218), .A3(new_n219), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n202), .A2(G101), .A3(new_n200), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n203), .B2(new_n201), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n212), .A2(new_n214), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n232), .B(new_n239), .C1(new_n241), .C2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n231), .A2(new_n244), .A3(KEYINPUT6), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n247), .B(new_n190), .C1(new_n215), .C2(new_n230), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n231), .A2(new_n244), .A3(KEYINPUT83), .A4(KEYINPUT6), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .A4(G128), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT1), .B1(new_n254), .B2(G146), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n253), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(G128), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n253), .A2(new_n255), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G125), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n264), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT0), .A3(G128), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G125), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G224), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n275), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n251), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT84), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n235), .B1(new_n236), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n227), .A2(KEYINPUT84), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n222), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n198), .A2(new_n218), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT85), .B(new_n222), .C1(new_n283), .C2(new_n284), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OR2_X1    g104(.A1(new_n190), .A2(KEYINPUT8), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n237), .A2(new_n233), .B1(KEYINPUT8), .B2(new_n190), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT86), .B(KEYINPUT7), .Z(new_n294));
  OAI21_X1  g108(.A(new_n275), .B1(new_n277), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n278), .A2(KEYINPUT87), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n277), .B2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n267), .A2(new_n274), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n300), .A3(new_n244), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n281), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n279), .B1(new_n249), .B2(new_n250), .ZN(new_n305));
  NOR4_X1   g119(.A1(new_n305), .A2(G902), .A3(new_n188), .A4(new_n302), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G214), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n254), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT64), .B(G131), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT17), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT64), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT64), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G131), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n311), .A2(new_n312), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n315), .A2(new_n316), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT16), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n324), .B2(G125), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n266), .A2(KEYINPUT74), .A3(G140), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n329), .A2(new_n330), .B1(G125), .B2(new_n324), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n331), .B2(new_n326), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G146), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n252), .B(new_n327), .C1(new_n331), .C2(new_n326), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n313), .A2(KEYINPUT17), .A3(new_n314), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n323), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n266), .A2(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n325), .A2(new_n337), .A3(KEYINPUT75), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT75), .B1(new_n325), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n252), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n252), .B2(new_n331), .ZN(new_n342));
  NAND2_X1  g156(.A1(KEYINPUT18), .A2(G131), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n311), .A2(new_n312), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n313), .A2(KEYINPUT18), .A3(G131), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n191), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n336), .A2(new_n346), .A3(new_n349), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XOR2_X1   g167(.A(KEYINPUT90), .B(G475), .Z(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G475), .ZN(new_n357));
  INV_X1    g171(.A(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n315), .A2(new_n322), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT19), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n339), .B2(new_n340), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n329), .A2(new_n330), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n325), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT19), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n361), .A2(new_n364), .A3(KEYINPUT89), .A4(new_n252), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n361), .A2(new_n252), .A3(new_n364), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT89), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n332), .B2(G146), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n359), .B(new_n365), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n349), .B1(new_n369), .B2(new_n346), .ZN(new_n370));
  INV_X1    g184(.A(new_n352), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n357), .B(new_n358), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n372), .A2(KEYINPUT20), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(KEYINPUT20), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n356), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT9), .B(G234), .Z(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G217), .ZN(new_n378));
  NOR3_X1   g192(.A1(new_n377), .A2(new_n378), .A3(G953), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n225), .A2(KEYINPUT14), .A3(G122), .ZN(new_n381));
  XOR2_X1   g195(.A(G116), .B(G122), .Z(new_n382));
  OAI211_X1 g196(.A(G107), .B(new_n381), .C1(new_n382), .C2(KEYINPUT14), .ZN(new_n383));
  XNOR2_X1  g197(.A(G116), .B(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n194), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n254), .A2(G128), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n387));
  INV_X1    g201(.A(G128), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(G143), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n254), .A2(KEYINPUT91), .A3(G128), .ZN(new_n390));
  AOI211_X1 g204(.A(G134), .B(new_n386), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G134), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n390), .ZN(new_n393));
  INV_X1    g207(.A(new_n386), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n383), .B(new_n385), .C1(new_n391), .C2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n397));
  OAI21_X1  g211(.A(G134), .B1(new_n386), .B2(KEYINPUT13), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n382), .A2(G107), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n385), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n398), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT92), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n396), .B2(new_n403), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n380), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n403), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT92), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n379), .A3(new_n405), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n411), .A3(new_n358), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT93), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(new_n416), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n412), .A2(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n375), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  NAND2_X1  g238(.A1(G234), .A2(G237), .ZN(new_n425));
  INV_X1    g239(.A(G953), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G952), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT21), .B(G898), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(G902), .A3(G953), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n308), .A2(new_n423), .A3(new_n424), .A4(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n378), .B1(G234), .B2(new_n358), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT23), .B1(new_n388), .B2(G119), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n223), .A2(G128), .ZN(new_n439));
  MUX2_X1   g253(.A(new_n438), .B(KEYINPUT23), .S(new_n439), .Z(new_n440));
  AOI22_X1  g254(.A1(new_n333), .A2(new_n334), .B1(G110), .B2(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT24), .B(G110), .Z(new_n442));
  XNOR2_X1  g256(.A(G119), .B(G128), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT73), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  OAI22_X1  g260(.A1(new_n440), .A2(G110), .B1(new_n443), .B2(new_n442), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n341), .A3(new_n333), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT22), .B(G137), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n426), .A2(G221), .A3(G234), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n446), .B2(new_n448), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT25), .B1(new_n456), .B2(new_n358), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT25), .ZN(new_n458));
  NOR4_X1   g272(.A1(new_n454), .A2(new_n455), .A3(new_n458), .A4(G902), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n437), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n437), .A2(G902), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n392), .B2(G137), .ZN(new_n465));
  INV_X1    g279(.A(G137), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(KEYINPUT11), .A3(G134), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n392), .A2(G137), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT65), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(new_n467), .A3(new_n471), .A4(new_n468), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(G131), .A3(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n321), .A2(new_n467), .A3(new_n468), .A4(new_n465), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n273), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n466), .A3(G134), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT66), .B1(new_n466), .B2(G134), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n392), .A2(G137), .ZN(new_n481));
  OAI211_X1 g295(.A(G131), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT69), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n388), .B1(new_n259), .B2(new_n260), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n271), .B1(new_n485), .B2(new_n262), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n483), .B(new_n484), .C1(new_n258), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n474), .A2(new_n482), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT69), .B1(new_n265), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n477), .A2(new_n487), .A3(new_n489), .A4(new_n243), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n309), .A2(G210), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n196), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n492), .B(new_n493), .Z(new_n494));
  AOI21_X1  g308(.A(new_n273), .B1(new_n473), .B2(new_n474), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n263), .A2(new_n264), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n488), .B1(new_n496), .B2(new_n257), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT30), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n477), .A2(new_n487), .A3(new_n489), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n498), .B1(KEYINPUT30), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n490), .B(new_n494), .C1(new_n500), .C2(new_n243), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT31), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(KEYINPUT30), .ZN(new_n503));
  INV_X1    g317(.A(new_n498), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n242), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT31), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n490), .A4(new_n494), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n469), .A2(new_n314), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n317), .B1(new_n469), .B2(KEYINPUT65), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n472), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n512), .A2(new_n273), .B1(new_n265), .B2(new_n488), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n509), .B1(new_n513), .B2(new_n242), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n242), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n514), .B(new_n515), .C1(new_n490), .C2(new_n509), .ZN(new_n516));
  INV_X1    g330(.A(new_n494), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT70), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n516), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n502), .A2(new_n508), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT32), .B1(new_n522), .B2(new_n523), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n516), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n494), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n243), .B1(new_n503), .B2(new_n504), .ZN(new_n530));
  INV_X1    g344(.A(new_n490), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n517), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT71), .B1(new_n516), .B2(new_n517), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n529), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n499), .A2(new_n242), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT72), .A3(new_n490), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n499), .A2(new_n538), .A3(new_n242), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(KEYINPUT28), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(KEYINPUT29), .A3(new_n494), .A4(new_n514), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n358), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n463), .B1(new_n526), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n426), .A2(G227), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT76), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G140), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT10), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT79), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n388), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n257), .B1(new_n551), .B2(new_n271), .ZN(new_n552));
  AND4_X1   g366(.A1(new_n550), .A2(new_n552), .A3(new_n198), .A4(new_n218), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n550), .B1(new_n288), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n265), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(KEYINPUT10), .A3(new_n234), .A4(new_n238), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n204), .A2(new_n205), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n559), .B2(new_n476), .ZN(new_n560));
  AOI211_X1 g374(.A(KEYINPUT78), .B(new_n273), .C1(new_n204), .C2(new_n205), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n555), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n548), .B1(new_n562), .B2(new_n475), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT82), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT12), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n288), .A2(new_n552), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT79), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n288), .A2(new_n550), .A3(new_n552), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n567), .A2(new_n568), .B1(new_n233), .B2(new_n265), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n565), .B1(new_n569), .B2(new_n512), .ZN(new_n570));
  OAI22_X1  g384(.A1(new_n553), .A2(new_n554), .B1(new_n556), .B2(new_n288), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(KEYINPUT12), .A3(new_n475), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT81), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT81), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n575), .A3(new_n572), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT82), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n548), .C1(new_n562), .C2(new_n475), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n564), .A2(new_n574), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n562), .A2(new_n475), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT78), .B1(new_n241), .B2(new_n273), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n559), .A2(new_n558), .A3(new_n476), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(new_n512), .A3(new_n555), .A4(new_n557), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n548), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G469), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n358), .ZN(new_n589));
  NAND2_X1  g403(.A1(G469), .A2(G902), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n584), .A3(new_n548), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n573), .A2(new_n584), .ZN(new_n592));
  OAI211_X1 g406(.A(G469), .B(new_n591), .C1(new_n592), .C2(new_n548), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G221), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n376), .B2(new_n358), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n436), .A2(new_n544), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n522), .A2(new_n358), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n601), .A2(G472), .B1(new_n523), .B2(new_n522), .ZN(new_n602));
  INV_X1    g416(.A(new_n463), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n602), .A2(new_n594), .A3(new_n603), .A4(new_n597), .ZN(new_n604));
  INV_X1    g418(.A(new_n187), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n281), .B2(new_n303), .ZN(new_n606));
  NOR4_X1   g420(.A1(new_n305), .A2(G902), .A3(new_n187), .A4(new_n302), .ZN(new_n607));
  INV_X1    g421(.A(new_n424), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OR2_X1    g424(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n406), .A2(new_n380), .A3(new_n407), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n379), .B1(new_n410), .B2(new_n405), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(KEYINPUT33), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n408), .A2(new_n411), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n615), .A2(G478), .A3(new_n358), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n412), .A2(new_n414), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n369), .A2(new_n346), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n352), .B1(new_n622), .B2(new_n349), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT20), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n357), .A4(new_n358), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n372), .A2(KEYINPUT20), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n355), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT95), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT95), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n621), .B2(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n611), .A2(new_n433), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT34), .B(G104), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  XOR2_X1   g449(.A(new_n355), .B(KEYINPUT96), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n625), .A2(new_n626), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n422), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n638), .A2(new_n639), .A3(new_n433), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n611), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n461), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n453), .A2(KEYINPUT36), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n449), .B(new_n646), .Z(new_n647));
  OAI21_X1  g461(.A(new_n460), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n602), .A2(new_n594), .A3(new_n597), .A4(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(new_n435), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  INV_X1    g466(.A(new_n648), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n526), .B2(new_n543), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n428), .B1(new_n432), .B2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n638), .A2(new_n639), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n654), .A2(new_n598), .A3(new_n609), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  XNOR2_X1  g473(.A(new_n656), .B(KEYINPUT39), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n598), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n375), .A2(new_n422), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n307), .B(KEYINPUT38), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n537), .A2(new_n539), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n358), .B1(new_n668), .B2(new_n494), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n494), .B1(new_n530), .B2(new_n531), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n648), .B1(new_n526), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n608), .B1(new_n662), .B2(KEYINPUT40), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n665), .A2(new_n667), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  NOR3_X1   g490(.A1(new_n621), .A2(new_n627), .A3(new_n656), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT97), .B1(new_n610), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT97), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n609), .A2(new_n680), .A3(new_n677), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n654), .A2(new_n679), .A3(new_n598), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  NOR2_X1   g497(.A1(new_n632), .A2(new_n433), .ZN(new_n684));
  INV_X1    g498(.A(new_n578), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n577), .B1(new_n584), .B2(new_n548), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n576), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n575), .B1(new_n570), .B2(new_n572), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n585), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n597), .A3(new_n589), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n610), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n544), .A2(new_n684), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND3_X1  g511(.A1(new_n544), .A2(new_n694), .A3(new_n640), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT98), .B(G116), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G18));
  NAND4_X1  g514(.A1(new_n654), .A2(new_n694), .A3(new_n423), .A4(new_n434), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NOR2_X1   g516(.A1(new_n610), .A2(new_n664), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n601), .A2(G472), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n523), .B(KEYINPUT99), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n502), .A2(new_n508), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n494), .B1(new_n540), .B2(new_n514), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n603), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n693), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n703), .A2(new_n709), .A3(new_n710), .A4(new_n434), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  AND4_X1   g526(.A1(new_n704), .A2(new_n677), .A3(new_n648), .A4(new_n708), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n694), .A2(KEYINPUT100), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n609), .A2(new_n597), .A3(new_n692), .A4(new_n589), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n704), .A2(new_n677), .A3(new_n648), .A4(new_n708), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NOR3_X1   g534(.A1(new_n304), .A2(new_n306), .A3(new_n608), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n594), .A2(new_n597), .A3(new_n677), .A4(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n544), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n522), .A2(new_n523), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT32), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n543), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n603), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n725), .B1(new_n731), .B2(new_n722), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n724), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NAND4_X1  g548(.A1(new_n544), .A2(new_n657), .A3(new_n598), .A4(new_n721), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n375), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n627), .A2(KEYINPUT102), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n619), .A2(new_n620), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT43), .A4(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT101), .B(KEYINPUT43), .Z(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n375), .B2(new_n621), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n704), .A2(new_n726), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n744), .A2(KEYINPUT44), .A3(new_n745), .A4(new_n648), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n721), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT45), .B(new_n591), .C1(new_n592), .C2(new_n548), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  INV_X1    g565(.A(new_n591), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n548), .B1(new_n573), .B2(new_n584), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n754), .A3(G469), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n590), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n589), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT46), .B1(new_n755), .B2(new_n590), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n597), .B(new_n661), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n744), .A2(new_n745), .A3(new_n648), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n746), .A2(KEYINPUT103), .A3(new_n721), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n749), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  OAI21_X1  g579(.A(new_n597), .B1(new_n757), .B2(new_n758), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n597), .B(new_n767), .C1(new_n757), .C2(new_n758), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n730), .ZN(new_n772));
  INV_X1    g586(.A(new_n721), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n773), .A2(new_n678), .A3(new_n603), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT105), .B(G140), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G42));
  INV_X1    g591(.A(new_n656), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n673), .A2(new_n598), .A3(new_n778), .A4(new_n703), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n719), .A2(new_n658), .A3(new_n682), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT52), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n701), .A2(new_n695), .A3(new_n698), .A4(new_n711), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT42), .B1(new_n723), .B2(new_n544), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n731), .A2(new_n722), .A3(new_n725), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n730), .A2(new_n603), .A3(new_n597), .A4(new_n594), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n435), .B1(new_n787), .B2(new_n649), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n308), .A2(new_n424), .A3(new_n434), .ZN(new_n789));
  INV_X1    g603(.A(new_n423), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n627), .B2(new_n740), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n604), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n772), .A2(new_n653), .A3(new_n656), .ZN(new_n794));
  INV_X1    g608(.A(new_n638), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n594), .A2(new_n597), .A3(new_n721), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n639), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n735), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n704), .A2(new_n648), .A3(new_n708), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT107), .B1(new_n722), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT107), .ZN(new_n801));
  INV_X1    g615(.A(new_n799), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n723), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n798), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n786), .A2(new_n793), .A3(new_n797), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(KEYINPUT53), .B1(new_n781), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT100), .B1(new_n694), .B2(new_n713), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n716), .A2(new_n717), .A3(new_n715), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n658), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT108), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n779), .A2(KEYINPUT52), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n719), .A2(new_n812), .A3(new_n658), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n682), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n780), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n695), .A2(new_n711), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n733), .A3(new_n698), .A4(new_n701), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n803), .A2(new_n800), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n793), .A2(new_n797), .A3(new_n821), .A4(new_n735), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n806), .A2(new_n824), .A3(KEYINPUT54), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT109), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n427), .B1(new_n741), .B2(new_n743), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n709), .A3(new_n608), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n666), .A2(new_n710), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT50), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n710), .A2(KEYINPUT112), .A3(new_n721), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT112), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n693), .B2(new_n773), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n834), .A3(new_n802), .A4(new_n828), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n692), .A2(new_n589), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n597), .B1(new_n837), .B2(KEYINPUT111), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(KEYINPUT111), .B2(new_n837), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n769), .A2(new_n839), .A3(new_n770), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n828), .A2(new_n709), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n721), .A3(new_n841), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT50), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n832), .A2(new_n834), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n526), .A2(new_n603), .A3(new_n672), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n375), .A2(new_n740), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n844), .A2(new_n428), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n836), .A2(new_n842), .A3(new_n843), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n544), .A3(new_n828), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n844), .A2(new_n853), .A3(new_n544), .A4(new_n828), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n841), .A2(new_n694), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n850), .A2(new_n857), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n844), .A2(new_n428), .A3(new_n845), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n632), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n848), .A2(new_n849), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n818), .B1(new_n781), .B2(new_n805), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n822), .B1(KEYINPUT110), .B2(new_n786), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT110), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n818), .B1(new_n820), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n817), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n867), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n806), .A2(new_n824), .A3(KEYINPUT109), .A4(KEYINPUT54), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n827), .A2(new_n866), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(G952), .B(new_n426), .C1(new_n875), .C2(KEYINPUT113), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n738), .A2(new_n740), .A3(new_n739), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n667), .A2(new_n608), .A3(new_n596), .A4(new_n877), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n837), .B(KEYINPUT49), .Z(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n845), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT106), .Z(new_n881));
  INV_X1    g695(.A(KEYINPUT113), .ZN(new_n882));
  OAI21_X1  g696(.A(G953), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n876), .A2(new_n881), .A3(new_n883), .ZN(G75));
  XNOR2_X1  g698(.A(new_n279), .B(KEYINPUT55), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n251), .B(KEYINPUT116), .Z(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT117), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n358), .B1(new_n867), .B2(new_n871), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT56), .B(new_n888), .C1(new_n889), .C2(G210), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n817), .A2(new_n868), .A3(new_n870), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n780), .B(new_n815), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n892), .B2(new_n823), .ZN(new_n893));
  OAI211_X1 g707(.A(G210), .B(G902), .C1(new_n891), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n885), .B1(new_n890), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(G210), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n898), .B(new_n358), .C1(new_n867), .C2(new_n871), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n888), .B1(new_n899), .B2(KEYINPUT56), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n895), .A3(new_n887), .ZN(new_n901));
  INV_X1    g715(.A(new_n885), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n426), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n897), .A2(new_n903), .A3(new_n905), .ZN(G51));
  INV_X1    g720(.A(new_n755), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n889), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n590), .A2(KEYINPUT57), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n590), .A2(KEYINPUT57), .ZN(new_n911));
  INV_X1    g725(.A(new_n873), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n872), .B1(new_n867), .B2(new_n871), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n587), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n904), .B1(new_n909), .B2(new_n915), .ZN(G54));
  NAND3_X1  g730(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  INV_X1    g731(.A(new_n623), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n904), .ZN(G60));
  AND2_X1   g735(.A1(new_n615), .A2(new_n618), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n827), .A2(new_n873), .A3(new_n874), .ZN(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT59), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n922), .B(new_n925), .C1(new_n912), .C2(new_n913), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n928), .A3(new_n904), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT60), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n867), .B2(new_n871), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n647), .ZN(new_n934));
  OR2_X1    g748(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n905), .B(new_n935), .C1(new_n932), .C2(new_n456), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT120), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n939), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n934), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(G66));
  OAI21_X1  g757(.A(G953), .B1(new_n430), .B2(new_n276), .ZN(new_n944));
  INV_X1    g758(.A(new_n793), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n782), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n946), .B2(G953), .ZN(new_n947));
  INV_X1    g761(.A(new_n886), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(G898), .B2(new_n426), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  AOI21_X1  g764(.A(new_n426), .B1(G227), .B2(G900), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n426), .A2(KEYINPUT122), .A3(G900), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT122), .B1(new_n426), .B2(G900), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n957), .B(new_n735), .C1(new_n783), .C2(new_n784), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n733), .B2(new_n735), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n810), .A2(new_n682), .A3(new_n813), .ZN(new_n962));
  INV_X1    g776(.A(new_n759), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n544), .A3(new_n703), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n764), .A2(new_n775), .A3(new_n964), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n961), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n955), .B(new_n956), .C1(new_n966), .C2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n361), .A2(new_n364), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n500), .B(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n962), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT123), .B1(new_n785), .B2(new_n798), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n958), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n764), .A2(new_n775), .A3(new_n964), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n426), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n976), .A2(new_n977), .A3(new_n955), .A4(new_n956), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n968), .A2(new_n970), .A3(new_n978), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n970), .B(KEYINPUT121), .Z(new_n980));
  OR4_X1    g794(.A1(new_n787), .A2(new_n660), .A3(new_n773), .A4(new_n791), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n764), .A2(new_n775), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n971), .A2(KEYINPUT62), .A3(new_n675), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  INV_X1    g798(.A(new_n675), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n962), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n982), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n980), .B1(new_n987), .B2(G953), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n953), .B(new_n954), .C1(new_n979), .C2(new_n988), .ZN(new_n989));
  AND4_X1   g803(.A1(new_n952), .A2(new_n979), .A3(new_n951), .A4(new_n988), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(G72));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n966), .B2(new_n946), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n530), .A2(new_n531), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n517), .ZN(new_n997));
  OAI211_X1 g811(.A(KEYINPUT126), .B(new_n905), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n971), .A2(new_n974), .A3(new_n973), .A4(new_n946), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n997), .B1(new_n1000), .B2(new_n993), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n999), .B1(new_n1001), .B2(new_n904), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n997), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1004), .A2(new_n671), .A3(new_n994), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n806), .A2(new_n824), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n946), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n1007), .B(new_n982), .C1(new_n983), .C2(new_n986), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n671), .B1(new_n1008), .B2(new_n994), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1003), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT127), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1003), .A2(new_n1012), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(G57));
endmodule


