

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741;

  XNOR2_X1 U370 ( .A(n528), .B(KEYINPUT39), .ZN(n572) );
  AND2_X1 U371 ( .A1(n527), .A2(n548), .ZN(n528) );
  XNOR2_X1 U372 ( .A(n471), .B(n470), .ZN(n502) );
  XNOR2_X2 U373 ( .A(n435), .B(KEYINPUT92), .ZN(n546) );
  XNOR2_X2 U374 ( .A(n518), .B(n517), .ZN(n710) );
  XOR2_X2 U375 ( .A(n530), .B(KEYINPUT41), .Z(n659) );
  NOR2_X1 U376 ( .A1(n736), .A2(n741), .ZN(n542) );
  NOR2_X1 U377 ( .A1(n602), .A2(n709), .ZN(n604) );
  NOR2_X1 U378 ( .A1(n618), .A2(n709), .ZN(n620) );
  BUF_X1 U379 ( .A(n594), .Z(n621) );
  XNOR2_X1 U380 ( .A(n378), .B(KEYINPUT0), .ZN(n468) );
  OR2_X1 U381 ( .A1(n550), .A2(n377), .ZN(n378) );
  XNOR2_X1 U382 ( .A(n581), .B(n520), .ZN(n644) );
  BUF_X1 U383 ( .A(n519), .Z(n581) );
  XNOR2_X1 U384 ( .A(n401), .B(n400), .ZN(n631) );
  OR2_X1 U385 ( .A1(n698), .A2(G902), .ZN(n429) );
  XNOR2_X1 U386 ( .A(n522), .B(n521), .ZN(n526) );
  XNOR2_X1 U387 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n521) );
  INV_X1 U388 ( .A(KEYINPUT46), .ZN(n541) );
  AND2_X1 U389 ( .A1(n631), .A2(n632), .ZN(n627) );
  INV_X1 U390 ( .A(KEYINPUT1), .ZN(n430) );
  OR2_X1 U391 ( .A1(n598), .A2(G902), .ZN(n414) );
  XNOR2_X1 U392 ( .A(n439), .B(n394), .ZN(n395) );
  XNOR2_X1 U393 ( .A(n418), .B(n417), .ZN(n424) );
  NOR2_X1 U394 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U395 ( .A(n481), .B(KEYINPUT34), .Z(n349) );
  AND2_X1 U396 ( .A1(n555), .A2(n554), .ZN(n350) );
  AND2_X1 U397 ( .A1(n556), .A2(n350), .ZN(n351) );
  NAND2_X1 U398 ( .A1(n648), .A2(n683), .ZN(n553) );
  NOR2_X1 U399 ( .A1(G953), .A2(G237), .ZN(n441) );
  AND2_X1 U400 ( .A1(n589), .A2(n588), .ZN(n593) );
  INV_X1 U401 ( .A(KEYINPUT48), .ZN(n570) );
  XNOR2_X1 U402 ( .A(n422), .B(KEYINPUT79), .ZN(n394) );
  XNOR2_X1 U403 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U404 ( .A1(n365), .A2(n590), .ZN(n368) );
  OR2_X1 U405 ( .A1(n519), .A2(n643), .ZN(n562) );
  XNOR2_X1 U406 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U407 ( .A(n368), .B(n367), .ZN(n519) );
  INV_X1 U408 ( .A(n544), .ZN(n485) );
  XNOR2_X1 U409 ( .A(n452), .B(n451), .ZN(n484) );
  BUF_X1 U410 ( .A(n695), .Z(n705) );
  NOR2_X1 U411 ( .A1(n464), .A2(n483), .ZN(n689) );
  INV_X1 U412 ( .A(KEYINPUT63), .ZN(n603) );
  NOR2_X1 U413 ( .A1(n612), .A2(n709), .ZN(n613) );
  XNOR2_X2 U414 ( .A(G143), .B(G128), .ZN(n454) );
  XNOR2_X1 U415 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n454), .B(n352), .ZN(n723) );
  XNOR2_X1 U417 ( .A(KEYINPUT69), .B(G101), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n723), .B(n353), .ZN(n425) );
  XNOR2_X1 U419 ( .A(KEYINPUT3), .B(G119), .ZN(n716) );
  XNOR2_X1 U420 ( .A(n425), .B(n716), .ZN(n411) );
  INV_X2 U421 ( .A(G953), .ZN(n419) );
  NAND2_X1 U422 ( .A1(n419), .A2(G224), .ZN(n354) );
  XNOR2_X1 U423 ( .A(n354), .B(KEYINPUT85), .ZN(n358) );
  INV_X1 U424 ( .A(G146), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n355), .B(G125), .ZN(n390) );
  XNOR2_X1 U426 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n356) );
  XNOR2_X1 U427 ( .A(n390), .B(n356), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n363) );
  XNOR2_X1 U429 ( .A(G122), .B(G113), .ZN(n359) );
  INV_X1 U430 ( .A(G104), .ZN(n415) );
  XNOR2_X1 U431 ( .A(n359), .B(n415), .ZN(n446) );
  INV_X1 U432 ( .A(n446), .ZN(n362) );
  XNOR2_X1 U433 ( .A(G116), .B(G107), .ZN(n458) );
  XNOR2_X1 U434 ( .A(KEYINPUT16), .B(G110), .ZN(n360) );
  XNOR2_X1 U435 ( .A(n458), .B(n360), .ZN(n361) );
  XNOR2_X1 U436 ( .A(n362), .B(n361), .ZN(n718) );
  XNOR2_X1 U437 ( .A(n363), .B(n718), .ZN(n364) );
  XNOR2_X1 U438 ( .A(n411), .B(n364), .ZN(n615) );
  INV_X1 U439 ( .A(n615), .ZN(n365) );
  XNOR2_X1 U440 ( .A(G902), .B(KEYINPUT15), .ZN(n590) );
  INV_X1 U441 ( .A(G902), .ZN(n450) );
  INV_X1 U442 ( .A(G237), .ZN(n366) );
  NAND2_X1 U443 ( .A1(n450), .A2(n366), .ZN(n369) );
  NAND2_X1 U444 ( .A1(n369), .A2(G210), .ZN(n367) );
  NAND2_X1 U445 ( .A1(n369), .A2(G214), .ZN(n370) );
  XNOR2_X1 U446 ( .A(n370), .B(KEYINPUT87), .ZN(n643) );
  INV_X1 U447 ( .A(KEYINPUT19), .ZN(n371) );
  XNOR2_X1 U448 ( .A(n562), .B(n371), .ZN(n550) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n372) );
  XNOR2_X1 U450 ( .A(n372), .B(KEYINPUT14), .ZN(n625) );
  NOR2_X1 U451 ( .A1(G902), .A2(n419), .ZN(n374) );
  NOR2_X1 U452 ( .A1(G953), .A2(G952), .ZN(n373) );
  NOR2_X1 U453 ( .A1(n374), .A2(n373), .ZN(n375) );
  NAND2_X1 U454 ( .A1(n625), .A2(n375), .ZN(n523) );
  AND2_X1 U455 ( .A1(G953), .A2(G898), .ZN(n376) );
  OR2_X1 U456 ( .A1(n523), .A2(n376), .ZN(n377) );
  XNOR2_X1 U457 ( .A(KEYINPUT89), .B(G140), .ZN(n380) );
  XNOR2_X1 U458 ( .A(G128), .B(G119), .ZN(n379) );
  XNOR2_X1 U459 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U460 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n382) );
  XNOR2_X1 U461 ( .A(G137), .B(KEYINPUT90), .ZN(n381) );
  XNOR2_X1 U462 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U463 ( .A(n384), .B(n383), .ZN(n387) );
  NAND2_X1 U464 ( .A1(G234), .A2(n419), .ZN(n385) );
  XOR2_X1 U465 ( .A(KEYINPUT8), .B(n385), .Z(n453) );
  NAND2_X1 U466 ( .A1(G221), .A2(n453), .ZN(n386) );
  XNOR2_X1 U467 ( .A(n387), .B(n386), .ZN(n396) );
  INV_X1 U468 ( .A(n390), .ZN(n388) );
  NAND2_X1 U469 ( .A1(n388), .A2(KEYINPUT10), .ZN(n392) );
  INV_X1 U470 ( .A(KEYINPUT10), .ZN(n389) );
  NAND2_X1 U471 ( .A1(n390), .A2(n389), .ZN(n391) );
  NAND2_X1 U472 ( .A1(n392), .A2(n391), .ZN(n439) );
  INV_X1 U473 ( .A(G110), .ZN(n393) );
  XNOR2_X1 U474 ( .A(n393), .B(KEYINPUT70), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n396), .B(n395), .ZN(n706) );
  NOR2_X1 U476 ( .A1(n706), .A2(G902), .ZN(n401) );
  XOR2_X1 U477 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n399) );
  NAND2_X1 U478 ( .A1(n590), .A2(G234), .ZN(n397) );
  XNOR2_X1 U479 ( .A(n397), .B(KEYINPUT20), .ZN(n402) );
  NAND2_X1 U480 ( .A1(n402), .A2(G217), .ZN(n398) );
  XNOR2_X1 U481 ( .A(n399), .B(n398), .ZN(n400) );
  AND2_X1 U482 ( .A1(n402), .A2(G221), .ZN(n403) );
  XNOR2_X1 U483 ( .A(n403), .B(KEYINPUT21), .ZN(n632) );
  XOR2_X1 U484 ( .A(G131), .B(KEYINPUT5), .Z(n405) );
  NAND2_X1 U485 ( .A1(n441), .A2(G210), .ZN(n404) );
  XNOR2_X1 U486 ( .A(n405), .B(n404), .ZN(n408) );
  XNOR2_X1 U487 ( .A(G113), .B(G116), .ZN(n406) );
  XNOR2_X1 U488 ( .A(n406), .B(KEYINPUT76), .ZN(n407) );
  XNOR2_X1 U489 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U490 ( .A(G137), .B(G134), .ZN(n726) );
  XNOR2_X1 U491 ( .A(n726), .B(n355), .ZN(n417) );
  XNOR2_X1 U492 ( .A(n409), .B(n417), .ZN(n410) );
  XNOR2_X1 U493 ( .A(n411), .B(n410), .ZN(n598) );
  XNOR2_X1 U494 ( .A(KEYINPUT94), .B(G472), .ZN(n412) );
  XNOR2_X1 U495 ( .A(n412), .B(KEYINPUT74), .ZN(n413) );
  XNOR2_X2 U496 ( .A(n414), .B(n413), .ZN(n634) );
  NAND2_X1 U497 ( .A1(n627), .A2(n634), .ZN(n431) );
  XNOR2_X1 U498 ( .A(G140), .B(G131), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n415), .B(G107), .ZN(n416) );
  XNOR2_X1 U500 ( .A(n440), .B(n416), .ZN(n418) );
  NAND2_X1 U501 ( .A1(n419), .A2(G227), .ZN(n420) );
  XNOR2_X1 U502 ( .A(n420), .B(KEYINPUT88), .ZN(n421) );
  XNOR2_X1 U503 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U504 ( .A(n426), .B(n425), .ZN(n698) );
  XNOR2_X1 U505 ( .A(KEYINPUT73), .B(G469), .ZN(n427) );
  XNOR2_X1 U506 ( .A(n427), .B(KEYINPUT72), .ZN(n428) );
  XNOR2_X1 U507 ( .A(n429), .B(n428), .ZN(n434) );
  XNOR2_X1 U508 ( .A(n434), .B(n430), .ZN(n626) );
  INV_X1 U509 ( .A(n626), .ZN(n577) );
  OR2_X1 U510 ( .A1(n431), .A2(n577), .ZN(n638) );
  OR2_X1 U511 ( .A1(n468), .A2(n638), .ZN(n433) );
  XOR2_X1 U512 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n432) );
  XNOR2_X1 U513 ( .A(n433), .B(n432), .ZN(n690) );
  INV_X1 U514 ( .A(n690), .ZN(n438) );
  INV_X1 U515 ( .A(n434), .ZN(n538) );
  NAND2_X1 U516 ( .A1(n627), .A2(n538), .ZN(n435) );
  OR2_X1 U517 ( .A1(n468), .A2(n546), .ZN(n436) );
  XNOR2_X1 U518 ( .A(n436), .B(KEYINPUT93), .ZN(n437) );
  INV_X1 U519 ( .A(n634), .ZN(n535) );
  NAND2_X1 U520 ( .A1(n437), .A2(n535), .ZN(n671) );
  NAND2_X1 U521 ( .A1(n438), .A2(n671), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n439), .B(n440), .ZN(n724) );
  XOR2_X1 U523 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n443) );
  NAND2_X1 U524 ( .A1(G214), .A2(n441), .ZN(n442) );
  XNOR2_X1 U525 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U526 ( .A(n444), .B(KEYINPUT96), .Z(n448) );
  XNOR2_X1 U527 ( .A(G143), .B(KEYINPUT97), .ZN(n445) );
  XNOR2_X1 U528 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U529 ( .A(n724), .B(n449), .ZN(n609) );
  NAND2_X1 U530 ( .A1(n609), .A2(n450), .ZN(n452) );
  XNOR2_X1 U531 ( .A(KEYINPUT13), .B(G475), .ZN(n451) );
  INV_X1 U532 ( .A(n484), .ZN(n464) );
  NAND2_X1 U533 ( .A1(G217), .A2(n453), .ZN(n456) );
  XNOR2_X1 U534 ( .A(n454), .B(G134), .ZN(n455) );
  XNOR2_X1 U535 ( .A(n456), .B(n455), .ZN(n460) );
  XOR2_X1 U536 ( .A(G122), .B(KEYINPUT9), .Z(n457) );
  XNOR2_X1 U537 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U538 ( .A(n460), .B(n459), .Z(n462) );
  XNOR2_X1 U539 ( .A(KEYINPUT7), .B(KEYINPUT98), .ZN(n461) );
  XNOR2_X1 U540 ( .A(n462), .B(n461), .ZN(n702) );
  NOR2_X1 U541 ( .A1(G902), .A2(n702), .ZN(n463) );
  XNOR2_X1 U542 ( .A(G478), .B(n463), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT99), .B(n689), .ZN(n573) );
  INV_X1 U544 ( .A(n483), .ZN(n465) );
  OR2_X1 U545 ( .A1(n484), .A2(n465), .ZN(n672) );
  NAND2_X1 U546 ( .A1(n573), .A2(n672), .ZN(n648) );
  NAND2_X1 U547 ( .A1(n466), .A2(n648), .ZN(n467) );
  XNOR2_X1 U548 ( .A(n467), .B(KEYINPUT100), .ZN(n474) );
  INV_X1 U549 ( .A(n468), .ZN(n480) );
  AND2_X1 U550 ( .A1(n484), .A2(n483), .ZN(n645) );
  AND2_X1 U551 ( .A1(n645), .A2(n632), .ZN(n469) );
  NAND2_X1 U552 ( .A1(n480), .A2(n469), .ZN(n471) );
  XNOR2_X1 U553 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n470) );
  XNOR2_X1 U554 ( .A(n634), .B(KEYINPUT6), .ZN(n496) );
  AND2_X1 U555 ( .A1(n631), .A2(n577), .ZN(n472) );
  AND2_X1 U556 ( .A1(n496), .A2(n472), .ZN(n473) );
  NAND2_X1 U557 ( .A1(n502), .A2(n473), .ZN(n669) );
  NAND2_X1 U558 ( .A1(n474), .A2(n669), .ZN(n493) );
  NAND2_X1 U559 ( .A1(n626), .A2(n627), .ZN(n475) );
  OR2_X1 U560 ( .A1(n475), .A2(n496), .ZN(n479) );
  XNOR2_X1 U561 ( .A(KEYINPUT101), .B(KEYINPUT33), .ZN(n477) );
  INV_X1 U562 ( .A(KEYINPUT84), .ZN(n476) );
  XNOR2_X1 U563 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U564 ( .A(n479), .B(n478), .ZN(n651) );
  NAND2_X1 U565 ( .A1(n480), .A2(n651), .ZN(n482) );
  INV_X1 U566 ( .A(KEYINPUT77), .ZN(n481) );
  XNOR2_X1 U567 ( .A(n482), .B(n349), .ZN(n486) );
  OR2_X1 U568 ( .A1(n484), .A2(n483), .ZN(n544) );
  NAND2_X1 U569 ( .A1(n486), .A2(n485), .ZN(n489) );
  INV_X1 U570 ( .A(KEYINPUT80), .ZN(n487) );
  XNOR2_X1 U571 ( .A(n487), .B(KEYINPUT35), .ZN(n488) );
  XNOR2_X2 U572 ( .A(n489), .B(n488), .ZN(n606) );
  NAND2_X1 U573 ( .A1(n606), .A2(KEYINPUT44), .ZN(n491) );
  INV_X1 U574 ( .A(KEYINPUT44), .ZN(n507) );
  NAND2_X1 U575 ( .A1(n507), .A2(KEYINPUT66), .ZN(n490) );
  AND2_X1 U576 ( .A1(n491), .A2(n490), .ZN(n492) );
  NOR2_X1 U577 ( .A1(n493), .A2(n492), .ZN(n516) );
  AND2_X1 U578 ( .A1(n507), .A2(KEYINPUT82), .ZN(n494) );
  NAND2_X1 U579 ( .A1(n606), .A2(n494), .ZN(n495) );
  AND2_X1 U580 ( .A1(n495), .A2(KEYINPUT66), .ZN(n504) );
  XNOR2_X1 U581 ( .A(n577), .B(KEYINPUT86), .ZN(n567) );
  INV_X1 U582 ( .A(n496), .ZN(n560) );
  OR2_X1 U583 ( .A1(n560), .A2(n631), .ZN(n497) );
  NOR2_X1 U584 ( .A1(n567), .A2(n497), .ZN(n498) );
  NAND2_X1 U585 ( .A1(n502), .A2(n498), .ZN(n499) );
  XNOR2_X1 U586 ( .A(n499), .B(KEYINPUT32), .ZN(n608) );
  OR2_X1 U587 ( .A1(n631), .A2(n634), .ZN(n500) );
  NOR2_X1 U588 ( .A1(n500), .A2(n626), .ZN(n501) );
  NAND2_X1 U589 ( .A1(n502), .A2(n501), .ZN(n605) );
  AND2_X1 U590 ( .A1(n608), .A2(n605), .ZN(n503) );
  NAND2_X1 U591 ( .A1(n504), .A2(n503), .ZN(n514) );
  INV_X1 U592 ( .A(KEYINPUT82), .ZN(n505) );
  AND2_X1 U593 ( .A1(n505), .A2(KEYINPUT66), .ZN(n506) );
  NAND2_X1 U594 ( .A1(n606), .A2(n506), .ZN(n510) );
  INV_X1 U595 ( .A(KEYINPUT66), .ZN(n508) );
  OR2_X1 U596 ( .A1(n508), .A2(n507), .ZN(n509) );
  AND2_X1 U597 ( .A1(n510), .A2(n509), .ZN(n512) );
  NAND2_X1 U598 ( .A1(n608), .A2(n605), .ZN(n511) );
  NAND2_X1 U599 ( .A1(n512), .A2(n511), .ZN(n513) );
  NAND2_X1 U600 ( .A1(n514), .A2(n513), .ZN(n515) );
  NAND2_X1 U601 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U602 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n517) );
  INV_X1 U603 ( .A(KEYINPUT38), .ZN(n520) );
  NOR2_X1 U604 ( .A1(n644), .A2(n546), .ZN(n527) );
  INV_X1 U605 ( .A(n643), .ZN(n576) );
  NAND2_X1 U606 ( .A1(n634), .A2(n576), .ZN(n522) );
  INV_X1 U607 ( .A(n523), .ZN(n525) );
  NAND2_X1 U608 ( .A1(G953), .A2(G900), .ZN(n524) );
  NAND2_X1 U609 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U610 ( .A1(n526), .A2(n531), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n572), .A2(n672), .ZN(n529) );
  XNOR2_X1 U612 ( .A(n529), .B(KEYINPUT40), .ZN(n736) );
  NOR2_X1 U613 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U614 ( .A1(n645), .A2(n647), .ZN(n530) );
  INV_X1 U615 ( .A(n632), .ZN(n532) );
  NOR2_X1 U616 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U617 ( .A(KEYINPUT71), .B(n533), .ZN(n534) );
  OR2_X1 U618 ( .A1(n631), .A2(n534), .ZN(n558) );
  NOR2_X1 U619 ( .A1(n558), .A2(n535), .ZN(n537) );
  XNOR2_X1 U620 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n536) );
  XNOR2_X1 U621 ( .A(n537), .B(n536), .ZN(n539) );
  NAND2_X1 U622 ( .A1(n539), .A2(n538), .ZN(n551) );
  NOR2_X1 U623 ( .A1(n659), .A2(n551), .ZN(n540) );
  XNOR2_X1 U624 ( .A(n540), .B(KEYINPUT42), .ZN(n741) );
  XNOR2_X1 U625 ( .A(n542), .B(n541), .ZN(n543) );
  INV_X1 U626 ( .A(n543), .ZN(n557) );
  OR2_X1 U627 ( .A1(n544), .A2(n581), .ZN(n545) );
  NOR2_X1 U628 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U629 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U630 ( .A(KEYINPUT105), .B(n549), .Z(n737) );
  XNOR2_X1 U631 ( .A(KEYINPUT78), .B(n737), .ZN(n556) );
  NOR2_X1 U632 ( .A1(n551), .A2(n550), .ZN(n683) );
  NOR2_X1 U633 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n552) );
  XNOR2_X1 U634 ( .A(n553), .B(n552), .ZN(n555) );
  NAND2_X1 U635 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n554) );
  NAND2_X1 U636 ( .A1(n557), .A2(n351), .ZN(n569) );
  NOR2_X1 U637 ( .A1(n558), .A2(n672), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U639 ( .A(n561), .B(KEYINPUT102), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT107), .ZN(n564) );
  INV_X1 U641 ( .A(n562), .ZN(n563) );
  NAND2_X1 U642 ( .A1(n564), .A2(n563), .ZN(n566) );
  XOR2_X1 U643 ( .A(KEYINPUT83), .B(KEYINPUT36), .Z(n565) );
  XNOR2_X1 U644 ( .A(n566), .B(n565), .ZN(n568) );
  NOR2_X1 U645 ( .A1(n568), .A2(n567), .ZN(n693) );
  NOR2_X1 U646 ( .A1(n569), .A2(n693), .ZN(n571) );
  XNOR2_X1 U647 ( .A(n571), .B(n570), .ZN(n586) );
  NOR2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U649 ( .A(KEYINPUT108), .ZN(n574) );
  XNOR2_X1 U650 ( .A(n575), .B(n574), .ZN(n739) );
  NAND2_X1 U651 ( .A1(n577), .A2(n576), .ZN(n578) );
  OR2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT43), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT103), .ZN(n738) );
  INV_X1 U656 ( .A(n738), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n739), .A2(n584), .ZN(n585) );
  NOR2_X2 U658 ( .A1(n586), .A2(n585), .ZN(n731) );
  NAND2_X1 U659 ( .A1(n710), .A2(n731), .ZN(n594) );
  NAND2_X1 U660 ( .A1(KEYINPUT2), .A2(KEYINPUT68), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n594), .A2(n587), .ZN(n589) );
  INV_X1 U662 ( .A(n590), .ZN(n588) );
  INV_X1 U663 ( .A(KEYINPUT2), .ZN(n595) );
  NOR2_X1 U664 ( .A1(n590), .A2(n595), .ZN(n591) );
  NOR2_X1 U665 ( .A1(n591), .A2(KEYINPUT68), .ZN(n592) );
  NOR2_X1 U666 ( .A1(n593), .A2(n592), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n621), .A2(n595), .ZN(n623) );
  NOR2_X2 U668 ( .A1(n596), .A2(n623), .ZN(n695) );
  NAND2_X1 U669 ( .A1(n695), .A2(G472), .ZN(n600) );
  XOR2_X1 U670 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n597) );
  XNOR2_X1 U671 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n600), .B(n599), .ZN(n602) );
  INV_X1 U673 ( .A(G952), .ZN(n601) );
  AND2_X1 U674 ( .A1(n601), .A2(G953), .ZN(n709) );
  XNOR2_X1 U675 ( .A(n604), .B(n603), .ZN(G57) );
  XNOR2_X1 U676 ( .A(n605), .B(G110), .ZN(G12) );
  XNOR2_X1 U677 ( .A(G122), .B(KEYINPUT125), .ZN(n607) );
  XOR2_X1 U678 ( .A(n607), .B(n606), .Z(G24) );
  XNOR2_X1 U679 ( .A(n608), .B(G119), .ZN(G21) );
  NAND2_X1 U680 ( .A1(n695), .A2(G475), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT59), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U684 ( .A1(n695), .A2(G210), .ZN(n617) );
  XOR2_X1 U685 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n619) );
  XNOR2_X1 U689 ( .A(n620), .B(n619), .ZN(G51) );
  INV_X1 U690 ( .A(n621), .ZN(n622) );
  NOR2_X1 U691 ( .A1(n622), .A2(KEYINPUT2), .ZN(n624) );
  NOR2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n664) );
  NAND2_X1 U693 ( .A1(G952), .A2(n625), .ZN(n657) );
  XNOR2_X1 U694 ( .A(KEYINPUT120), .B(KEYINPUT51), .ZN(n641) );
  NOR2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n630) );
  XOR2_X1 U696 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n628) );
  XOR2_X1 U697 ( .A(n628), .B(KEYINPUT118), .Z(n629) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(n637) );
  NOR2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U700 ( .A(KEYINPUT49), .B(n633), .Z(n635) );
  NOR2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U702 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U703 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U704 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X1 U705 ( .A1(n659), .A2(n642), .ZN(n654) );
  NAND2_X1 U706 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U707 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U708 ( .A1(n648), .A2(n647), .ZN(n649) );
  AND2_X1 U709 ( .A1(n650), .A2(n649), .ZN(n652) );
  INV_X1 U710 ( .A(n651), .ZN(n658) );
  NOR2_X1 U711 ( .A1(n652), .A2(n658), .ZN(n653) );
  NOR2_X1 U712 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U713 ( .A(n655), .B(KEYINPUT52), .ZN(n656) );
  NOR2_X1 U714 ( .A1(n657), .A2(n656), .ZN(n661) );
  NOR2_X1 U715 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U716 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U717 ( .A(n662), .B(KEYINPUT121), .ZN(n663) );
  XNOR2_X1 U718 ( .A(n665), .B(KEYINPUT122), .ZN(n666) );
  NAND2_X1 U719 ( .A1(n666), .A2(n419), .ZN(n668) );
  XNOR2_X1 U720 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n667) );
  XNOR2_X1 U721 ( .A(n668), .B(n667), .ZN(G75) );
  XNOR2_X1 U722 ( .A(G101), .B(KEYINPUT110), .ZN(n670) );
  XNOR2_X1 U723 ( .A(n670), .B(n669), .ZN(G3) );
  INV_X1 U724 ( .A(n671), .ZN(n674) );
  INV_X1 U725 ( .A(n672), .ZN(n686) );
  NAND2_X1 U726 ( .A1(n674), .A2(n686), .ZN(n673) );
  XNOR2_X1 U727 ( .A(n673), .B(G104), .ZN(G6) );
  XOR2_X1 U728 ( .A(G107), .B(KEYINPUT27), .Z(n676) );
  NAND2_X1 U729 ( .A1(n674), .A2(n689), .ZN(n675) );
  XNOR2_X1 U730 ( .A(n676), .B(n675), .ZN(n678) );
  XOR2_X1 U731 ( .A(KEYINPUT26), .B(KEYINPUT111), .Z(n677) );
  XNOR2_X1 U732 ( .A(n678), .B(n677), .ZN(G9) );
  XOR2_X1 U733 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n680) );
  NAND2_X1 U734 ( .A1(n683), .A2(n689), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n680), .B(n679), .ZN(n682) );
  XOR2_X1 U736 ( .A(G128), .B(KEYINPUT112), .Z(n681) );
  XNOR2_X1 U737 ( .A(n682), .B(n681), .ZN(G30) );
  NAND2_X1 U738 ( .A1(n683), .A2(n686), .ZN(n684) );
  XNOR2_X1 U739 ( .A(n684), .B(KEYINPUT114), .ZN(n685) );
  XNOR2_X1 U740 ( .A(G146), .B(n685), .ZN(G48) );
  XOR2_X1 U741 ( .A(G113), .B(KEYINPUT115), .Z(n688) );
  NAND2_X1 U742 ( .A1(n690), .A2(n686), .ZN(n687) );
  XNOR2_X1 U743 ( .A(n688), .B(n687), .ZN(G15) );
  NAND2_X1 U744 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U745 ( .A(n691), .B(KEYINPUT116), .ZN(n692) );
  XNOR2_X1 U746 ( .A(G116), .B(n692), .ZN(G18) );
  XNOR2_X1 U747 ( .A(G125), .B(n693), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n694), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U749 ( .A1(n705), .A2(G469), .ZN(n700) );
  XOR2_X1 U750 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n696) );
  XNOR2_X1 U751 ( .A(n696), .B(KEYINPUT124), .ZN(n697) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n709), .A2(n701), .ZN(G54) );
  NAND2_X1 U755 ( .A1(n705), .A2(G478), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n709), .A2(n704), .ZN(G63) );
  NAND2_X1 U758 ( .A1(n705), .A2(G217), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(G66) );
  AND2_X1 U761 ( .A1(n710), .A2(n419), .ZN(n715) );
  INV_X1 U762 ( .A(G898), .ZN(n713) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n711) );
  XOR2_X1 U764 ( .A(KEYINPUT61), .B(n711), .Z(n712) );
  NOR2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n722) );
  XNOR2_X1 U767 ( .A(n716), .B(G101), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U769 ( .A1(G898), .A2(n419), .ZN(n719) );
  NOR2_X1 U770 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U771 ( .A(n722), .B(n721), .Z(G69) );
  XOR2_X1 U772 ( .A(n724), .B(KEYINPUT70), .Z(n725) );
  XNOR2_X1 U773 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U774 ( .A(n723), .B(n727), .ZN(n730) );
  XOR2_X1 U775 ( .A(G227), .B(n730), .Z(n728) );
  NAND2_X1 U776 ( .A1(G900), .A2(n728), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(G953), .ZN(n734) );
  XNOR2_X1 U778 ( .A(n731), .B(n730), .ZN(n732) );
  NAND2_X1 U779 ( .A1(n732), .A2(n419), .ZN(n733) );
  NAND2_X1 U780 ( .A1(n734), .A2(n733), .ZN(G72) );
  XOR2_X1 U781 ( .A(G131), .B(KEYINPUT126), .Z(n735) );
  XNOR2_X1 U782 ( .A(n736), .B(n735), .ZN(G33) );
  XNOR2_X1 U783 ( .A(G143), .B(n737), .ZN(G45) );
  XOR2_X1 U784 ( .A(G140), .B(n738), .Z(G42) );
  XOR2_X1 U785 ( .A(G134), .B(n739), .Z(n740) );
  XNOR2_X1 U786 ( .A(KEYINPUT117), .B(n740), .ZN(G36) );
  XOR2_X1 U787 ( .A(n741), .B(G137), .Z(G39) );
endmodule

