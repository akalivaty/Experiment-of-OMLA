//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n462), .A2(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n467), .A2(G136), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n462), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  INV_X1    g053(.A(G138), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n480), .B(new_n483), .C1(new_n465), .C2(new_n464), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n486), .A2(new_n490), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n482), .B2(new_n484), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT66), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n506), .A2(KEYINPUT67), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n506), .A2(KEYINPUT67), .B1(G75), .B2(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n500), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n505), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n503), .A2(KEYINPUT68), .A3(new_n504), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n518), .A2(KEYINPUT69), .A3(new_n519), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  INV_X1    g101(.A(G51), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n511), .A2(new_n526), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n518), .A2(new_n519), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n511), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n510), .A2(G543), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(G90), .B1(new_n541), .B2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND3_X1  g119(.A1(new_n505), .A2(new_n510), .A3(G81), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n510), .A2(G43), .A3(G543), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT71), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT71), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n518), .A2(G56), .A3(new_n519), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n500), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n547), .A2(new_n548), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT72), .B1(new_n556), .B2(new_n553), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  XNOR2_X1  g140(.A(KEYINPUT74), .B(G65), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n505), .A2(new_n566), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n500), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n513), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n510), .A2(new_n571), .A3(G53), .A4(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n540), .A2(G91), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n568), .A2(new_n573), .A3(new_n574), .ZN(G299));
  AOI21_X1  g150(.A(KEYINPUT75), .B1(new_n525), .B2(new_n532), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n525), .A2(new_n532), .A3(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n500), .B1(new_n536), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n511), .A2(new_n584), .B1(new_n513), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n583), .A2(new_n586), .ZN(G288));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n503), .B2(new_n504), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  INV_X1    g165(.A(G73), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n589), .A2(new_n590), .B1(new_n591), .B2(new_n502), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n505), .A2(new_n590), .A3(G61), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n511), .A2(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n536), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT77), .B(G85), .Z(new_n605));
  AOI22_X1  g180(.A1(new_n540), .A2(new_n605), .B1(new_n541), .B2(G47), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n540), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n511), .B2(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n513), .A2(KEYINPUT78), .ZN(new_n613));
  INV_X1    g188(.A(G54), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(new_n513), .B2(KEYINPUT78), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n609), .A2(new_n612), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n505), .A2(G66), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT79), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n617), .A2(new_n621), .A3(new_n618), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n620), .A2(G651), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n608), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n608), .B1(new_n625), .B2(G868), .ZN(G321));
  AND3_X1   g202(.A1(new_n568), .A2(new_n573), .A3(new_n574), .ZN(new_n628));
  OAI21_X1  g203(.A(KEYINPUT80), .B1(new_n628), .B2(G868), .ZN(new_n629));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n579), .A2(new_n630), .ZN(new_n631));
  MUX2_X1   g206(.A(new_n629), .B(KEYINPUT80), .S(new_n631), .Z(G297));
  XOR2_X1   g207(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n625), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n558), .A2(new_n630), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n624), .A2(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n630), .B2(new_n637), .ZN(G323));
  XOR2_X1   g213(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n639));
  XNOR2_X1  g214(.A(G323), .B(new_n639), .ZN(G282));
  NAND2_X1  g215(.A1(new_n460), .A2(new_n468), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g220(.A1(G123), .A2(new_n473), .B1(new_n467), .B2(G135), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n647), .A2(new_n462), .A3(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n462), .B2(G111), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n649), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n643), .A2(new_n644), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n645), .A2(new_n652), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  INV_X1    g230(.A(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2430), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(KEYINPUT14), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT86), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n666), .B(new_n667), .Z(new_n668));
  OR2_X1    g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(G14), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G401));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  NOR2_X1   g255(.A1(G2072), .A2(G2078), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n442), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n678), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n682), .B(KEYINPUT17), .Z(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n680), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n678), .A3(new_n679), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT18), .Z(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n680), .A3(new_n678), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(new_n644), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT88), .B(G2096), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G227));
  XOR2_X1   g268(.A(G1971), .B(G1976), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT20), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n697), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n695), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n695), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT89), .Z(new_n705));
  XOR2_X1   g280(.A(G1981), .B(G1986), .Z(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n705), .B(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G23), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n583), .A2(new_n586), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT33), .B(G1976), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1971), .ZN(new_n718));
  NAND2_X1  g293(.A1(G166), .A2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G16), .B2(G22), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n712), .A2(G6), .ZN(new_n722));
  INV_X1    g297(.A(G305), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n712), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT32), .B(G1981), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT90), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n720), .A2(new_n718), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n721), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(KEYINPUT34), .ZN(new_n731));
  MUX2_X1   g306(.A(G24), .B(G290), .S(G16), .Z(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(G1986), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(G1986), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n467), .A2(G131), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n473), .A2(G119), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n462), .A2(G107), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n735), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G25), .B(new_n739), .S(G29), .Z(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n733), .A2(new_n734), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n730), .A2(new_n731), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT36), .ZN(new_n746));
  INV_X1    g321(.A(G29), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G32), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n473), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n747), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n747), .B1(new_n758), .B2(G34), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(KEYINPUT92), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(G34), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n759), .B2(KEYINPUT92), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n470), .A2(new_n747), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT30), .B(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n747), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n651), .B2(new_n747), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n765), .B1(KEYINPUT93), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n757), .B(new_n771), .C1(KEYINPUT93), .C2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n747), .A2(G33), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n467), .A2(G139), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(G115), .A2(G2104), .ZN(new_n778));
  INV_X1    g353(.A(G127), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n466), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n777), .B1(G2105), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n773), .B1(new_n781), .B2(new_n747), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n782), .A2(G2072), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n755), .A2(new_n756), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n782), .A2(G2072), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n763), .A2(new_n764), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n747), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n467), .A2(G140), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n473), .A2(G128), .ZN(new_n791));
  OR2_X1    g366(.A1(G104), .A2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n792), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n747), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT91), .B(G2067), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n747), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n747), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G2078), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n772), .A2(new_n787), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n625), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G4), .B2(G16), .ZN(new_n804));
  INV_X1    g379(.A(G1348), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n712), .A2(G5), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G171), .B2(new_n712), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n804), .A2(new_n805), .B1(G1961), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G168), .A2(new_n712), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n712), .B2(G21), .ZN(new_n810));
  INV_X1    g385(.A(G1966), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n747), .A2(G35), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT94), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n747), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n810), .A2(new_n811), .B1(new_n815), .B2(G2090), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n802), .A2(new_n808), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n810), .A2(new_n811), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n804), .A2(new_n805), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n800), .A2(G2078), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n807), .A2(G1961), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n712), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n559), .B2(new_n712), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(G1341), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n817), .B(new_n825), .C1(G1341), .C2(new_n824), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n712), .A2(G20), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT23), .Z(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G299), .B2(G16), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT95), .Z(new_n830));
  INV_X1    g405(.A(G1956), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n815), .A2(G2090), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT96), .Z(new_n836));
  NOR2_X1   g411(.A1(new_n826), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n746), .A2(new_n837), .ZN(G150));
  INV_X1    g413(.A(G150), .ZN(G311));
  XOR2_X1   g414(.A(KEYINPUT97), .B(G93), .Z(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n511), .A2(new_n840), .B1(new_n513), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  INV_X1    g418(.A(G67), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n536), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(new_n845), .B2(G651), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n558), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n549), .A3(new_n554), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n625), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n847), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(G145));
  NAND2_X1  g434(.A1(new_n492), .A2(KEYINPUT98), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n485), .A2(new_n861), .A3(new_n491), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n794), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n781), .B(new_n754), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n739), .B(new_n642), .Z(new_n868));
  AOI22_X1  g443(.A1(G130), .A2(new_n473), .B1(new_n467), .B2(G142), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  INV_X1    g445(.A(G118), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n870), .A2(KEYINPUT99), .B1(new_n871), .B2(G2105), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n872), .B1(KEYINPUT99), .B2(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n868), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n867), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n651), .B(new_n470), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n477), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n866), .A2(new_n876), .A3(new_n875), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n881), .B1(new_n879), .B2(new_n882), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n885), .B2(new_n887), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(G395));
  XOR2_X1   g468(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n637), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n848), .B2(new_n849), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n846), .B1(new_n555), .B2(new_n557), .ZN(new_n898));
  INV_X1    g473(.A(new_n849), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n898), .A2(new_n637), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(G299), .A2(new_n616), .A3(new_n623), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n902), .ZN(new_n905));
  AOI21_X1  g480(.A(G299), .B1(new_n623), .B2(new_n616), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n907), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G288), .B(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G305), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n714), .B(KEYINPUT103), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n723), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(G166), .B(G290), .Z(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n915), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n624), .A2(new_n628), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n903), .B1(new_n920), .B2(new_n902), .ZN(new_n921));
  INV_X1    g496(.A(new_n904), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT41), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n907), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n923), .B(new_n925), .C1(new_n897), .C2(new_n900), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n909), .A2(new_n919), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n919), .B1(new_n909), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n895), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n909), .A2(new_n926), .ZN(new_n930));
  INV_X1    g505(.A(new_n919), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n909), .A2(new_n919), .A3(new_n926), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n894), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(new_n934), .A3(G868), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT105), .B1(new_n847), .B2(new_n630), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n929), .A2(new_n934), .A3(KEYINPUT105), .A4(G868), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(G295));
  AND2_X1   g514(.A1(new_n937), .A2(new_n938), .ZN(G331));
  INV_X1    g515(.A(new_n578), .ZN(new_n941));
  OAI21_X1  g516(.A(G171), .B1(new_n941), .B2(new_n576), .ZN(new_n942));
  NAND2_X1  g517(.A1(G301), .A2(new_n533), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n848), .A2(new_n942), .A3(new_n849), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(G301), .B1(new_n577), .B2(new_n578), .ZN(new_n945));
  INV_X1    g520(.A(new_n943), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n945), .A2(new_n946), .B1(new_n898), .B2(new_n899), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n947), .A3(KEYINPUT106), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n850), .B(new_n949), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n948), .A2(new_n950), .A3(new_n923), .A4(new_n925), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n944), .A3(new_n908), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n953), .B2(new_n931), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n919), .A3(new_n952), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n908), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n948), .B2(new_n950), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n908), .A2(new_n924), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n902), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT107), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n959), .A2(new_n961), .B1(new_n947), .B2(new_n944), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n931), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  AND4_X1   g538(.A1(KEYINPUT43), .A2(new_n963), .A3(new_n884), .A4(new_n955), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT44), .B1(new_n956), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n954), .B2(new_n955), .ZN(new_n968));
  AND4_X1   g543(.A1(new_n967), .A2(new_n963), .A3(new_n884), .A4(new_n955), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(G397));
  AND3_X1   g546(.A1(new_n463), .A2(G40), .A3(new_n469), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT111), .B1(new_n492), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  AOI211_X1 g550(.A(new_n975), .B(G1384), .C1(new_n485), .C2(new_n491), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(G2067), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n496), .B2(G1384), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(new_n484), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n483), .B1(new_n460), .B2(new_n480), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT111), .B(new_n973), .C1(new_n983), .C2(new_n495), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n485), .A2(KEYINPUT66), .A3(new_n491), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT66), .B1(new_n485), .B2(new_n491), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT50), .B(new_n973), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n972), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n978), .B1(new_n990), .B2(new_n805), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT120), .B1(new_n991), .B2(new_n624), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT120), .ZN(new_n993));
  AOI21_X1  g568(.A(G1348), .B1(new_n989), .B2(new_n972), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n993), .B(new_n625), .C1(new_n994), .C2(new_n978), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n979), .A2(KEYINPUT50), .A3(new_n984), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n980), .B(new_n973), .C1(new_n986), .C2(new_n987), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n972), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT117), .B(G1956), .Z(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n973), .B1(new_n986), .B2(new_n987), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT108), .B(G1384), .Z(new_n1004));
  NAND4_X1  g579(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n862), .A4(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT56), .B(G2072), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1003), .A2(new_n972), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(KEYINPUT57), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(KEYINPUT57), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT119), .Z(new_n1013));
  NAND3_X1  g588(.A1(new_n628), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1013), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(G299), .B2(new_n1010), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(KEYINPUT121), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(KEYINPUT121), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1008), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n992), .A2(new_n995), .A3(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1000), .A2(new_n1007), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1022), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1023), .A2(new_n1026), .A3(KEYINPUT61), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT61), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1008), .A2(new_n1028), .A3(new_n1017), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT60), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n994), .B2(new_n978), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n463), .A2(G40), .A3(new_n469), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n985), .B2(new_n988), .ZN(new_n1034));
  OAI221_X1 g609(.A(KEYINPUT60), .B1(G2067), .B2(new_n977), .C1(new_n1034), .C2(G1348), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1035), .A3(new_n625), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n991), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1033), .A2(G1996), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1003), .A2(new_n1005), .A3(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT58), .B(G1341), .Z(new_n1040));
  NAND2_X1  g615(.A1(new_n977), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n558), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT123), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT124), .Z(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1036), .A2(new_n1037), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1025), .B1(new_n1030), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT112), .B(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1002), .A2(G1384), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1033), .B1(new_n498), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n979), .A2(new_n1002), .A3(new_n984), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1966), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n972), .A2(new_n764), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n985), .B2(new_n988), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n533), .B(new_n1053), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n989), .A2(new_n764), .A3(new_n972), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1054), .B1(new_n986), .B2(new_n987), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1056), .A2(new_n1063), .A3(new_n972), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n811), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G168), .A2(new_n1052), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1060), .B(KEYINPUT51), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G2078), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1003), .A2(new_n1069), .A3(new_n972), .A4(new_n1005), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1961), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n990), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1071), .A2(G2078), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1055), .A2(new_n1056), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(G301), .B(KEYINPUT54), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n1053), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1071), .A2(new_n1070), .B1(new_n990), .B2(new_n1073), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n863), .A2(new_n1004), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1002), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n469), .A2(KEYINPUT125), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1087), .A2(G40), .A3(new_n1075), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n463), .B1(KEYINPUT125), .B2(new_n469), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1090), .A2(new_n1005), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1078), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1068), .A2(new_n1079), .A3(new_n1083), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n504), .ZN(new_n1095));
  NOR2_X1   g670(.A1(KEYINPUT5), .A2(G543), .ZN(new_n1096));
  OAI21_X1  g671(.A(G61), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1097), .A2(KEYINPUT76), .B1(G73), .B2(G543), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n500), .B1(new_n1098), .B2(new_n593), .ZN(new_n1099));
  OAI21_X1  g674(.A(G1981), .B1(new_n1099), .B2(new_n598), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n595), .A2(new_n599), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1102), .A3(KEYINPUT113), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n1105));
  NAND3_X1  g680(.A1(G305), .A2(new_n1105), .A3(G1981), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1103), .A2(KEYINPUT114), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n979), .A2(new_n984), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1052), .B1(new_n1112), .B2(new_n972), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(KEYINPUT115), .A3(KEYINPUT49), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT115), .B1(new_n1114), .B2(KEYINPUT49), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1111), .B(new_n1113), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT55), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(G166), .B2(new_n1061), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT55), .B(G8), .C1(new_n509), .C2(new_n515), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G2090), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n996), .A2(new_n997), .A3(new_n972), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1384), .B1(new_n494), .B2(new_n497), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n972), .B(new_n1005), .C1(new_n1125), .C2(KEYINPUT45), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT110), .B(G1971), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1123), .A2(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1122), .B1(new_n1128), .B2(new_n1052), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n714), .A2(G1976), .ZN(new_n1130));
  INV_X1    g705(.A(G1976), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT52), .B1(G288), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1113), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n977), .A2(new_n1053), .A3(new_n1130), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1034), .A2(new_n1123), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1122), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(G8), .A3(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1118), .A2(new_n1129), .A3(new_n1137), .A4(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1094), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1051), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1080), .A2(new_n579), .A3(new_n1053), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1140), .A2(G8), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT116), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1140), .A2(new_n1151), .A3(G8), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1122), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1104), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT115), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1113), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1136), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1061), .B(new_n1122), .C1(new_n1139), .C2(new_n1138), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1080), .A2(KEYINPUT63), .A3(new_n579), .A4(new_n1053), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1148), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1077), .A2(G171), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1143), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1068), .A2(new_n1083), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1068), .A2(KEYINPUT62), .A3(new_n1083), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1165), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1118), .A2(new_n1131), .A3(new_n714), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1102), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1172), .A2(new_n1113), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1145), .A2(new_n1163), .A3(new_n1170), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1085), .A2(new_n1002), .A3(new_n972), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT109), .B1(new_n1175), .B2(G1996), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1175), .A2(KEYINPUT109), .A3(G1996), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n754), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1175), .ZN(new_n1180));
  INV_X1    g755(.A(G2067), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n794), .B(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(G1996), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(new_n754), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n739), .B(new_n741), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1179), .B(new_n1185), .C1(new_n1175), .C2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(G290), .B(G1986), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1187), .B1(new_n1180), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1174), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n739), .A2(new_n742), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT126), .Z(new_n1192));
  NAND3_X1  g767(.A1(new_n1179), .A2(new_n1185), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n795), .A2(new_n1181), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1175), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1175), .A2(G1986), .A3(G290), .ZN(new_n1196));
  XOR2_X1   g771(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1197));
  XNOR2_X1  g772(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1187), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1175), .B1(new_n754), .B2(new_n1182), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT46), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1178), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1203), .A2(KEYINPUT46), .A3(new_n1176), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1200), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT47), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1208));
  AOI211_X1 g783(.A(new_n1195), .B(new_n1199), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1190), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g785(.A1(new_n968), .A2(new_n969), .ZN(new_n1212));
  NOR3_X1   g786(.A1(G229), .A2(G227), .A3(new_n458), .ZN(new_n1213));
  OAI211_X1 g787(.A(new_n676), .B(new_n1213), .C1(new_n885), .C2(new_n887), .ZN(new_n1214));
  NOR2_X1   g788(.A1(new_n1212), .A2(new_n1214), .ZN(G308));
  AND2_X1   g789(.A1(new_n676), .A2(new_n1213), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n886), .A2(new_n888), .ZN(new_n1217));
  OAI211_X1 g791(.A(new_n1216), .B(new_n1217), .C1(new_n968), .C2(new_n969), .ZN(G225));
endmodule


