//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT67), .B(G120gat), .Z(new_n204));
  XOR2_X1   g003(.A(KEYINPUT68), .B(G113gat), .Z(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n203), .A2(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(G127gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n207), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n210), .B(KEYINPUT65), .Z(new_n213));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G127gat), .Z(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(new_n209), .ZN(new_n215));
  XNOR2_X1  g014(.A(G113gat), .B(G120gat), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n213), .A2(new_n215), .B1(KEYINPUT1), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT69), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n212), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G155gat), .B(G162gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT79), .ZN(new_n223));
  INV_X1    g022(.A(G155gat), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT2), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G141gat), .ZN(new_n227));
  INV_X1    g026(.A(G148gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n226), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n231), .A2(new_n222), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(KEYINPUT81), .A3(new_n233), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n239));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n212), .A2(new_n217), .A3(new_n232), .A4(new_n233), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n238), .A2(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n234), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n234), .A2(KEYINPUT3), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n218), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n202), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n218), .A2(new_n234), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n250), .A2(new_n241), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n202), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT39), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT0), .ZN(new_n256));
  XNOR2_X1  g055(.A(G57gat), .B(G85gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(new_n257), .Z(new_n258));
  INV_X1    g057(.A(KEYINPUT39), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n254), .A2(KEYINPUT40), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n202), .B1(new_n251), .B2(KEYINPUT5), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n242), .A2(KEYINPUT82), .A3(new_n240), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n241), .B2(KEYINPUT4), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n238), .A2(new_n239), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n248), .A2(KEYINPUT5), .A3(new_n202), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n262), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n243), .A2(new_n248), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n258), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n270), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT40), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n254), .A2(new_n258), .A3(new_n260), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280));
  INV_X1    g079(.A(G226gat), .ZN(new_n281));
  INV_X1    g080(.A(G233gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G169gat), .ZN(new_n287));
  INV_X1    g086(.A(G176gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT23), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n286), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n293), .A2(new_n294), .B1(new_n285), .B2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT24), .ZN(new_n296));
  INV_X1    g095(.A(G183gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(G190gat), .A3(new_n292), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n291), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT27), .B(G183gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT64), .B1(new_n303), .B2(new_n294), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n286), .A2(KEYINPUT26), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n286), .B1(new_n289), .B2(KEYINPUT26), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n307), .A2(new_n308), .B1(G183gat), .B2(G190gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n284), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT75), .B(new_n284), .C1(new_n311), .C2(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n310), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n283), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT71), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n322), .B1(KEYINPUT22), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n326), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n280), .B1(new_n320), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n320), .A2(new_n280), .A3(new_n332), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n283), .B1(new_n318), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n331), .A3(new_n319), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n339), .A2(new_n340), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n334), .A2(new_n335), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(KEYINPUT30), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n342), .A2(new_n341), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n320), .A2(new_n280), .A3(new_n332), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n333), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n346), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n349), .B(new_n347), .C1(new_n350), .C2(new_n333), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n246), .A2(new_n312), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G228gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(new_n282), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT3), .B1(new_n331), .B2(new_n336), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n358), .B(new_n360), .C1(new_n361), .C2(new_n244), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n236), .A2(new_n237), .ZN(new_n364));
  INV_X1    g163(.A(new_n329), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n326), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n326), .A2(new_n365), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n313), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n368), .B2(KEYINPUT3), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n360), .B1(new_n369), .B2(new_n358), .ZN(new_n370));
  OAI21_X1  g169(.A(G22gat), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n370), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n362), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n376), .B(KEYINPUT84), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(G50gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n377), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n371), .A2(new_n374), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n380), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n371), .A2(new_n374), .A3(new_n381), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n381), .B1(new_n371), .B2(new_n374), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n279), .A2(new_n356), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT37), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n349), .B(new_n389), .C1(new_n350), .C2(new_n333), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n347), .A2(KEYINPUT38), .ZN(new_n391));
  INV_X1    g190(.A(new_n319), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT85), .B(new_n332), .C1(new_n392), .C2(new_n337), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n332), .B1(new_n392), .B2(new_n337), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n393), .B(new_n396), .C1(new_n320), .C2(new_n332), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n391), .B1(new_n397), .B2(KEYINPUT37), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT86), .B1(new_n390), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n265), .A2(new_n263), .B1(new_n238), .B2(new_n239), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n248), .A2(KEYINPUT5), .A3(new_n202), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n401), .A2(new_n402), .B1(new_n403), .B2(new_n202), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT5), .B1(new_n243), .B2(new_n248), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n258), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n275), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n270), .A2(new_n273), .A3(KEYINPUT6), .A4(new_n274), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n408), .A2(new_n353), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n390), .A2(KEYINPUT86), .A3(new_n398), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n400), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n343), .A2(new_n389), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n390), .A2(new_n346), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT38), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n353), .A3(new_n409), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n399), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n411), .B1(new_n419), .B2(new_n412), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n388), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n219), .A2(new_n221), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n311), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n219), .A2(new_n318), .A3(new_n221), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(G227gat), .A3(G233gat), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(KEYINPUT32), .ZN(new_n428));
  XOR2_X1   g227(.A(G15gat), .B(G43gat), .Z(new_n429));
  XNOR2_X1  g228(.A(G71gat), .B(G99gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n431), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n425), .B(KEYINPUT32), .C1(new_n426), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n423), .A2(new_n424), .ZN(new_n436));
  NAND2_X1  g235(.A1(G227gat), .A2(G233gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT34), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n437), .B2(KEYINPUT70), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n440), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n432), .A2(new_n441), .A3(new_n442), .A4(new_n434), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT36), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448));
  INV_X1    g247(.A(new_n352), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n353), .A2(new_n354), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n348), .A2(KEYINPUT78), .A3(new_n352), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n408), .A2(new_n409), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n453), .A2(new_n355), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n387), .A2(new_n383), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n447), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n446), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT35), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n356), .ZN(new_n462));
  INV_X1    g261(.A(new_n453), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n462), .A2(new_n456), .A3(new_n464), .A4(new_n459), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n421), .A2(new_n458), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G113gat), .B(G141gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT11), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(new_n287), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(G197gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT12), .ZN(new_n471));
  INV_X1    g270(.A(G197gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n469), .B(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g275(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n478));
  INV_X1    g277(.A(G1gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT16), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n373), .A2(G15gat), .ZN(new_n481));
  INV_X1    g280(.A(G15gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G22gat), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(G1gat), .B1(new_n481), .B2(new_n483), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n477), .B(new_n478), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n482), .A2(G22gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n373), .A2(G15gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n479), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT90), .A4(G8gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(G29gat), .ZN(new_n499));
  INV_X1    g298(.A(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n499), .A2(new_n500), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G43gat), .A2(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(G43gat), .A2(G50gat), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT15), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n512), .A2(new_n513), .B1(new_n494), .B2(new_n501), .ZN(new_n514));
  OR2_X1    g313(.A1(G43gat), .A2(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n503), .B1(new_n516), .B2(KEYINPUT15), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT91), .B1(new_n493), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n505), .A2(new_n510), .B1(new_n514), .B2(new_n517), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n521), .A2(new_n492), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT92), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n493), .A2(new_n519), .A3(KEYINPUT91), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n522), .B1(new_n521), .B2(new_n492), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n492), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n531), .B(KEYINPUT13), .Z(new_n532));
  AND2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(new_n526), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n511), .A2(KEYINPUT17), .A3(new_n518), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n501), .A2(new_n494), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n515), .A2(new_n513), .A3(new_n506), .ZN(new_n538));
  AND4_X1   g337(.A1(new_n509), .A2(new_n537), .A3(new_n538), .A4(new_n504), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n509), .B1(new_n502), .B2(new_n504), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n535), .A2(new_n541), .A3(new_n492), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n534), .A2(new_n531), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n531), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n476), .B1(new_n533), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n471), .A2(new_n475), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n532), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n549), .A2(new_n550), .A3(new_n545), .A4(new_n546), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n466), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G183gat), .B(G211gat), .Z(new_n554));
  INV_X1    g353(.A(G71gat), .ZN(new_n555));
  INV_X1    g354(.A(G78gat), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT93), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G57gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G64gat), .ZN(new_n567));
  INV_X1    g366(.A(G64gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n568), .A2(G57gat), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n567), .A2(new_n569), .B1(KEYINPUT9), .B2(new_n561), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n563), .A3(new_n557), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n493), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n579), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n582), .B1(new_n580), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n554), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  INV_X1    g387(.A(new_n554), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT8), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n593), .A2(new_n596), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G99gat), .B(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n597), .B2(new_n598), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(new_n602), .A3(new_n596), .A4(new_n600), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n535), .A2(new_n541), .A3(KEYINPUT94), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n511), .B2(new_n518), .ZN(new_n609));
  NAND3_X1  g408(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT95), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n613), .B(new_n610), .C1(new_n521), .C2(new_n607), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n535), .A2(new_n541), .A3(new_n607), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT94), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND4_X1   g419(.A1(new_n608), .A2(new_n615), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n612), .A2(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n622), .B2(new_n608), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT96), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n615), .A2(new_n608), .A3(new_n618), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n619), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n622), .A2(new_n608), .A3(new_n620), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n624), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n630), .A2(new_n631), .A3(new_n627), .A4(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n591), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n560), .A2(new_n564), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n563), .B1(new_n570), .B2(new_n557), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n606), .B(new_n604), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n607), .A2(new_n565), .A3(new_n571), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n606), .A4(new_n604), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n642), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n647), .A2(new_n650), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n637), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n553), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n453), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n479), .ZN(G1324gat));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n462), .ZN(new_n663));
  INV_X1    g462(.A(G8gat), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT42), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  MUX2_X1   g466(.A(KEYINPUT42), .B(new_n665), .S(new_n667), .Z(G1325gat));
  INV_X1    g467(.A(new_n660), .ZN(new_n669));
  AOI21_X1  g468(.A(G15gat), .B1(new_n669), .B2(new_n459), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n447), .A2(G15gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT97), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n669), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n660), .A2(new_n456), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  NOR3_X1   g475(.A1(new_n591), .A2(new_n636), .A3(new_n658), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT98), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n553), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(G29gat), .A3(new_n453), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n421), .A2(new_n458), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n461), .A2(new_n465), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n636), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(KEYINPUT44), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n636), .A2(KEYINPUT99), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n634), .A2(new_n689), .A3(new_n635), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n687), .B1(new_n466), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n591), .A2(new_n552), .A3(new_n658), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n499), .B1(new_n696), .B2(new_n463), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n681), .A2(new_n697), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n679), .A2(G36gat), .A3(new_n462), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n356), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G36gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(G1329gat));
  NAND3_X1  g505(.A1(new_n696), .A2(G43gat), .A3(new_n447), .ZN(new_n707));
  INV_X1    g506(.A(G43gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n679), .B2(new_n446), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n712), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1330gat));
  XNOR2_X1  g513(.A(new_n679), .B(KEYINPUT101), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n456), .A2(G50gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n694), .A2(new_n457), .A3(new_n695), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(G50gat), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT102), .B1(new_n717), .B2(G50gat), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(G50gat), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n679), .A2(KEYINPUT101), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n553), .B2(new_n678), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n716), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n722), .B(new_n726), .C1(new_n727), .C2(new_n719), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n721), .A2(new_n729), .ZN(G1331gat));
  NAND2_X1  g529(.A1(new_n548), .A2(new_n551), .ZN(new_n731));
  INV_X1    g530(.A(new_n658), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n637), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n684), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n453), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n566), .ZN(G1332gat));
  AOI211_X1 g535(.A(new_n462), .B(new_n734), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  XOR2_X1   g538(.A(new_n446), .B(KEYINPUT103), .Z(new_n740));
  NOR2_X1   g539(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n555), .B1(new_n741), .B2(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n447), .A2(G71gat), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n742), .A2(new_n743), .B1(new_n734), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g545(.A1(new_n734), .A2(new_n456), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n556), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n591), .A2(new_n731), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n732), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n694), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n453), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n636), .B1(new_n682), .B2(new_n683), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT51), .B1(new_n754), .B2(new_n749), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n466), .A2(new_n756), .A3(new_n636), .A4(new_n750), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT105), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n463), .A2(new_n597), .A3(new_n658), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT106), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n753), .B1(new_n759), .B2(new_n761), .ZN(G1336gat));
  OAI21_X1  g561(.A(G92gat), .B1(new_n752), .B2(new_n462), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n758), .A2(new_n598), .A3(new_n356), .A4(new_n658), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g565(.A(new_n447), .ZN(new_n767));
  OAI21_X1  g566(.A(G99gat), .B1(new_n752), .B2(new_n767), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n446), .A2(G99gat), .A3(new_n732), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n759), .B2(new_n769), .ZN(G1338gat));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n686), .A2(new_n693), .A3(new_n457), .A4(new_n751), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G106gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n456), .A2(G106gat), .A3(new_n732), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT107), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n755), .B2(new_n757), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n771), .B1(new_n777), .B2(KEYINPUT53), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779));
  AOI211_X1 g578(.A(KEYINPUT108), .B(new_n779), .C1(new_n773), .C2(new_n776), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n755), .B2(new_n757), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n694), .A2(KEYINPUT110), .A3(new_n457), .A4(new_n751), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n772), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT111), .B(new_n784), .C1(new_n788), .C2(G106gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n772), .A2(new_n786), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n772), .A2(new_n786), .ZN(new_n792));
  OAI21_X1  g591(.A(G106gat), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n784), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n781), .B1(new_n789), .B2(new_n795), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n643), .A2(new_n644), .A3(new_n649), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n649), .B1(new_n643), .B2(new_n644), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n656), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n657), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n801), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g606(.A(KEYINPUT112), .B(KEYINPUT55), .C1(new_n798), .C2(new_n801), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810));
  INV_X1    g609(.A(new_n532), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n524), .A2(new_n811), .A3(new_n528), .A4(new_n529), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n534), .A2(new_n542), .ZN(new_n813));
  INV_X1    g612(.A(new_n531), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n810), .B1(new_n816), .B2(new_n470), .ZN(new_n817));
  AOI211_X1 g616(.A(KEYINPUT113), .B(new_n473), .C1(new_n812), .C2(new_n815), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n551), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n809), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n634), .A2(new_n689), .A3(new_n635), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n689), .B1(new_n634), .B2(new_n635), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n691), .A2(KEYINPUT114), .A3(new_n820), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n805), .A2(new_n806), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT112), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n805), .A2(new_n804), .A3(new_n806), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n731), .A3(new_n803), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n551), .B(new_n658), .C1(new_n817), .C2(new_n818), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT115), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n692), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n591), .B1(new_n827), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n591), .A2(new_n552), .A3(new_n636), .A4(new_n732), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT116), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n836), .B1(new_n832), .B2(new_n833), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n691), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n837), .A2(new_n845), .B1(new_n825), .B2(new_n826), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n843), .B(new_n840), .C1(new_n846), .C2(new_n591), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n356), .A2(new_n453), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n460), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n731), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n205), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(G113gat), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n851), .A3(new_n658), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G120gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n204), .B2(new_n858), .ZN(G1341gat));
  NAND3_X1  g659(.A1(new_n850), .A2(new_n851), .A3(new_n591), .ZN(new_n861));
  INV_X1    g660(.A(new_n214), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT118), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  MUX2_X1   g663(.A(new_n863), .B(KEYINPUT118), .S(new_n864), .Z(G1342gat));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n685), .A3(new_n849), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(G134gat), .A3(new_n460), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n866), .B2(new_n460), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n867), .B2(new_n869), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n874), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n876), .B(new_n877), .C1(new_n871), .C2(new_n870), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(new_n878), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n803), .A2(new_n828), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n833), .B1(new_n552), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n636), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n827), .ZN(new_n884));
  INV_X1    g683(.A(new_n591), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n841), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n456), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n842), .A2(new_n847), .A3(new_n457), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n767), .A2(new_n849), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(new_n227), .A3(new_n552), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n447), .A2(new_n456), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n850), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(G141gat), .B1(new_n896), .B2(new_n731), .ZN(new_n897));
  OR3_X1    g696(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n893), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1344gat));
  NAND3_X1  g699(.A1(new_n896), .A2(new_n228), .A3(new_n658), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n892), .A2(new_n732), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(KEYINPUT59), .A3(new_n228), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n840), .B(KEYINPUT122), .Z(new_n906));
  NAND2_X1  g705(.A1(new_n820), .A2(new_n685), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n591), .B1(new_n907), .B2(new_n882), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n887), .B(new_n457), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n732), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n767), .A3(new_n849), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n904), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n901), .B1(new_n903), .B2(new_n913), .ZN(G1345gat));
  OAI21_X1  g713(.A(G155gat), .B1(new_n892), .B2(new_n885), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n896), .A2(new_n224), .A3(new_n591), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n892), .B2(new_n692), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n895), .A2(new_n225), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n866), .B2(new_n919), .ZN(G1347gat));
  NAND2_X1  g719(.A1(new_n356), .A2(new_n453), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n740), .A2(new_n457), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n848), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n287), .A3(new_n552), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n848), .A2(new_n453), .A3(new_n851), .A4(new_n356), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n926), .A2(new_n552), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n927), .B2(new_n287), .ZN(G1348gat));
  OAI21_X1  g727(.A(G176gat), .B1(new_n924), .B2(new_n732), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n658), .A2(new_n288), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n926), .B2(new_n930), .ZN(G1349gat));
  INV_X1    g730(.A(new_n303), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n926), .A2(new_n932), .A3(new_n885), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n297), .B1(new_n923), .B2(new_n591), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g735(.A(new_n294), .B1(new_n923), .B2(new_n685), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT61), .Z(new_n938));
  NOR3_X1   g737(.A1(new_n926), .A2(G190gat), .A3(new_n692), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT123), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1351gat));
  NOR3_X1   g740(.A1(new_n910), .A2(new_n447), .A3(new_n921), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n552), .A2(new_n472), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n848), .A2(new_n453), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n447), .A2(new_n462), .A3(new_n456), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n731), .A3(new_n945), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n942), .A2(new_n943), .B1(new_n946), .B2(new_n472), .ZN(G1352gat));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(new_n945), .ZN(new_n949));
  XOR2_X1   g748(.A(KEYINPUT124), .B(G204gat), .Z(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n732), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n948), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n944), .A2(KEYINPUT62), .A3(new_n945), .A4(new_n952), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n921), .A2(new_n447), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n911), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n951), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT125), .ZN(G1353gat));
  NAND4_X1  g760(.A1(new_n905), .A2(new_n591), .A3(new_n909), .A4(new_n957), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n962), .A2(new_n965), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n962), .A2(G211gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n944), .A2(new_n323), .A3(new_n591), .A4(new_n945), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(KEYINPUT127), .A3(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1354gat));
  AOI21_X1  g775(.A(new_n324), .B1(new_n942), .B2(new_n685), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n949), .A2(G218gat), .A3(new_n692), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n977), .A2(new_n978), .ZN(G1355gat));
endmodule


