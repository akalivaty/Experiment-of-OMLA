

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(KEYINPUT33), .A2(n682), .ZN(n687) );
  NOR2_X1 U554 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U555 ( .A1(n680), .A2(n695), .ZN(n517) );
  AND2_X1 U556 ( .A1(n944), .A2(n747), .ZN(n518) );
  NOR2_X1 U557 ( .A1(n736), .A2(n518), .ZN(n519) );
  OR2_X1 U558 ( .A1(n632), .A2(n757), .ZN(n633) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n658) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n654) );
  XNOR2_X1 U561 ( .A(n659), .B(n658), .ZN(n667) );
  NAND2_X1 U562 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U563 ( .A1(n702), .A2(n597), .ZN(n661) );
  NAND2_X1 U564 ( .A1(G8), .A2(n661), .ZN(n695) );
  AND2_X1 U565 ( .A1(n687), .A2(n686), .ZN(n699) );
  NOR2_X2 U566 ( .A1(G2105), .A2(n525), .ZN(n873) );
  NOR2_X2 U567 ( .A1(G651), .A2(n580), .ZN(n786) );
  INV_X1 U568 ( .A(G2104), .ZN(n525) );
  NAND2_X1 U569 ( .A1(G102), .A2(n873), .ZN(n522) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X2 U571 ( .A(KEYINPUT17), .B(n520), .Z(n870) );
  NAND2_X1 U572 ( .A1(G138), .A2(n870), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n522), .A2(n521), .ZN(n529) );
  INV_X1 U574 ( .A(G2105), .ZN(n524) );
  NOR2_X1 U575 ( .A1(n524), .A2(G2104), .ZN(n523) );
  XNOR2_X2 U576 ( .A(n523), .B(KEYINPUT64), .ZN(n866) );
  NAND2_X1 U577 ( .A1(G126), .A2(n866), .ZN(n527) );
  NOR2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n865) );
  NAND2_X1 U579 ( .A1(G114), .A2(n865), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U581 ( .A1(n529), .A2(n528), .ZN(G164) );
  NAND2_X1 U582 ( .A1(n873), .A2(G101), .ZN(n532) );
  XNOR2_X1 U583 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n530) );
  XNOR2_X1 U584 ( .A(n530), .B(KEYINPUT66), .ZN(n531) );
  XNOR2_X1 U585 ( .A(n532), .B(n531), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n866), .A2(G125), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U588 ( .A1(G137), .A2(n870), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G113), .A2(n865), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G160) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n580) );
  NAND2_X1 U593 ( .A1(n786), .A2(G51), .ZN(n539) );
  XOR2_X1 U594 ( .A(KEYINPUT75), .B(n539), .Z(n543) );
  INV_X1 U595 ( .A(G651), .ZN(n546) );
  NOR2_X1 U596 ( .A1(G543), .A2(n546), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n540), .Z(n782) );
  NAND2_X1 U598 ( .A1(n782), .A2(G63), .ZN(n541) );
  XNOR2_X1 U599 ( .A(KEYINPUT74), .B(n541), .ZN(n542) );
  AND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U601 ( .A(KEYINPUT6), .B(n544), .ZN(n551) );
  NOR2_X1 U602 ( .A1(G651), .A2(G543), .ZN(n779) );
  NAND2_X1 U603 ( .A1(n779), .A2(G89), .ZN(n545) );
  XNOR2_X1 U604 ( .A(n545), .B(KEYINPUT4), .ZN(n548) );
  NOR2_X1 U605 ( .A1(n580), .A2(n546), .ZN(n778) );
  NAND2_X1 U606 ( .A1(G76), .A2(n778), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n549), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT7), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT76), .ZN(G168) );
  NAND2_X1 U612 ( .A1(G52), .A2(n786), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G64), .A2(n782), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G77), .A2(n778), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G90), .A2(n779), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U619 ( .A1(n560), .A2(n559), .ZN(G171) );
  NAND2_X1 U620 ( .A1(G78), .A2(n778), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G91), .A2(n779), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U623 ( .A(KEYINPUT68), .B(n563), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G53), .A2(n786), .ZN(n564) );
  XNOR2_X1 U625 ( .A(KEYINPUT69), .B(n564), .ZN(n565) );
  NOR2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n782), .A2(G65), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U629 ( .A(KEYINPUT70), .B(n569), .ZN(G299) );
  XOR2_X1 U630 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U631 ( .A1(G75), .A2(n778), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G88), .A2(n779), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G50), .A2(n786), .ZN(n573) );
  NAND2_X1 U635 ( .A1(G62), .A2(n782), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U637 ( .A1(n575), .A2(n574), .ZN(G166) );
  XNOR2_X1 U638 ( .A(KEYINPUT85), .B(G166), .ZN(G303) );
  NAND2_X1 U639 ( .A1(G49), .A2(n786), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G74), .A2(G651), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n782), .A2(n578), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT80), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G87), .A2(n580), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U646 ( .A1(G86), .A2(n779), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G61), .A2(n782), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n778), .A2(G73), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT2), .B(n585), .Z(n586) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n786), .A2(G48), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(G305) );
  NAND2_X1 U654 ( .A1(G72), .A2(n778), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G85), .A2(n779), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G60), .A2(n782), .ZN(n592) );
  XNOR2_X1 U658 ( .A(KEYINPUT67), .B(n592), .ZN(n593) );
  NOR2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n786), .A2(G47), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(G290) );
  XOR2_X1 U662 ( .A(G2078), .B(KEYINPUT25), .Z(n993) );
  NOR2_X1 U663 ( .A1(G164), .A2(G1384), .ZN(n702) );
  NAND2_X1 U664 ( .A1(G160), .A2(G40), .ZN(n701) );
  INV_X1 U665 ( .A(n701), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n993), .A2(n661), .ZN(n599) );
  INV_X1 U667 ( .A(n661), .ZN(n613) );
  NOR2_X1 U668 ( .A1(n613), .A2(G1961), .ZN(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U670 ( .A(KEYINPUT93), .B(n600), .ZN(n651) );
  NAND2_X1 U671 ( .A1(n651), .A2(G171), .ZN(n645) );
  NAND2_X1 U672 ( .A1(n613), .A2(G2072), .ZN(n601) );
  XNOR2_X1 U673 ( .A(KEYINPUT27), .B(n601), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G1956), .A2(n661), .ZN(n602) );
  XOR2_X1 U675 ( .A(KEYINPUT94), .B(n602), .Z(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n639) );
  INV_X1 U677 ( .A(G299), .ZN(n638) );
  NAND2_X1 U678 ( .A1(n639), .A2(n638), .ZN(n637) );
  NAND2_X1 U679 ( .A1(G66), .A2(n782), .ZN(n611) );
  NAND2_X1 U680 ( .A1(G79), .A2(n778), .ZN(n606) );
  NAND2_X1 U681 ( .A1(G92), .A2(n779), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G54), .A2(n786), .ZN(n607) );
  XNOR2_X1 U684 ( .A(KEYINPUT73), .B(n607), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X2 U687 ( .A(n612), .B(KEYINPUT15), .ZN(n953) );
  INV_X1 U688 ( .A(n953), .ZN(n757) );
  NOR2_X1 U689 ( .A1(n613), .A2(G1348), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G2067), .A2(n661), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n632) );
  NAND2_X1 U692 ( .A1(n757), .A2(n632), .ZN(n631) );
  INV_X1 U693 ( .A(G1996), .ZN(n997) );
  NOR2_X1 U694 ( .A1(n661), .A2(n997), .ZN(n617) );
  INV_X1 U695 ( .A(KEYINPUT26), .ZN(n616) );
  XNOR2_X1 U696 ( .A(n617), .B(n616), .ZN(n629) );
  AND2_X1 U697 ( .A1(n661), .A2(G1341), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G56), .A2(n782), .ZN(n618) );
  XOR2_X1 U699 ( .A(KEYINPUT14), .B(n618), .Z(n624) );
  NAND2_X1 U700 ( .A1(n779), .A2(G81), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G68), .A2(n778), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U704 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n786), .A2(G43), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n954) );
  NOR2_X1 U708 ( .A1(n627), .A2(n954), .ZN(n628) );
  AND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U712 ( .A(KEYINPUT95), .B(n635), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n642) );
  NOR2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U715 ( .A(n640), .B(KEYINPUT28), .Z(n641) );
  AND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U717 ( .A(KEYINPUT29), .B(n643), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n657) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n695), .ZN(n673) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n661), .ZN(n670) );
  INV_X1 U721 ( .A(n670), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n646), .A2(G8), .ZN(n647) );
  OR2_X1 U723 ( .A1(n673), .A2(n647), .ZN(n648) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n648), .ZN(n649) );
  NOR2_X1 U725 ( .A1(G168), .A2(n649), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n650), .B(KEYINPUT96), .ZN(n653) );
  NOR2_X1 U727 ( .A1(n651), .A2(G171), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n674) );
  NAND2_X1 U731 ( .A1(n674), .A2(G286), .ZN(n659) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n695), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT98), .ZN(n663) );
  NOR2_X1 U734 ( .A1(n661), .A2(G2090), .ZN(n662) );
  NOR2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U736 ( .A(KEYINPUT99), .B(n664), .Z(n665) );
  NAND2_X1 U737 ( .A1(G303), .A2(n665), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n668), .A2(G8), .ZN(n669) );
  XNOR2_X1 U739 ( .A(n669), .B(KEYINPUT32), .ZN(n677) );
  NAND2_X1 U740 ( .A1(G8), .A2(n670), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT92), .B(n671), .Z(n672) );
  NOR2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n690) );
  NOR2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n947) );
  NOR2_X1 U746 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n947), .A2(n678), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n690), .A2(n679), .ZN(n681) );
  NAND2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n951) );
  INV_X1 U750 ( .A(n951), .ZN(n680) );
  AND2_X1 U751 ( .A1(n681), .A2(n517), .ZN(n682) );
  NAND2_X1 U752 ( .A1(n947), .A2(KEYINPUT33), .ZN(n683) );
  NOR2_X1 U753 ( .A1(n683), .A2(n695), .ZN(n685) );
  XOR2_X1 U754 ( .A(G1981), .B(G305), .Z(n939) );
  INV_X1 U755 ( .A(n939), .ZN(n684) );
  NOR2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U757 ( .A1(G2090), .A2(G303), .ZN(n688) );
  NAND2_X1 U758 ( .A1(G8), .A2(n688), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT100), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n692), .A2(n695), .ZN(n697) );
  NOR2_X1 U762 ( .A1(G1981), .A2(G305), .ZN(n693) );
  XOR2_X1 U763 ( .A(n693), .B(KEYINPUT24), .Z(n694) );
  OR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U766 ( .A(n700), .B(KEYINPUT101), .ZN(n737) );
  NOR2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n747) );
  XNOR2_X1 U768 ( .A(KEYINPUT37), .B(G2067), .ZN(n745) );
  NAND2_X1 U769 ( .A1(G104), .A2(n873), .ZN(n704) );
  NAND2_X1 U770 ( .A1(G140), .A2(n870), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n705), .ZN(n710) );
  NAND2_X1 U773 ( .A1(G116), .A2(n865), .ZN(n707) );
  NAND2_X1 U774 ( .A1(G128), .A2(n866), .ZN(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U776 ( .A(KEYINPUT35), .B(n708), .Z(n709) );
  NOR2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U778 ( .A(KEYINPUT36), .B(n711), .ZN(n886) );
  NOR2_X1 U779 ( .A1(n745), .A2(n886), .ZN(n918) );
  NAND2_X1 U780 ( .A1(n747), .A2(n918), .ZN(n743) );
  XOR2_X1 U781 ( .A(KEYINPUT89), .B(G1991), .Z(n1003) );
  INV_X1 U782 ( .A(n1003), .ZN(n722) );
  NAND2_X1 U783 ( .A1(G107), .A2(n865), .ZN(n713) );
  NAND2_X1 U784 ( .A1(G119), .A2(n866), .ZN(n712) );
  NAND2_X1 U785 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U786 ( .A(KEYINPUT86), .B(n714), .ZN(n717) );
  NAND2_X1 U787 ( .A1(G131), .A2(n870), .ZN(n715) );
  XNOR2_X1 U788 ( .A(KEYINPUT87), .B(n715), .ZN(n716) );
  NOR2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U790 ( .A1(n873), .A2(G95), .ZN(n718) );
  NAND2_X1 U791 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U792 ( .A(KEYINPUT88), .B(n720), .ZN(n885) );
  INV_X1 U793 ( .A(n885), .ZN(n721) );
  NOR2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U795 ( .A(n723), .B(KEYINPUT90), .ZN(n732) );
  NAND2_X1 U796 ( .A1(G117), .A2(n865), .ZN(n725) );
  NAND2_X1 U797 ( .A1(G129), .A2(n866), .ZN(n724) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n873), .A2(G105), .ZN(n726) );
  XOR2_X1 U800 ( .A(KEYINPUT38), .B(n726), .Z(n727) );
  NOR2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n730) );
  NAND2_X1 U802 ( .A1(n870), .A2(G141), .ZN(n729) );
  NAND2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n881) );
  AND2_X1 U804 ( .A1(G1996), .A2(n881), .ZN(n731) );
  NOR2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n924) );
  INV_X1 U806 ( .A(n747), .ZN(n733) );
  NOR2_X1 U807 ( .A1(n924), .A2(n733), .ZN(n740) );
  INV_X1 U808 ( .A(n740), .ZN(n734) );
  NAND2_X1 U809 ( .A1(n743), .A2(n734), .ZN(n735) );
  XOR2_X1 U810 ( .A(KEYINPUT91), .B(n735), .Z(n736) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n944) );
  NAND2_X1 U812 ( .A1(n737), .A2(n519), .ZN(n750) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n881), .ZN(n913) );
  NOR2_X1 U814 ( .A1(n1003), .A2(n885), .ZN(n922) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n738) );
  NOR2_X1 U816 ( .A1(n922), .A2(n738), .ZN(n739) );
  NOR2_X1 U817 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U818 ( .A1(n913), .A2(n741), .ZN(n742) );
  XNOR2_X1 U819 ( .A(KEYINPUT39), .B(n742), .ZN(n744) );
  NAND2_X1 U820 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n745), .A2(n886), .ZN(n926) );
  NAND2_X1 U822 ( .A1(n746), .A2(n926), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U826 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U827 ( .A(G132), .ZN(G219) );
  INV_X1 U828 ( .A(G82), .ZN(G220) );
  INV_X1 U829 ( .A(G57), .ZN(G237) );
  XOR2_X1 U830 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n753) );
  NAND2_X1 U831 ( .A1(G7), .A2(G661), .ZN(n752) );
  XNOR2_X1 U832 ( .A(n753), .B(n752), .ZN(G223) );
  XOR2_X1 U833 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n755) );
  INV_X1 U834 ( .A(G223), .ZN(n818) );
  NAND2_X1 U835 ( .A1(G567), .A2(n818), .ZN(n754) );
  XNOR2_X1 U836 ( .A(n755), .B(n754), .ZN(G234) );
  INV_X1 U837 ( .A(n954), .ZN(n756) );
  NAND2_X1 U838 ( .A1(n756), .A2(G860), .ZN(G153) );
  INV_X1 U839 ( .A(G171), .ZN(G301) );
  NAND2_X1 U840 ( .A1(G868), .A2(G301), .ZN(n759) );
  INV_X1 U841 ( .A(G868), .ZN(n800) );
  NAND2_X1 U842 ( .A1(n757), .A2(n800), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n759), .A2(n758), .ZN(G284) );
  NAND2_X1 U844 ( .A1(G868), .A2(G286), .ZN(n761) );
  NAND2_X1 U845 ( .A1(G299), .A2(n800), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n761), .A2(n760), .ZN(G297) );
  INV_X1 U847 ( .A(G559), .ZN(n762) );
  NOR2_X1 U848 ( .A1(G860), .A2(n762), .ZN(n763) );
  XNOR2_X1 U849 ( .A(KEYINPUT77), .B(n763), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n764), .A2(n953), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n765), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U852 ( .A1(G868), .A2(n954), .ZN(n768) );
  NAND2_X1 U853 ( .A1(G868), .A2(n953), .ZN(n766) );
  NOR2_X1 U854 ( .A1(G559), .A2(n766), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(G282) );
  NAND2_X1 U856 ( .A1(G99), .A2(n873), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G111), .A2(n865), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n866), .A2(G123), .ZN(n771) );
  XOR2_X1 U860 ( .A(KEYINPUT18), .B(n771), .Z(n772) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n870), .A2(G135), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n915) );
  XNOR2_X1 U864 ( .A(G2096), .B(n915), .ZN(n776) );
  NOR2_X1 U865 ( .A1(G2100), .A2(n776), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT78), .B(n777), .Z(G156) );
  NAND2_X1 U867 ( .A1(G80), .A2(n778), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G93), .A2(n779), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G67), .A2(n782), .ZN(n783) );
  XNOR2_X1 U871 ( .A(KEYINPUT79), .B(n783), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U873 ( .A1(n786), .A2(G55), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n799) );
  NAND2_X1 U875 ( .A1(G559), .A2(n953), .ZN(n789) );
  XNOR2_X1 U876 ( .A(n789), .B(n954), .ZN(n797) );
  NOR2_X1 U877 ( .A1(G860), .A2(n797), .ZN(n790) );
  XOR2_X1 U878 ( .A(n799), .B(n790), .Z(G145) );
  XOR2_X1 U879 ( .A(G290), .B(G305), .Z(n791) );
  XNOR2_X1 U880 ( .A(G288), .B(n791), .ZN(n794) );
  XOR2_X1 U881 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n792) );
  XNOR2_X1 U882 ( .A(n799), .B(n792), .ZN(n793) );
  XOR2_X1 U883 ( .A(n794), .B(n793), .Z(n796) );
  XNOR2_X1 U884 ( .A(G299), .B(G166), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n796), .B(n795), .ZN(n891) );
  XNOR2_X1 U886 ( .A(n797), .B(n891), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n798), .A2(G868), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U890 ( .A(KEYINPUT82), .B(n803), .ZN(G295) );
  NAND2_X1 U891 ( .A1(G2078), .A2(G2084), .ZN(n804) );
  XOR2_X1 U892 ( .A(KEYINPUT20), .B(n804), .Z(n805) );
  NAND2_X1 U893 ( .A1(G2090), .A2(n805), .ZN(n806) );
  XNOR2_X1 U894 ( .A(KEYINPUT21), .B(n806), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n807), .A2(G2072), .ZN(G158) );
  XOR2_X1 U896 ( .A(KEYINPUT83), .B(G44), .Z(n808) );
  XNOR2_X1 U897 ( .A(KEYINPUT3), .B(n808), .ZN(G218) );
  NAND2_X1 U898 ( .A1(G108), .A2(G120), .ZN(n809) );
  NOR2_X1 U899 ( .A1(G237), .A2(n809), .ZN(n810) );
  NAND2_X1 U900 ( .A1(G69), .A2(n810), .ZN(n823) );
  NAND2_X1 U901 ( .A1(n823), .A2(G567), .ZN(n816) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n811) );
  XNOR2_X1 U903 ( .A(KEYINPUT22), .B(n811), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n812), .A2(G96), .ZN(n813) );
  NOR2_X1 U905 ( .A1(G218), .A2(n813), .ZN(n814) );
  XOR2_X1 U906 ( .A(KEYINPUT84), .B(n814), .Z(n824) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n824), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n825) );
  NAND2_X1 U909 ( .A1(G661), .A2(G483), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n825), .A2(n817), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n822), .A2(G36), .ZN(G176) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U914 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n820) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n820), .Z(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(G188) );
  XOR2_X1 U918 ( .A(G120), .B(KEYINPUT104), .Z(G236) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(G325) );
  XNOR2_X1 U920 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U922 ( .A(G108), .ZN(G238) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(n825), .ZN(G319) );
  XNOR2_X1 U925 ( .A(G1961), .B(G2474), .ZN(n835) );
  XOR2_X1 U926 ( .A(G1976), .B(G1971), .Z(n827) );
  XNOR2_X1 U927 ( .A(G1986), .B(G1966), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U929 ( .A(G1981), .B(G1956), .Z(n829) );
  XNOR2_X1 U930 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U931 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U932 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U933 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(G229) );
  XOR2_X1 U936 ( .A(KEYINPUT107), .B(G2678), .Z(n837) );
  XNOR2_X1 U937 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2090), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U942 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2096), .B(G2100), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U945 ( .A(G2078), .B(G2084), .Z(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(G227) );
  NAND2_X1 U947 ( .A1(G100), .A2(n873), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G112), .A2(n865), .ZN(n846) );
  NAND2_X1 U949 ( .A1(n847), .A2(n846), .ZN(n853) );
  NAND2_X1 U950 ( .A1(n866), .A2(G124), .ZN(n848) );
  XOR2_X1 U951 ( .A(KEYINPUT44), .B(n848), .Z(n849) );
  XNOR2_X1 U952 ( .A(n849), .B(KEYINPUT109), .ZN(n851) );
  NAND2_X1 U953 ( .A1(G136), .A2(n870), .ZN(n850) );
  NAND2_X1 U954 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U955 ( .A1(n853), .A2(n852), .ZN(G162) );
  NAND2_X1 U956 ( .A1(G130), .A2(n866), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n854), .B(KEYINPUT110), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G118), .A2(n865), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n857), .B(KEYINPUT111), .ZN(n863) );
  XNOR2_X1 U961 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G106), .A2(n873), .ZN(n859) );
  NAND2_X1 U963 ( .A1(G142), .A2(n870), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U965 ( .A(n861), .B(n860), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n889) );
  XOR2_X1 U967 ( .A(G160), .B(G162), .Z(n864) );
  XNOR2_X1 U968 ( .A(n915), .B(n864), .ZN(n880) );
  XOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n878) );
  NAND2_X1 U970 ( .A1(G115), .A2(n865), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G127), .A2(n866), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n869), .B(KEYINPUT47), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G139), .A2(n870), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G103), .A2(n873), .ZN(n874) );
  XNOR2_X1 U977 ( .A(KEYINPUT113), .B(n874), .ZN(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n928) );
  XNOR2_X1 U979 ( .A(n928), .B(KEYINPUT114), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(n880), .B(n879), .Z(n883) );
  XOR2_X1 U982 ( .A(G164), .B(n881), .Z(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U987 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U988 ( .A(n954), .B(n891), .ZN(n893) );
  XNOR2_X1 U989 ( .A(G171), .B(n953), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U991 ( .A(n894), .B(G286), .Z(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(G397) );
  XOR2_X1 U993 ( .A(KEYINPUT102), .B(G2446), .Z(n897) );
  XNOR2_X1 U994 ( .A(G2443), .B(G2454), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(n898), .B(G2451), .Z(n900) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U999 ( .A(G2435), .B(G2427), .Z(n902) );
  XNOR2_X1 U1000 ( .A(G2430), .B(G2438), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1003 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  INV_X1 U1012 ( .A(n911), .ZN(G401) );
  XNOR2_X1 U1013 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1023) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n912) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1016 ( .A(KEYINPUT51), .B(n914), .Z(n920) );
  XNOR2_X1 U1017 ( .A(G160), .B(G2084), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT115), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1025 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT50), .B(n931), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n934), .ZN(n936) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n937), .A2(G29), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT116), .B(n938), .ZN(n1021) );
  XNOR2_X1 U1035 ( .A(G16), .B(KEYINPUT56), .ZN(n964) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G168), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(n941), .B(KEYINPUT57), .ZN(n962) );
  XNOR2_X1 U1039 ( .A(G1956), .B(G299), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(n942), .B(KEYINPUT121), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G1961), .B(G301), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n960) );
  XNOR2_X1 U1044 ( .A(G303), .B(G1971), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(n947), .B(KEYINPUT122), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n952), .B(KEYINPUT123), .ZN(n958) );
  XOR2_X1 U1049 ( .A(G1348), .B(n953), .Z(n956) );
  XNOR2_X1 U1050 ( .A(n954), .B(G1341), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n991) );
  INV_X1 U1056 ( .A(G16), .ZN(n989) );
  XNOR2_X1 U1057 ( .A(G1348), .B(KEYINPUT59), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n965), .B(G4), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(G1341), .B(G19), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1981), .B(G6), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT124), .B(G1956), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(G20), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT60), .B(n973), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G21), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G1961), .B(G5), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n985) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G23), .B(G1976), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(G1986), .B(KEYINPUT125), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(G24), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT58), .B(n983), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(KEYINPUT61), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT126), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n1019) );
  XNOR2_X1 U1083 ( .A(KEYINPUT117), .B(G2067), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(n992), .B(G26), .ZN(n1002) );
  XNOR2_X1 U1085 ( .A(n993), .B(G27), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(G2072), .B(G33), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(G28), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(G32), .B(n997), .Z(n998) );
  XNOR2_X1 U1090 ( .A(KEYINPUT118), .B(n998), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G25), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT53), .B(n1006), .Z(n1010) );
  XNOR2_X1 U1096 ( .A(KEYINPUT54), .B(G34), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT119), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(G2084), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(G35), .B(G2090), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1013), .B(KEYINPUT55), .ZN(n1015) );
  INV_X1 U1103 ( .A(G29), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(G11), .A2(n1016), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(KEYINPUT120), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(n1023), .B(n1022), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

