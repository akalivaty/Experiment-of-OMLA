//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1323, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n204), .A2(G50), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT66), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT67), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n215), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  XNOR2_X1  g0044(.A(KEYINPUT3), .B(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(G222), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(G223), .A3(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G77), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n247), .A2(new_n248), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  INV_X1    g0058(.A(G45), .ZN(new_n259));
  AOI21_X1  g0059(.A(G1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n262), .A3(G274), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT68), .B(G226), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G179), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n218), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n210), .B1(new_n201), .B2(new_n203), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n251), .A2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G150), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI22_X1  g0082(.A1(new_n277), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n275), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n275), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n209), .B2(G20), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n287), .A2(new_n289), .B1(new_n288), .B2(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n273), .B(new_n291), .C1(G169), .C2(new_n271), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n245), .A2(G238), .A3(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n245), .A2(G232), .A3(new_n246), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n253), .A2(G107), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n256), .ZN(new_n297));
  INV_X1    g0097(.A(G244), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n263), .B1(new_n298), .B2(new_n266), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n299), .B1(new_n296), .B2(new_n256), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n272), .ZN(new_n305));
  INV_X1    g0105(.A(new_n275), .ZN(new_n306));
  INV_X1    g0106(.A(G87), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT15), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT15), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT69), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(KEYINPUT70), .A3(new_n278), .A4(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n277), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(new_n278), .A3(new_n314), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n306), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n209), .B2(G20), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n287), .A2(new_n324), .B1(new_n323), .B2(new_n286), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n303), .B(new_n305), .C1(new_n322), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT71), .B(G200), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n301), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n321), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n315), .A2(new_n317), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n275), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n304), .A2(G190), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n332), .A3(new_n325), .A4(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n292), .A2(new_n327), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n270), .A2(new_n328), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT9), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n291), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n257), .A2(new_n269), .A3(G190), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n284), .A2(KEYINPUT9), .A3(new_n290), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n336), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT10), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n341), .A2(KEYINPUT10), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n335), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G226), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n246), .ZN(new_n346));
  INV_X1    g0146(.A(G232), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G1698), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n250), .A2(new_n346), .A3(new_n252), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n256), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n267), .A2(G238), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n263), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G238), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n263), .B1(new_n356), .B2(new_n266), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n262), .B1(new_n349), .B2(new_n350), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT13), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n359), .A3(G190), .ZN(new_n360));
  INV_X1    g0160(.A(G68), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n281), .A2(G50), .B1(G20), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n279), .B2(new_n323), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n275), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT11), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n368));
  OR3_X1    g0168(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n361), .B1(new_n209), .B2(G20), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n368), .A2(new_n369), .B1(new_n287), .B2(new_n370), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n366), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n355), .B2(new_n359), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT72), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT72), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n360), .A4(new_n372), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n372), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n355), .A2(new_n359), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT14), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(G169), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n355), .A2(new_n359), .A3(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n382), .B2(G169), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n381), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n344), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n277), .B1(new_n209), .B2(G20), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(new_n287), .B1(new_n286), .B2(new_n277), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(G58), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(new_n361), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n203), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n281), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n249), .A2(KEYINPUT73), .A3(G33), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n252), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT73), .B1(new_n249), .B2(G33), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n399), .B(new_n210), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G68), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT73), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(new_n400), .A3(new_n252), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n399), .B1(new_n407), .B2(new_n210), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT16), .B(new_n398), .C1(new_n404), .C2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n409), .A2(new_n275), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n399), .B1(new_n245), .B2(G20), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n361), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n398), .B1(new_n414), .B2(KEYINPUT74), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT74), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n416), .B(new_n361), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n392), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n262), .A2(G232), .A3(new_n265), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n263), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n345), .A2(G1698), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G223), .B2(G1698), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n407), .A2(new_n423), .B1(new_n251), .B2(new_n307), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n421), .B1(new_n424), .B2(new_n256), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G179), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n302), .B2(new_n425), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT18), .B1(new_n419), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT7), .B1(new_n253), .B2(new_n210), .ZN(new_n430));
  AOI211_X1 g0230(.A(new_n399), .B(G20), .C1(new_n250), .C2(new_n252), .ZN(new_n431));
  OAI21_X1  g0231(.A(G68), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n397), .B1(new_n432), .B2(new_n416), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n414), .A2(KEYINPUT74), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT16), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n409), .A2(new_n275), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n391), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT18), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n427), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n440), .B(new_n421), .C1(new_n256), .C2(new_n424), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n424), .A2(new_n256), .ZN(new_n442));
  INV_X1    g0242(.A(new_n421), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n374), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n391), .B(new_n445), .C1(new_n435), .C2(new_n436), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT17), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n410), .A2(new_n418), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n449), .A2(KEYINPUT17), .A3(new_n391), .A4(new_n445), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n429), .A2(new_n439), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n389), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n274), .A2(new_n218), .B1(G20), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n210), .C1(G33), .C2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT20), .B1(new_n455), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n285), .A2(new_n454), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n209), .A2(G33), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n285), .A2(new_n464), .A3(new_n218), .A4(new_n274), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(G116), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT78), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n455), .A2(new_n458), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  INV_X1    g0273(.A(new_n465), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n462), .B1(new_n474), .B2(new_n454), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n209), .A2(G45), .ZN(new_n479));
  OR2_X1    g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(new_n256), .ZN(new_n483));
  INV_X1    g0283(.A(G274), .ZN(new_n484));
  INV_X1    g0284(.A(new_n218), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n261), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n483), .A2(G270), .B1(new_n486), .B2(new_n482), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n253), .A2(G303), .ZN(new_n488));
  INV_X1    g0288(.A(G264), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G1698), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(G257), .B2(G1698), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n407), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n256), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n400), .A2(new_n252), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G257), .A2(G1698), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n489), .B2(G1698), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n406), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n262), .B1(new_n499), .B2(new_n488), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT5), .B(G41), .ZN(new_n501));
  INV_X1    g0301(.A(new_n479), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(G270), .A3(new_n262), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n482), .A2(new_n486), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G190), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n478), .A2(new_n495), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n302), .B1(new_n487), .B2(new_n493), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT78), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n473), .B1(new_n472), .B2(new_n475), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n494), .A2(new_n272), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n477), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n477), .A2(KEYINPUT21), .A3(new_n510), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n509), .A2(new_n515), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G107), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT25), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n285), .B2(G107), .ZN(new_n523));
  AOI22_X1  g0323(.A1(G107), .A2(new_n474), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n210), .A2(G87), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n253), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G20), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n210), .B2(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n520), .A2(KEYINPUT23), .A3(G20), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n406), .A2(new_n400), .A3(new_n210), .A4(new_n252), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n525), .A2(new_n307), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT24), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n496), .A2(new_n210), .A3(new_n406), .A4(new_n536), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(new_n527), .A4(new_n533), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT79), .B1(new_n543), .B2(new_n275), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT79), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n545), .B(new_n306), .C1(new_n539), .C2(new_n542), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n524), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g0347(.A1(G250), .A2(G1698), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G257), .B2(new_n246), .ZN(new_n549));
  INV_X1    g0349(.A(G294), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n407), .A2(new_n549), .B1(new_n251), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(new_n256), .B1(new_n483), .B2(G264), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n505), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G179), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n302), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n374), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n256), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n483), .A2(G264), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n558), .A2(new_n440), .A3(new_n505), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT80), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT80), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n552), .A2(new_n562), .A3(new_n440), .A4(new_n505), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n564), .B(new_n524), .C1(new_n544), .C2(new_n546), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n503), .A2(G257), .A3(new_n262), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n505), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT4), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n298), .A2(G1698), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n407), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n569), .A2(new_n298), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n245), .A2(new_n246), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n250), .A2(new_n252), .A3(G250), .A4(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n456), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n568), .B1(new_n576), .B2(new_n256), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n272), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n406), .A2(new_n400), .A3(new_n252), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT4), .B1(new_n579), .B2(new_n570), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n456), .A3(new_n575), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n256), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n568), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n302), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n520), .A2(KEYINPUT6), .A3(G97), .ZN(new_n586));
  XNOR2_X1  g0386(.A(G97), .B(G107), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT6), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n589), .A2(new_n210), .B1(new_n323), .B2(new_n282), .ZN(new_n590));
  OAI21_X1  g0390(.A(G107), .B1(new_n430), .B2(new_n431), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(KEYINPUT75), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n520), .B1(new_n412), .B2(new_n413), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT75), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n306), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT76), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n285), .B2(G97), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n285), .A2(new_n597), .A3(G97), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(new_n600), .B1(new_n457), .B2(new_n465), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n578), .B(new_n585), .C1(new_n596), .C2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n210), .B1(new_n350), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G97), .A2(G107), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n307), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(new_n606), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n361), .B2(new_n535), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n275), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n313), .A2(new_n314), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n286), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n465), .A2(new_n307), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT77), .ZN(new_n616));
  NOR2_X1   g0416(.A1(G238), .A2(G1698), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n298), .B2(G1698), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n496), .A2(new_n406), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(new_n528), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n298), .A2(G1698), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G238), .B2(G1698), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n616), .B(new_n528), .C1(new_n407), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n256), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n486), .A2(new_n502), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n479), .A2(G250), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n262), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n328), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n528), .B1(new_n407), .B2(new_n622), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT77), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n262), .B1(new_n632), .B2(new_n623), .ZN(new_n633));
  INV_X1    g0433(.A(new_n629), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n633), .A2(G190), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n615), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n457), .A2(new_n520), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n588), .B1(new_n637), .B2(new_n605), .ZN(new_n638));
  INV_X1    g0438(.A(new_n586), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n594), .B2(new_n593), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n591), .A2(KEYINPUT75), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n275), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n601), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n582), .A2(new_n440), .A3(new_n583), .ZN(new_n646));
  AOI21_X1  g0446(.A(G200), .B1(new_n582), .B2(new_n583), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n302), .B1(new_n633), .B2(new_n634), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n609), .A2(new_n275), .B1(new_n286), .B2(new_n611), .ZN(new_n650));
  INV_X1    g0450(.A(new_n611), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n474), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n625), .A2(new_n629), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n649), .B(new_n653), .C1(new_n654), .C2(G179), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n602), .A2(new_n636), .A3(new_n648), .A4(new_n655), .ZN(new_n656));
  NOR4_X1   g0456(.A1(new_n453), .A2(new_n519), .A3(new_n566), .A4(new_n656), .ZN(G372));
  INV_X1    g0457(.A(new_n292), .ZN(new_n658));
  INV_X1    g0458(.A(new_n388), .ZN(new_n659));
  INV_X1    g0459(.A(new_n327), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n380), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n448), .A2(new_n450), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n429), .B(new_n439), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT82), .ZN(new_n664));
  INV_X1    g0464(.A(new_n342), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n341), .A2(KEYINPUT10), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n343), .A2(KEYINPUT82), .A3(new_n342), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n658), .B1(new_n663), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n328), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n633), .B2(new_n634), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n654), .B2(G190), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT81), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n613), .B2(new_n614), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n650), .B(KEYINPUT81), .C1(new_n307), .C2(new_n465), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n585), .A2(new_n578), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n591), .A2(KEYINPUT75), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n595), .A3(new_n641), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n601), .B1(new_n681), .B2(new_n275), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n678), .A2(new_n683), .A3(new_n655), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n636), .A2(new_n655), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(KEYINPUT26), .A3(new_n683), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n678), .A2(new_n602), .A3(new_n648), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n556), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n692), .A3(new_n565), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n693), .A3(new_n655), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n670), .B1(new_n453), .B2(new_n695), .ZN(G369));
  OR2_X1    g0496(.A1(new_n519), .A2(KEYINPUT84), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT83), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n698), .B(KEYINPUT83), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(new_n704), .A3(G213), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n478), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n519), .B2(KEYINPUT84), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n697), .A2(new_n710), .B1(new_n691), .B2(new_n709), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n547), .A2(new_n707), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n566), .A2(new_n712), .B1(new_n556), .B2(new_n708), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(G330), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n547), .A2(new_n555), .A3(new_n708), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n556), .A2(new_n565), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n708), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n714), .A2(new_n715), .A3(new_n720), .ZN(G399));
  NOR2_X1   g0521(.A1(new_n606), .A2(G116), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT85), .ZN(new_n723));
  INV_X1    g0523(.A(new_n213), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G41), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n723), .A2(new_n725), .A3(new_n209), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n217), .B2(new_n725), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  NOR2_X1   g0528(.A1(new_n633), .A2(new_n634), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n272), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n649), .A2(new_n653), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n730), .A2(new_n731), .B1(new_n673), .B2(new_n677), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT26), .B1(new_n732), .B2(new_n683), .ZN(new_n733));
  AND4_X1   g0533(.A1(KEYINPUT26), .A2(new_n683), .A3(new_n636), .A4(new_n655), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n717), .B1(new_n547), .B2(new_n555), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n565), .A2(new_n678), .A3(new_n602), .A4(new_n648), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n655), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n708), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT88), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n694), .A2(KEYINPUT88), .A3(new_n708), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n684), .A2(KEYINPUT26), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n687), .A2(new_n685), .A3(new_n683), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(KEYINPUT29), .B(new_n708), .C1(new_n738), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT87), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT30), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n577), .A2(new_n507), .A3(G179), .A4(new_n552), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(new_n654), .ZN(new_n753));
  AOI21_X1  g0553(.A(G179), .B1(new_n487), .B2(new_n493), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n584), .A2(new_n754), .A3(new_n553), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT86), .B1(new_n755), .B2(new_n729), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n558), .A2(new_n505), .A3(new_n559), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n272), .B1(new_n500), .B2(new_n506), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT86), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n759), .A2(new_n760), .A3(new_n654), .A4(new_n584), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n582), .A2(new_n552), .A3(new_n583), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(new_n729), .A3(new_n516), .A4(KEYINPUT30), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n753), .A2(new_n756), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n707), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n753), .B(new_n763), .C1(new_n729), .C2(new_n755), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n708), .A2(new_n766), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n519), .ZN(new_n770));
  AND4_X1   g0570(.A1(new_n636), .A2(new_n602), .A3(new_n648), .A4(new_n655), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n716), .A2(new_n770), .A3(new_n771), .A4(new_n708), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n750), .B1(new_n773), .B2(G330), .ZN(new_n774));
  INV_X1    g0574(.A(G330), .ZN(new_n775));
  AOI211_X1 g0575(.A(KEYINPUT87), .B(new_n775), .C1(new_n769), .C2(new_n772), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n749), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT89), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n749), .A2(KEYINPUT89), .A3(new_n777), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n728), .B1(new_n782), .B2(G1), .ZN(G364));
  NAND2_X1  g0583(.A1(new_n711), .A2(G330), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n210), .A2(G13), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n209), .B1(new_n785), .B2(G45), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n725), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n711), .A2(G330), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OR3_X1    g0592(.A1(KEYINPUT91), .A2(G13), .A3(G33), .ZN(new_n793));
  OAI21_X1  g0593(.A(KEYINPUT91), .B1(G13), .B2(G33), .ZN(new_n794));
  AOI21_X1  g0594(.A(G20), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT97), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n711), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n724), .A2(new_n253), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n454), .B2(new_n724), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT90), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n217), .A2(new_n259), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n724), .A2(new_n579), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n243), .C2(new_n259), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(KEYINPUT90), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n801), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n218), .B1(G20), .B2(new_n302), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n795), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n788), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(G20), .A2(G179), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT92), .Z(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G190), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n374), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n812), .A2(G190), .A3(new_n374), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n288), .B1(new_n393), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G190), .A2(G200), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n374), .A2(G190), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n820), .A2(new_n323), .B1(new_n361), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n440), .A2(G179), .A3(G200), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n210), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n457), .ZN(new_n826));
  NOR4_X1   g0626(.A1(new_n210), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G159), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT32), .ZN(new_n829));
  OR3_X1    g0629(.A1(new_n823), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n328), .A2(new_n272), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT93), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n210), .B1(new_n831), .B2(KEYINPUT93), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n440), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n245), .B1(new_n836), .B2(new_n307), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n817), .B(new_n830), .C1(KEYINPUT94), .C2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n832), .A2(new_n440), .A3(new_n833), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n839), .A2(KEYINPUT95), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(KEYINPUT95), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n838), .B1(KEYINPUT94), .B2(new_n837), .C1(new_n520), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n245), .B1(new_n835), .B2(G303), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT96), .ZN(new_n845));
  INV_X1    g0645(.A(new_n825), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n846), .A2(G294), .B1(G329), .B2(new_n827), .ZN(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n820), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n822), .ZN(new_n850));
  XNOR2_X1  g0650(.A(KEYINPUT33), .B(G317), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n816), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G326), .A2(new_n814), .B1(new_n853), .B2(G322), .ZN(new_n854));
  INV_X1    g0654(.A(G283), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n852), .B(new_n854), .C1(new_n842), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n843), .B1(new_n845), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n810), .B1(new_n857), .B2(new_n807), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n792), .B1(new_n797), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G396));
  OAI21_X1  g0660(.A(new_n707), .B1(new_n322), .B2(new_n326), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n327), .A2(new_n334), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT99), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n327), .A2(new_n334), .A3(new_n861), .A4(KEYINPUT99), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT100), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n660), .A2(new_n867), .A3(new_n707), .ZN(new_n868));
  OAI21_X1  g0668(.A(KEYINPUT100), .B1(new_n327), .B2(new_n708), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n741), .A2(new_n743), .A3(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n708), .B(new_n871), .C1(new_n735), .C2(new_n738), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n773), .A2(G330), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT87), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n773), .A2(new_n750), .A3(G330), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT101), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(new_n873), .A3(KEYINPUT101), .A4(new_n874), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n789), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT102), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n873), .A2(new_n874), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n777), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT101), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n884), .B2(new_n777), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT102), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n789), .A4(new_n881), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n842), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(G87), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n850), .A2(G283), .ZN(new_n893));
  AOI22_X1  g0693(.A1(G303), .A2(new_n814), .B1(new_n853), .B2(G294), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n819), .A2(G116), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n245), .B(new_n826), .C1(G311), .C2(new_n827), .ZN(new_n896));
  AND4_X1   g0696(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n892), .B(new_n897), .C1(new_n520), .C2(new_n836), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n891), .A2(G68), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n825), .A2(new_n393), .ZN(new_n900));
  INV_X1    g0700(.A(new_n827), .ZN(new_n901));
  INV_X1    g0701(.A(G132), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n579), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n900), .B(new_n903), .C1(new_n835), .C2(G50), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT98), .Z(new_n906));
  AOI22_X1  g0706(.A1(G150), .A2(new_n850), .B1(new_n819), .B2(G159), .ZN(new_n907));
  INV_X1    g0707(.A(G143), .ZN(new_n908));
  INV_X1    g0708(.A(G137), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n907), .B1(new_n908), .B2(new_n816), .C1(new_n909), .C2(new_n815), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT34), .Z(new_n911));
  OAI21_X1  g0711(.A(new_n898), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n807), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n793), .A2(new_n794), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n872), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n807), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n789), .B1(new_n323), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n890), .A2(new_n918), .ZN(G384));
  OR2_X1    g0719(.A1(new_n640), .A2(KEYINPUT35), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n640), .A2(KEYINPUT35), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n920), .A2(G116), .A3(new_n219), .A4(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT36), .Z(new_n923));
  OAI211_X1 g0723(.A(new_n217), .B(G77), .C1(new_n393), .C2(new_n361), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n201), .A2(G68), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n209), .B(G13), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n744), .A2(new_n452), .A3(new_n748), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n670), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n381), .A2(new_n707), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n380), .A2(new_n388), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n380), .B2(new_n388), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n327), .A2(new_n707), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n874), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT7), .B1(new_n579), .B2(G20), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(G68), .A3(new_n403), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT16), .B1(new_n938), .B2(new_n398), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n391), .B1(new_n436), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n705), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n451), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n427), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n942), .A3(new_n446), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT37), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n437), .A2(new_n427), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n437), .A2(new_n941), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT37), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n446), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n944), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT38), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n944), .A2(new_n952), .A3(KEYINPUT38), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n936), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT39), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n944), .A2(new_n952), .A3(KEYINPUT38), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n446), .B1(new_n419), .B2(new_n428), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n419), .A2(new_n705), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT37), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n951), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n429), .A2(new_n439), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n962), .B1(new_n965), .B2(new_n662), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT38), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n959), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n955), .A2(KEYINPUT39), .A3(new_n956), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n659), .A2(new_n708), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n965), .A2(new_n705), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n958), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n929), .B(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n960), .A2(new_n967), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n765), .A2(new_n766), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n772), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n380), .A2(new_n388), .ZN(new_n980));
  INV_X1    g0780(.A(new_n930), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n380), .A2(new_n388), .A3(new_n930), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(new_n866), .B2(new_n870), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT40), .B1(new_n976), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n864), .A2(new_n865), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n868), .A2(new_n869), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n987), .A2(new_n988), .B1(new_n931), .B2(new_n932), .ZN(new_n989));
  INV_X1    g0789(.A(new_n978), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT31), .B1(new_n764), .B2(new_n707), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n989), .B1(new_n772), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT40), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n957), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n986), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n452), .A3(new_n979), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n979), .B(new_n984), .C1(new_n960), .C2(new_n967), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n977), .A2(new_n978), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n566), .A2(new_n656), .A3(new_n519), .A4(new_n707), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n984), .B(new_n994), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(KEYINPUT40), .A2(new_n998), .B1(new_n1002), .B2(new_n957), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n979), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n453), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n997), .A2(new_n1005), .A3(G330), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n975), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n209), .B2(new_n785), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n975), .A2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n927), .B1(new_n1008), .B2(new_n1009), .ZN(G367));
  INV_X1    g0810(.A(KEYINPUT105), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n602), .B(new_n648), .C1(new_n682), .C2(new_n708), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n602), .B1(new_n1012), .B2(new_n556), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n708), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n683), .A2(new_n707), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT104), .B1(new_n720), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT104), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n716), .A3(new_n719), .A4(new_n1019), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n1018), .A2(KEYINPUT42), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT42), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1014), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n675), .A2(new_n676), .A3(new_n707), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT103), .B1(new_n655), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n732), .B2(new_n1024), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n655), .A2(new_n1024), .A3(KEYINPUT103), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(KEYINPUT43), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1011), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT42), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1018), .A2(KEYINPUT42), .A3(new_n1020), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1036), .A2(KEYINPUT105), .A3(new_n1029), .A4(new_n1014), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1028), .A2(KEYINPUT43), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1023), .A2(new_n1030), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1031), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT106), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n714), .A2(new_n1017), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1042), .A2(new_n1041), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1042), .A2(new_n1041), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1044), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n720), .B1(new_n713), .B2(new_n719), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n784), .B(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n720), .A2(new_n715), .A3(new_n1016), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n1052));
  AND2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n715), .B1(new_n566), .B2(new_n718), .ZN(new_n1055));
  AND3_X1   g0855(.A1(new_n1055), .A2(KEYINPUT44), .A3(new_n1017), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT44), .B1(new_n1055), .B2(new_n1017), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1053), .A2(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT109), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n1059), .A3(new_n714), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1051), .B(new_n1052), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n714), .A2(new_n1059), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n711), .A2(KEYINPUT109), .A3(G330), .A4(new_n713), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n780), .A2(new_n781), .B1(new_n1050), .B2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n725), .B(new_n1068), .Z(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n786), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1047), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT46), .B1(new_n835), .B2(G116), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n820), .A2(new_n855), .B1(new_n520), .B2(new_n825), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G294), .B2(new_n850), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n835), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G311), .A2(new_n814), .B1(new_n853), .B2(G303), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n891), .A2(G97), .ZN(new_n1079));
  INV_X1    g0879(.A(G317), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n407), .C1(new_n1080), .C2(new_n901), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT110), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1073), .B(new_n1078), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n846), .A2(G68), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n253), .B1(new_n827), .B2(G137), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n820), .C2(new_n201), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n815), .A2(new_n908), .B1(new_n280), .B2(new_n816), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G159), .C2(new_n850), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n891), .A2(G77), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n393), .C2(new_n836), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT47), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n807), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n809), .B1(new_n651), .B2(new_n724), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n803), .A2(new_n236), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n789), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1028), .B2(new_n796), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1072), .A2(new_n1100), .ZN(G387));
  AOI21_X1  g0901(.A(new_n1049), .B1(new_n780), .B2(new_n781), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n780), .A2(new_n781), .A3(new_n1049), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n725), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n713), .A2(new_n796), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n723), .A2(new_n798), .B1(new_n520), .B2(new_n724), .ZN(new_n1107));
  AOI211_X1 g0907(.A(G45), .B(new_n723), .C1(G68), .C2(G77), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT112), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n316), .A2(new_n288), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT50), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1110), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n803), .B1(new_n233), .B2(new_n259), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n808), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n788), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n835), .A2(G77), .ZN(new_n1119));
  INV_X1    g0919(.A(G159), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n815), .A2(new_n1120), .B1(new_n288), .B2(new_n816), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n651), .A2(new_n846), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n579), .C1(new_n280), .C2(new_n901), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n820), .A2(new_n361), .B1(new_n277), .B2(new_n822), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1079), .A2(new_n1119), .A3(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT113), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n579), .B1(G326), .B2(new_n827), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G311), .A2(new_n850), .B1(new_n819), .B2(G303), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n814), .A2(G322), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1129), .B(new_n1130), .C1(new_n1080), .C2(new_n816), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT48), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n835), .A2(G294), .B1(G283), .B2(new_n846), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT114), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT49), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1128), .B1(new_n454), .B2(new_n842), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1127), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1106), .B(new_n1118), .C1(new_n1141), .C2(new_n807), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT111), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1049), .B2(new_n786), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1050), .A2(KEYINPUT111), .A3(new_n787), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1105), .A2(new_n1146), .ZN(G393));
  AOI21_X1  g0947(.A(new_n786), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n407), .B1(G143), .B2(new_n827), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n892), .B(new_n1149), .C1(new_n361), .C2(new_n836), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT115), .Z(new_n1151));
  AOI22_X1  g0951(.A1(G150), .A2(new_n814), .B1(new_n853), .B2(G159), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT51), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n825), .A2(new_n323), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n819), .B2(new_n316), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n201), .B2(new_n822), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1151), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n815), .A2(new_n1080), .B1(new_n848), .B2(new_n816), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT52), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n245), .B1(new_n827), .B2(G322), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n454), .B2(new_n825), .C1(new_n820), .C2(new_n550), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G303), .B2(new_n850), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1159), .B(new_n1162), .C1(new_n855), .C2(new_n836), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G107), .B2(new_n891), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n807), .B1(new_n1157), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1017), .A2(new_n795), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n809), .B1(G97), .B2(new_n724), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n803), .A2(new_n240), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n789), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1165), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1148), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n782), .A2(new_n1050), .A3(new_n1066), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n725), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1102), .A2(new_n1066), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(G390));
  OAI21_X1  g0975(.A(new_n708), .B1(new_n738), .B2(new_n747), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n935), .B1(new_n1176), .B2(new_n872), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n979), .A2(G330), .A3(new_n871), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n933), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n933), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n871), .B(new_n1180), .C1(new_n774), .C2(new_n776), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n979), .A2(G330), .A3(new_n984), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n871), .B1(new_n774), .B2(new_n776), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n933), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n874), .A2(new_n935), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1182), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n452), .A2(new_n979), .A3(G330), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n928), .A2(new_n670), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n968), .A2(new_n969), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n971), .B2(new_n936), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n976), .A2(new_n971), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1198), .A3(new_n1181), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1187), .A2(new_n1180), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n970), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1201), .A2(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1199), .B1(new_n1202), .B2(new_n1183), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1193), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1183), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1206), .A2(new_n1189), .A3(new_n1199), .A4(new_n1192), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n725), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1205), .B1(new_n1202), .B2(new_n1181), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1194), .A2(new_n914), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n916), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n788), .B1(new_n316), .B2(new_n1211), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n815), .A2(new_n855), .B1(new_n454), .B2(new_n816), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n245), .B(new_n1154), .C1(G294), .C2(new_n827), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n457), .B2(new_n820), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G107), .C2(new_n850), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n899), .C1(new_n307), .C2(new_n836), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n253), .B1(new_n827), .B2(G125), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n842), .B2(new_n201), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT116), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n835), .A2(G150), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT53), .Z(new_n1222));
  INV_X1    g1022(.A(G128), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n815), .A2(new_n1223), .B1(new_n902), .B2(new_n816), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT117), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(KEYINPUT54), .B(G143), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n820), .A2(new_n1226), .B1(new_n1120), .B2(new_n825), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G137), .B2(new_n850), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1222), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1217), .B1(new_n1220), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1212), .B1(new_n1230), .B2(new_n807), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1209), .A2(new_n787), .B1(new_n1210), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1208), .A2(new_n1232), .ZN(G378));
  NAND3_X1  g1033(.A1(new_n667), .A2(new_n668), .A3(new_n292), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n941), .A2(new_n291), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n667), .A2(new_n668), .A3(new_n292), .A4(new_n1235), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1003), .B2(new_n775), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n974), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1242), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n996), .A2(G330), .A3(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1244), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n787), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n891), .A2(G58), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n815), .A2(new_n454), .B1(new_n520), .B2(new_n816), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1085), .B1(new_n855), .B2(new_n901), .C1(new_n822), .C2(new_n457), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n820), .A2(new_n611), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n407), .A2(new_n258), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1250), .A2(new_n1119), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT58), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1254), .B(new_n288), .C1(G33), .C2(G41), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n814), .A2(G125), .B1(G150), .B2(new_n846), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1261), .B1(new_n1223), .B2(new_n816), .C1(new_n836), .C2(new_n1226), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G132), .A2(new_n850), .B1(new_n819), .B2(G137), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT118), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT59), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT119), .ZN(new_n1267));
  AOI211_X1 g1067(.A(G33), .B(G41), .C1(new_n827), .C2(G124), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n842), .B2(new_n1120), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT120), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1267), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1266), .A2(KEYINPUT119), .ZN(new_n1274));
  OAI221_X1 g1074(.A(new_n1260), .B1(new_n1257), .B2(new_n1256), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n807), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1242), .A2(new_n914), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n788), .B1(new_n202), .B2(new_n1211), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(KEYINPUT121), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1249), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1191), .B1(new_n1209), .B2(new_n1189), .ZN(new_n1283));
  OAI21_X1  g1083(.A(KEYINPUT57), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n725), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1183), .B1(new_n1286), .B2(new_n1180), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1287), .A2(new_n1187), .B1(new_n1181), .B2(new_n1179), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1192), .B1(new_n1203), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1245), .B1(new_n996), .B2(G330), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n775), .B(new_n1242), .C1(new_n986), .C2(new_n995), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n974), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT57), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1282), .B1(new_n1285), .B2(new_n1295), .ZN(G375));
  OAI22_X1  g1096(.A1(new_n815), .A2(new_n550), .B1(new_n855), .B2(new_n816), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(G116), .A2(new_n850), .B1(new_n819), .B2(G107), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n245), .B1(new_n827), .B2(G303), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1122), .A3(new_n1299), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n1297), .B(new_n1300), .C1(G97), .C2(new_n835), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n836), .A2(new_n1120), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n579), .B1(new_n825), .B2(new_n288), .C1(new_n1223), .C2(new_n901), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n815), .A2(new_n902), .B1(new_n909), .B2(new_n816), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n820), .A2(new_n280), .B1(new_n822), .B2(new_n1226), .ZN(new_n1305));
  NOR4_X1   g1105(.A1(new_n1302), .A2(new_n1303), .A3(new_n1304), .A4(new_n1305), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1090), .A2(new_n1301), .B1(new_n1306), .B2(new_n1250), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n807), .ZN(new_n1308));
  OAI221_X1 g1108(.A(new_n788), .B1(G68), .B2(new_n1211), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n914), .B2(new_n933), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1189), .B2(new_n787), .ZN(new_n1311));
  XOR2_X1   g1111(.A(new_n1069), .B(KEYINPUT122), .Z(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1193), .A2(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1311), .B1(new_n1314), .B2(new_n1315), .ZN(G381));
  INV_X1    g1116(.A(G375), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1099), .B1(new_n1047), .B2(new_n1071), .ZN(new_n1318));
  INV_X1    g1118(.A(G378), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1105), .A2(new_n859), .A3(new_n1146), .ZN(new_n1320));
  NOR4_X1   g1120(.A1(new_n1320), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .A4(new_n1321), .ZN(G407));
  NAND2_X1  g1122(.A1(new_n1319), .A2(new_n706), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G407), .B(G213), .C1(G375), .C2(new_n1323), .ZN(G409));
  NAND2_X1  g1124(.A1(G393), .A2(G396), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1320), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1171), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1174), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n725), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1102), .B2(new_n1066), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1327), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(G387), .A2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1318), .A2(G390), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1326), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G387), .A2(new_n1331), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1318), .A2(G390), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1335), .A2(new_n1320), .A3(new_n1325), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1334), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT61), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1312), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1289), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT123), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1340), .A2(new_n1289), .A3(KEYINPUT123), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1282), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1319), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G378), .B(new_n1282), .C1(new_n1285), .C2(new_n1295), .ZN(new_n1347));
  AOI22_X1  g1147(.A1(new_n1346), .A2(new_n1347), .B1(G213), .B2(new_n706), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT60), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1349), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1350), .A2(new_n1315), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1287), .A2(new_n1187), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1352), .A2(KEYINPUT60), .A3(new_n1191), .A4(new_n1182), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n725), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1311), .B1(new_n1351), .B2(new_n1354), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n890), .A2(new_n918), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(G384), .B(new_n1311), .C1(new_n1351), .C2(new_n1354), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n706), .A2(G213), .A3(G2897), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1357), .A2(new_n1358), .A3(new_n1360), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1338), .B(new_n1339), .C1(new_n1348), .C2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n706), .A2(G213), .ZN(new_n1367));
  AND2_X1   g1167(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1347), .ZN(new_n1369));
  AOI21_X1  g1169(.A(KEYINPUT123), .B1(new_n1340), .B2(new_n1289), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1370), .A2(new_n1281), .ZN(new_n1371));
  AOI21_X1  g1171(.A(G378), .B1(new_n1371), .B2(new_n1344), .ZN(new_n1372));
  OAI211_X1 g1172(.A(new_n1367), .B(new_n1368), .C1(new_n1369), .C2(new_n1372), .ZN(new_n1373));
  XOR2_X1   g1173(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n1374));
  NAND3_X1  g1174(.A1(new_n1373), .A2(KEYINPUT125), .A3(new_n1374), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1348), .A2(KEYINPUT62), .A3(new_n1368), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1375), .A2(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(KEYINPUT125), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1366), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT126), .ZN(new_n1380));
  OAI21_X1  g1180(.A(new_n1367), .B1(new_n1369), .B2(new_n1372), .ZN(new_n1381));
  AND3_X1   g1181(.A1(new_n1357), .A2(new_n1358), .A3(new_n1360), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1360), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1383));
  NOR2_X1   g1183(.A1(new_n1382), .A2(new_n1383), .ZN(new_n1384));
  AOI21_X1  g1184(.A(KEYINPUT61), .B1(new_n1381), .B2(new_n1384), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1348), .A2(KEYINPUT63), .A3(new_n1368), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT63), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1373), .A2(new_n1387), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1385), .A2(new_n1386), .A3(new_n1388), .ZN(new_n1389));
  INV_X1    g1189(.A(new_n1338), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1389), .A2(new_n1390), .ZN(new_n1391));
  AND3_X1   g1191(.A1(new_n1379), .A2(new_n1380), .A3(new_n1391), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1380), .B1(new_n1379), .B2(new_n1391), .ZN(new_n1393));
  NOR2_X1   g1193(.A1(new_n1392), .A2(new_n1393), .ZN(G405));
  INV_X1    g1194(.A(KEYINPUT127), .ZN(new_n1395));
  NOR2_X1   g1195(.A1(new_n1368), .A2(new_n1395), .ZN(new_n1396));
  XNOR2_X1  g1196(.A(new_n1338), .B(new_n1396), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(G375), .A2(new_n1319), .ZN(new_n1398));
  OAI211_X1 g1198(.A(new_n1398), .B(new_n1347), .C1(KEYINPUT127), .C2(new_n1359), .ZN(new_n1399));
  XOR2_X1   g1199(.A(new_n1397), .B(new_n1399), .Z(G402));
endmodule


