//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT2), .B(G113), .Z(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(new_n191), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT75), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(KEYINPUT75), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n200), .A2(new_n203), .A3(KEYINPUT75), .A4(G104), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n199), .B1(new_n209), .B2(KEYINPUT76), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n211), .A3(new_n207), .A4(new_n208), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n205), .A2(new_n199), .A3(new_n207), .A4(new_n208), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n210), .A2(new_n212), .B1(KEYINPUT4), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n206), .A2(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n208), .A2(new_n207), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT76), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n221), .A2(new_n212), .A3(KEYINPUT4), .A4(G101), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n198), .B1(new_n214), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(new_n207), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n213), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT5), .ZN(new_n228));
  OAI21_X1  g042(.A(G113), .B1(new_n189), .B2(KEYINPUT5), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n194), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G110), .B(G122), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n233), .ZN(new_n235));
  INV_X1    g049(.A(new_n198), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n221), .A2(G101), .A3(new_n212), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n213), .A2(KEYINPUT4), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n239), .B2(new_n222), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n235), .B1(new_n240), .B2(new_n231), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n234), .A2(new_n241), .A3(KEYINPUT6), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT6), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(new_n235), .C1(new_n240), .C2(new_n231), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G143), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT64), .ZN(new_n251));
  XNOR2_X1  g065(.A(G143), .B(G146), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n249), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n246), .A2(new_n248), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(G125), .A3(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n247), .A2(KEYINPUT1), .A3(G146), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n261), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n246), .A3(new_n248), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G125), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G224), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n269), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n242), .A2(new_n244), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n271), .A2(KEYINPUT7), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n260), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n260), .B2(new_n268), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n230), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n213), .A2(new_n226), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n194), .B(KEYINPUT80), .C1(new_n228), .C2(new_n229), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT81), .A4(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n233), .B(KEYINPUT8), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT81), .B1(new_n227), .B2(new_n230), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n277), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n288), .B2(new_n234), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n187), .B1(new_n273), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n273), .A2(new_n187), .A3(new_n289), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G478), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(KEYINPUT15), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n262), .A2(G143), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n247), .A2(G128), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT90), .B1(new_n301), .B2(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G134), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT86), .B1(new_n190), .B2(G122), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n312));
  INV_X1    g126(.A(G122), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G116), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT87), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n313), .B2(G116), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n190), .A2(KEYINPUT87), .A3(G122), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT88), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n315), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n315), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n203), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n319), .A2(KEYINPUT14), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n315), .B1(new_n319), .B2(KEYINPUT14), .ZN(new_n325));
  OAI21_X1  g139(.A(G107), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n310), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n315), .A2(new_n319), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT88), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n315), .A2(new_n319), .A3(new_n320), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G107), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT91), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT13), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n302), .B1(new_n303), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(KEYINPUT89), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n301), .B2(KEYINPUT13), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n309), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n336), .A2(new_n339), .B1(new_n308), .B2(new_n309), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n332), .A2(new_n333), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n333), .B1(new_n332), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n327), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g157(.A(KEYINPUT9), .B(G234), .Z(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT74), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT70), .B(G217), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n270), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n327), .B(new_n350), .C1(new_n341), .C2(new_n342), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G902), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n300), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI211_X1 g168(.A(G902), .B(new_n299), .C1(new_n349), .C2(new_n351), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G952), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G953), .ZN(new_n359));
  INV_X1    g173(.A(G234), .ZN(new_n360));
  INV_X1    g174(.A(G237), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(G902), .B(G953), .C1(new_n360), .C2(new_n361), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT92), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT21), .B(G898), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n267), .A2(G140), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT16), .ZN(new_n372));
  OR3_X1    g186(.A1(new_n267), .A2(KEYINPUT16), .A3(G140), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G146), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT71), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n373), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(new_n245), .ZN(new_n378));
  AOI211_X1 g192(.A(KEYINPUT72), .B(G146), .C1(new_n372), .C2(new_n373), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n361), .A2(new_n270), .A3(G214), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n247), .ZN(new_n383));
  INV_X1    g197(.A(G131), .ZN(new_n384));
  NOR2_X1   g198(.A1(G237), .A2(G953), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(G143), .A3(G214), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n383), .A2(KEYINPUT82), .A3(new_n384), .A4(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n386), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT84), .B1(new_n393), .B2(KEYINPUT17), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n384), .B1(new_n383), .B2(new_n386), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n388), .B2(new_n387), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n390), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(KEYINPUT17), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n381), .A2(new_n394), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(new_n206), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n383), .A2(new_n386), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n370), .A2(new_n371), .A3(new_n245), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n370), .A2(new_n371), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G146), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n404), .A2(new_n405), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n391), .A2(KEYINPUT18), .A3(G131), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n401), .A2(new_n403), .A3(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT19), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT19), .B1(new_n370), .B2(new_n371), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n245), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n374), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n418), .A2(new_n393), .B1(new_n409), .B2(new_n410), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT83), .B1(new_n419), .B2(new_n403), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n421));
  INV_X1    g235(.A(new_n403), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n417), .B1(new_n396), .B2(new_n390), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n421), .B(new_n422), .C1(new_n423), .C2(new_n411), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n413), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G475), .A2(G902), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n413), .A2(new_n425), .A3(KEYINPUT85), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n429), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT20), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n431), .A2(KEYINPUT20), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n401), .A2(new_n412), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n422), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n413), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n353), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n438), .A2(G475), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n297), .A2(new_n368), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n385), .A2(G210), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT27), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT26), .B(G101), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT28), .ZN(new_n449));
  INV_X1    g263(.A(G137), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT65), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G137), .ZN(new_n453));
  AND2_X1   g267(.A1(KEYINPUT11), .A2(G134), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT11), .A2(G134), .ZN(new_n456));
  NOR2_X1   g270(.A1(KEYINPUT11), .A2(G134), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(G137), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n384), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(new_n453), .A3(new_n309), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n384), .B1(G134), .B2(G137), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT1), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n252), .A2(G128), .B1(new_n463), .B2(new_n248), .ZN(new_n464));
  INV_X1    g278(.A(new_n265), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n459), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n455), .A2(new_n384), .A3(new_n458), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n384), .B1(new_n455), .B2(new_n458), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n253), .B1(new_n252), .B2(new_n249), .ZN(new_n470));
  AND4_X1   g284(.A1(new_n253), .A2(new_n246), .A3(new_n248), .A4(new_n249), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n259), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n466), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n198), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n255), .B(new_n259), .C1(new_n467), .C2(new_n468), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n236), .A3(new_n466), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(KEYINPUT69), .A3(new_n198), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n449), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n477), .A2(KEYINPUT28), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n448), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n473), .A2(KEYINPUT30), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n476), .A2(new_n484), .A3(new_n466), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n236), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n476), .A2(new_n236), .A3(new_n466), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n447), .B1(new_n488), .B2(new_n445), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT67), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n236), .B1(new_n476), .B2(new_n466), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT28), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n481), .A2(new_n490), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n446), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n482), .B(new_n353), .C1(new_n489), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G472), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT67), .B1(new_n474), .B2(new_n477), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n494), .B(new_n446), .C1(new_n498), .C2(new_n449), .ZN(new_n499));
  INV_X1    g313(.A(new_n485), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n484), .B1(new_n476), .B2(new_n466), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n198), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT66), .B(KEYINPUT31), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n502), .A2(new_n477), .A3(new_n445), .A4(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n486), .A2(new_n487), .A3(new_n446), .ZN(new_n505));
  NOR2_X1   g319(.A1(KEYINPUT66), .A2(KEYINPUT31), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n499), .B(new_n504), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G472), .A2(G902), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(KEYINPUT32), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n497), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT32), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI211_X1 g328(.A(KEYINPUT68), .B(KEYINPUT32), .C1(new_n507), .C2(new_n508), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n188), .B2(G128), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n518), .B(new_n519), .C1(G119), .C2(new_n262), .ZN(new_n520));
  XNOR2_X1  g334(.A(G119), .B(G128), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G110), .Z(new_n522));
  AOI22_X1  g336(.A1(new_n520), .A2(G110), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n375), .B2(new_n380), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT73), .B(G110), .ZN(new_n525));
  OAI22_X1  g339(.A1(new_n520), .A2(new_n525), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n406), .A3(new_n374), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G137), .ZN(new_n529));
  INV_X1    g343(.A(G221), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n530), .A2(new_n360), .A3(G953), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n529), .B(new_n531), .Z(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n524), .A2(new_n527), .A3(new_n532), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n346), .B1(G234), .B2(new_n353), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G902), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n353), .A3(new_n535), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT25), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n534), .A2(KEYINPUT25), .A3(new_n353), .A4(new_n535), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n539), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n516), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT79), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G140), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n270), .A2(G227), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n464), .A2(new_n465), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n227), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n265), .A2(KEYINPUT77), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n252), .A2(new_n556), .A3(new_n264), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n263), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n213), .A3(new_n226), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n469), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT12), .ZN(new_n561));
  INV_X1    g375(.A(new_n472), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n214), .B2(new_n223), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT10), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n263), .A2(new_n555), .A3(new_n557), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n564), .B1(new_n565), .B2(new_n227), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n266), .A2(KEYINPUT10), .A3(new_n213), .A4(new_n226), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n568), .A3(new_n469), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n552), .B1(new_n561), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n469), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n472), .B1(new_n239), .B2(new_n222), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n567), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n569), .A2(new_n574), .A3(new_n552), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n353), .B1(new_n570), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n469), .B1(new_n563), .B2(new_n568), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n572), .A2(new_n573), .A3(new_n571), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n551), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n561), .A2(new_n569), .A3(new_n552), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT78), .B(G469), .ZN(new_n582));
  AOI22_X1  g396(.A1(G469), .A2(new_n576), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n530), .B1(new_n345), .B2(new_n353), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n548), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n581), .A2(new_n582), .ZN(new_n587));
  INV_X1    g401(.A(G469), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n560), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n551), .B1(new_n590), .B2(new_n578), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n569), .A2(new_n574), .A3(new_n552), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n588), .B1(new_n593), .B2(new_n353), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT79), .B(new_n586), .C1(new_n587), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n441), .A2(new_n547), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n292), .A2(KEYINPUT94), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n295), .B1(new_n600), .B2(new_n290), .ZN(new_n601));
  AOI211_X1 g415(.A(KEYINPUT94), .B(new_n187), .C1(new_n273), .C2(new_n289), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n291), .A2(KEYINPUT94), .A3(new_n292), .ZN(new_n604));
  INV_X1    g418(.A(new_n602), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(KEYINPUT95), .A3(new_n295), .A4(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n507), .A2(new_n353), .ZN(new_n608));
  NAND2_X1  g422(.A1(KEYINPUT93), .A2(G472), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n585), .B2(new_n595), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n545), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n298), .A2(G902), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n349), .A2(new_n615), .A3(new_n351), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n349), .B2(new_n351), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n352), .A2(new_n353), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT96), .B(G478), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n367), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n623), .B(new_n624), .C1(new_n434), .C2(new_n439), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n613), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT20), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n413), .A2(new_n425), .A3(KEYINPUT85), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT85), .B1(new_n413), .B2(new_n425), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n630), .B1(new_n633), .B2(new_n429), .ZN(new_n634));
  NOR4_X1   g448(.A1(new_n631), .A2(new_n632), .A3(KEYINPUT20), .A4(new_n432), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n631), .A2(new_n632), .A3(new_n432), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n630), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n431), .A2(KEYINPUT20), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT97), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n356), .A2(new_n439), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n624), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT98), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n641), .A2(new_n645), .A3(new_n624), .A4(new_n642), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n613), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  AND2_X1   g464(.A1(new_n544), .A2(new_n537), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n528), .B(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n538), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n441), .A2(new_n612), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  XNOR2_X1  g473(.A(KEYINPUT99), .B(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n365), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n362), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n641), .A2(new_n642), .A3(new_n656), .A4(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n514), .A2(new_n515), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n507), .A2(new_n508), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n666), .A2(KEYINPUT32), .B1(new_n496), .B2(G472), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n585), .A2(new_n595), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n607), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XOR2_X1   g484(.A(new_n293), .B(KEYINPUT38), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n426), .A2(new_n433), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n672), .B1(new_n637), .B2(new_n630), .ZN(new_n673));
  INV_X1    g487(.A(new_n439), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n356), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR4_X1   g490(.A1(new_n671), .A2(new_n676), .A3(new_n296), .A4(new_n656), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n662), .B(KEYINPUT39), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n596), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n445), .B1(new_n486), .B2(new_n487), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n478), .A2(new_n479), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n682), .B(new_n353), .C1(new_n683), .C2(new_n445), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G472), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n509), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n681), .B1(new_n665), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n512), .A2(new_n513), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT68), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n512), .A2(new_n511), .A3(new_n513), .ZN(new_n690));
  AND4_X1   g504(.A1(new_n681), .A2(new_n689), .A3(new_n690), .A4(new_n686), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n677), .A2(new_n680), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NAND3_X1  g510(.A1(new_n667), .A2(new_n689), .A3(new_n690), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n596), .A2(new_n603), .A3(new_n697), .A4(new_n606), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n673), .A2(new_n674), .B1(new_n622), .B2(new_n618), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n656), .A3(new_n662), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT101), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n623), .B1(new_n434), .B2(new_n439), .ZN(new_n703));
  INV_X1    g517(.A(new_n662), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n703), .A2(new_n655), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n607), .A2(new_n702), .A3(new_n668), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  NOR3_X1   g522(.A1(new_n590), .A2(new_n578), .A3(new_n551), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n552), .B1(new_n569), .B2(new_n574), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n353), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n581), .A2(new_n582), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n586), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n603), .A2(new_n606), .A3(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n516), .A2(new_n625), .A3(new_n546), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT102), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n603), .A2(new_n606), .A3(new_n715), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n697), .A2(new_n699), .A3(new_n624), .A4(new_n545), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND4_X1  g539(.A1(new_n603), .A2(new_n606), .A3(new_n697), .A4(new_n715), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n644), .A3(new_n545), .A4(new_n646), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NAND3_X1  g543(.A1(new_n368), .A2(new_n440), .A3(new_n656), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n188), .ZN(G21));
  NAND2_X1  g546(.A1(new_n608), .A2(G472), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n480), .A2(new_n481), .A3(new_n445), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n508), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n545), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n712), .A2(new_n713), .A3(new_n624), .A4(new_n586), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n603), .A2(new_n739), .A3(new_n606), .A4(new_n675), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  AND2_X1   g555(.A1(new_n733), .A2(new_n736), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n699), .A2(new_n656), .A3(new_n662), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n716), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  NOR2_X1   g560(.A1(new_n293), .A2(new_n296), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n575), .B1(new_n570), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n591), .A2(KEYINPUT104), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(G469), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(G469), .A2(G902), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT103), .Z(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n713), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n747), .A2(new_n586), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n703), .A2(new_n704), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n688), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n512), .A2(KEYINPUT105), .A3(new_n513), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n667), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n756), .A2(new_n757), .A3(new_n545), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n747), .A2(new_n586), .A3(new_n755), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n516), .A3(new_n546), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n703), .A2(KEYINPUT42), .A3(new_n704), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n762), .A2(KEYINPUT42), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NOR3_X1   g581(.A1(new_n634), .A2(new_n635), .A3(new_n629), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT97), .B1(new_n638), .B2(new_n639), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n642), .B(new_n662), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT106), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n764), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  INV_X1    g589(.A(new_n623), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n439), .A3(new_n434), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT43), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n611), .A3(new_n656), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n747), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n678), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n749), .A2(KEYINPUT45), .A3(new_n750), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n588), .B1(new_n593), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n753), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n713), .B1(new_n788), .B2(KEYINPUT46), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n586), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n784), .B(new_n791), .C1(new_n779), .C2(new_n780), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT107), .B(new_n747), .C1(new_n779), .C2(new_n780), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n783), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  XNOR2_X1  g609(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n791), .B(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n747), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n697), .A2(new_n798), .A3(new_n545), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n757), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NAND2_X1  g615(.A1(new_n712), .A2(new_n713), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT110), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n671), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n545), .A2(new_n295), .A3(new_n586), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n777), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT109), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(KEYINPUT109), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n805), .A2(new_n692), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n698), .A2(new_n663), .B1(new_n720), .B2(new_n743), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n755), .A2(new_n655), .A3(new_n586), .A4(new_n662), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n689), .A2(new_n686), .A3(new_n690), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT100), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n665), .A2(new_n681), .A3(new_n686), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n603), .A2(new_n606), .A3(new_n675), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND4_X1   g635(.A1(KEYINPUT114), .A2(new_n707), .A3(new_n814), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n815), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n687), .B2(new_n691), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n603), .A2(new_n606), .A3(new_n675), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n813), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT114), .B1(new_n827), .B2(new_n707), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n812), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n814), .A2(KEYINPUT113), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n814), .A2(KEYINPUT113), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n707), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n642), .A2(new_n673), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n703), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n546), .A2(new_n367), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n612), .A2(new_n297), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n597), .A2(new_n657), .A3(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n357), .A2(new_n439), .A3(new_n704), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n641), .A3(new_n747), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n641), .A3(KEYINPUT112), .A4(new_n747), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n656), .A3(new_n668), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n744), .A2(new_n756), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n766), .A2(new_n774), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n740), .B1(new_n726), .B2(new_n730), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n723), .A2(new_n728), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT111), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n849), .B1(new_n722), .B2(new_n718), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(KEYINPUT111), .A3(new_n728), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n840), .B(new_n848), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n835), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n840), .ZN(new_n859));
  INV_X1    g673(.A(new_n848), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n854), .A2(KEYINPUT111), .A3(new_n728), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT111), .B1(new_n854), .B2(new_n728), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n832), .B1(new_n822), .B2(new_n828), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n701), .A2(new_n706), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n669), .A2(new_n745), .A3(new_n821), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n827), .A2(KEYINPUT114), .A3(new_n707), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(KEYINPUT52), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n863), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n858), .B(KEYINPUT54), .C1(new_n871), .C2(new_n857), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n840), .A2(new_n857), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n860), .A2(new_n728), .A3(new_n874), .A4(new_n854), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n835), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n873), .B(new_n877), .C1(new_n871), .C2(KEYINPUT53), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n798), .A2(new_n546), .A3(new_n362), .A4(new_n714), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n692), .A3(new_n699), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT43), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n777), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n737), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n777), .A2(new_n881), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n882), .A2(new_n363), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n359), .B(new_n880), .C1(new_n885), .C2(new_n720), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n778), .A2(new_n363), .A3(new_n715), .A4(new_n747), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n761), .A2(new_n545), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n887), .A2(KEYINPUT48), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT48), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n879), .A2(new_n692), .A3(new_n440), .A4(new_n776), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n656), .A2(new_n742), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n885), .A2(new_n798), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n712), .A2(new_n584), .A3(new_n713), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n797), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n895), .A2(KEYINPUT51), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT50), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n671), .A2(new_n296), .A3(new_n715), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n901), .B1(new_n885), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n885), .A2(new_n901), .A3(new_n902), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n891), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n899), .A2(KEYINPUT116), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n894), .B1(new_n899), .B2(KEYINPUT116), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n906), .A2(KEYINPUT117), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n904), .A2(new_n911), .A3(new_n905), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n908), .B(new_n909), .C1(new_n910), .C2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n872), .A2(new_n878), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n872), .A2(new_n878), .A3(new_n915), .A4(KEYINPUT118), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n358), .A2(new_n270), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT119), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n811), .B1(new_n918), .B2(new_n922), .ZN(G75));
  NAND2_X1  g737(.A1(new_n864), .A2(new_n870), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT53), .B1(new_n924), .B2(new_n856), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n875), .B1(new_n829), .B2(new_n834), .ZN(new_n926));
  OAI211_X1 g740(.A(G210), .B(G902), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n242), .A2(new_n244), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n272), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(KEYINPUT120), .B2(new_n928), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n927), .A2(new_n928), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n927), .B2(new_n928), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n270), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  XNOR2_X1  g751(.A(new_n753), .B(KEYINPUT57), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n868), .A2(KEYINPUT52), .A3(new_n869), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT52), .B1(new_n868), .B2(new_n869), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n857), .B1(new_n941), .B2(new_n863), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n873), .B1(new_n942), .B2(new_n877), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n925), .A2(KEYINPUT54), .A3(new_n926), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n579), .A2(new_n580), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n924), .A2(new_n856), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n926), .B1(new_n948), .B2(new_n857), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n353), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n785), .A3(new_n787), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n936), .B1(new_n947), .B2(new_n951), .ZN(G54));
  INV_X1    g766(.A(new_n936), .ZN(new_n953));
  NAND2_X1  g767(.A1(KEYINPUT58), .A2(G475), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT121), .ZN(new_n955));
  OAI211_X1 g769(.A(G902), .B(new_n955), .C1(new_n925), .C2(new_n926), .ZN(new_n956));
  INV_X1    g770(.A(new_n633), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n956), .ZN(new_n959));
  OAI21_X1  g773(.A(KEYINPUT122), .B1(new_n959), .B2(new_n633), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n956), .A2(new_n961), .A3(new_n957), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n958), .B1(new_n960), .B2(new_n962), .ZN(G60));
  OR2_X1    g777(.A1(new_n616), .A2(new_n617), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n872), .A2(new_n878), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT59), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n964), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n964), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT54), .B1(new_n925), .B2(new_n926), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n878), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n969), .A2(new_n936), .A3(new_n972), .ZN(G63));
  INV_X1    g787(.A(new_n536), .ZN(new_n974));
  XNOR2_X1  g788(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n974), .B1(new_n949), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n653), .B(new_n977), .C1(new_n925), .C2(new_n926), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n953), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n979), .A2(KEYINPUT61), .A3(new_n953), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G66));
  INV_X1    g799(.A(G224), .ZN(new_n986));
  OAI21_X1  g800(.A(G953), .B1(new_n366), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n840), .B1(new_n853), .B2(new_n855), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(G953), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n929), .B1(G898), .B2(new_n270), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT124), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n989), .B(new_n991), .ZN(G69));
  NAND2_X1  g806(.A1(new_n483), .A2(new_n485), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT125), .Z(new_n994));
  NOR2_X1   g808(.A1(new_n414), .A2(new_n415), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n994), .B(new_n995), .Z(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT126), .Z(new_n997));
  INV_X1    g811(.A(new_n679), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n998), .A2(new_n547), .A3(new_n747), .A4(new_n837), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n794), .A2(new_n800), .A3(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n830), .A2(new_n707), .A3(new_n831), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n695), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1001), .A2(KEYINPUT62), .A3(new_n695), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n997), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  OR4_X1    g821(.A1(new_n784), .A2(new_n791), .A3(new_n825), .A4(new_n888), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n766), .A2(new_n800), .A3(new_n774), .A4(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n794), .A2(new_n1009), .A3(new_n1001), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n270), .ZN(new_n1011));
  INV_X1    g825(.A(new_n996), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(G900), .B2(G953), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n1014));
  AOI22_X1  g828(.A1(new_n1011), .A2(new_n1013), .B1(KEYINPUT127), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1007), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1014), .A2(KEYINPUT127), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(G72));
  NOR2_X1   g832(.A1(new_n488), .A2(new_n445), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1019), .A2(new_n505), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT63), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n936), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n682), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n486), .A2(new_n487), .A3(new_n445), .ZN(new_n1025));
  AOI22_X1  g839(.A1(new_n1006), .A2(new_n1024), .B1(new_n1010), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n988), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n948), .A2(KEYINPUT53), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n1029), .A2(new_n858), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G57));
endmodule


