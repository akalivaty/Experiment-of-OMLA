//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT66), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT64), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n218), .B1(new_n222), .B2(new_n223), .C1(new_n213), .C2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n215), .A2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(KEYINPUT76), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT74), .ZN(new_n242));
  INV_X1    g0042(.A(KEYINPUT69), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n243), .B1(new_n206), .B2(new_n244), .ZN(new_n245));
  NAND4_X1  g0045(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n245), .A2(new_n219), .A3(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(KEYINPUT70), .A3(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G77), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G68), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n248), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT11), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT67), .B(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT12), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G68), .ZN(new_n266));
  INV_X1    g0066(.A(new_n265), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(KEYINPUT12), .A3(new_n256), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n266), .B(new_n268), .C1(new_n258), .C2(KEYINPUT11), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT14), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n219), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G226), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G232), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n278), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n276), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G97), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n273), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT13), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(new_n293), .A3(G274), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n260), .A2(new_n292), .B1(new_n220), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n297), .B2(G238), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n288), .A2(new_n289), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n289), .B1(new_n288), .B2(new_n298), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n271), .B(G169), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n273), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n244), .ZN(new_n304));
  NAND2_X1  g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(G226), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n306), .B1(new_n310), .B2(new_n283), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n302), .B1(new_n311), .B2(new_n286), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n260), .A2(new_n292), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n313), .A2(new_n302), .A3(G238), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n294), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT13), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n288), .A2(new_n298), .A3(new_n289), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G179), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n301), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n271), .B1(new_n320), .B2(G169), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT73), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(G169), .B1(new_n299), .B2(new_n300), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT14), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n318), .A4(new_n301), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n270), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n320), .A2(G200), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n316), .A2(G190), .A3(new_n317), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n270), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n242), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT16), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n306), .B2(G20), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n249), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n256), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G58), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n256), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n201), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n255), .A2(G159), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n333), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n306), .A2(new_n334), .A3(G20), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT7), .B1(new_n276), .B2(new_n249), .ZN(new_n345));
  OAI21_X1  g0145(.A(G68), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n342), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n348), .A3(new_n247), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n265), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n262), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n351), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n295), .B1(new_n297), .B2(G232), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n306), .A2(G226), .A3(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n307), .A2(new_n308), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT75), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n306), .A2(new_n360), .A3(new_n361), .A4(G223), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n279), .B(new_n280), .C1(new_n274), .C2(new_n275), .ZN(new_n363));
  INV_X1    g0163(.A(G223), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT75), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n359), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n356), .B1(new_n366), .B2(new_n302), .ZN(new_n367));
  INV_X1    g0167(.A(G169), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(new_n356), .C1(new_n366), .C2(new_n302), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n355), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT18), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n367), .A2(G200), .ZN(new_n374));
  OAI211_X1 g0174(.A(G190), .B(new_n356), .C1(new_n366), .C2(new_n302), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n374), .A2(new_n349), .A3(new_n354), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT17), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n349), .A2(new_n354), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n379), .A2(KEYINPUT17), .A3(new_n375), .A4(new_n374), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n355), .A2(new_n381), .A3(new_n369), .A4(new_n371), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n373), .A2(new_n378), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n306), .A2(G238), .A3(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n276), .A2(G107), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(new_n282), .C2(new_n363), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n273), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n295), .B1(new_n297), .B2(G244), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G200), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G20), .A2(G77), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n351), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G87), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT15), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT15), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT15), .B(G87), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n391), .B(new_n394), .C1(new_n404), .C2(new_n250), .ZN(new_n405));
  INV_X1    g0205(.A(G77), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(new_n247), .B1(new_n406), .B2(new_n267), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n387), .A2(G190), .A3(new_n388), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n353), .A2(G77), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n390), .A2(new_n407), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n247), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n267), .A2(new_n406), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n389), .A2(new_n368), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n387), .A2(new_n370), .A3(new_n388), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n306), .A2(new_n360), .A3(G222), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n306), .A2(G223), .A3(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(new_n419), .C1(new_n406), .C2(new_n306), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n273), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n295), .B1(new_n297), .B2(G226), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n370), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n265), .A2(G50), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n255), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n252), .A2(new_n253), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n426), .B1(new_n427), .B2(new_n350), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n425), .B1(new_n428), .B2(new_n247), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n248), .A2(G50), .A3(new_n261), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n424), .B(new_n431), .C1(G169), .C2(new_n423), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT10), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n429), .A2(KEYINPUT9), .A3(new_n430), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n421), .A2(G190), .A3(new_n422), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT9), .B1(new_n429), .B2(new_n430), .ZN(new_n438));
  INV_X1    g0238(.A(G200), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(new_n421), .B2(new_n422), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n433), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  NOR4_X1   g0242(.A1(new_n436), .A2(new_n438), .A3(new_n440), .A4(KEYINPUT10), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n417), .B(new_n432), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n383), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n332), .A2(new_n445), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n327), .A2(new_n242), .A3(new_n331), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n241), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n322), .A2(new_n326), .ZN(new_n449));
  INV_X1    g0249(.A(new_n270), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n331), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT74), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT76), .A3(new_n332), .A4(new_n445), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n267), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(G33), .B2(G283), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n244), .A2(G97), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n457), .A2(new_n458), .B1(G20), .B2(new_n455), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n247), .A2(KEYINPUT20), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT20), .B1(new_n247), .B2(new_n459), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n260), .A2(G33), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n248), .A2(new_n265), .A3(new_n462), .ZN(new_n463));
  OAI221_X1 g0263(.A(new_n456), .B1(new_n460), .B2(new_n461), .C1(new_n455), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G257), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n304), .B2(new_n305), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(new_n360), .B1(new_n276), .B2(G303), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n306), .A2(G264), .A3(G1698), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n273), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT67), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G41), .ZN(new_n475));
  AND4_X1   g0275(.A1(G45), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(G274), .B1(new_n474), .B2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n273), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n478), .A3(KEYINPUT80), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n471), .A2(new_n473), .A3(new_n475), .A4(G45), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(G274), .C1(new_n272), .C2(new_n219), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n482), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n302), .B(G270), .C1(new_n481), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n470), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G190), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n464), .B(new_n490), .C1(G200), .C2(new_n488), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(new_n487), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n302), .B1(new_n467), .B2(new_n468), .ZN(new_n493));
  OAI211_X1 g0293(.A(KEYINPUT21), .B(G169), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n470), .A2(new_n485), .A3(G179), .A4(new_n487), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n464), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n464), .A2(new_n488), .A3(G169), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT84), .B(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n249), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT22), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT22), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n306), .A2(new_n505), .A3(new_n249), .A4(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT24), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n250), .A2(new_n455), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT23), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n249), .B2(G107), .ZN(new_n511));
  INV_X1    g0311(.A(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n508), .B1(new_n507), .B2(new_n514), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n247), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g0318(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n519));
  NAND3_X1  g0319(.A1(new_n267), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT85), .B(KEYINPUT25), .C1(new_n265), .C2(G107), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n463), .C2(new_n512), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n273), .B1(new_n476), .B2(new_n482), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G294), .ZN(new_n527));
  INV_X1    g0327(.A(G250), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n363), .C2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n525), .A2(G264), .B1(new_n529), .B2(new_n273), .ZN(new_n530));
  AOI21_X1  g0330(.A(G200), .B1(new_n530), .B2(new_n485), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n525), .A2(G264), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n273), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n485), .A3(new_n534), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n531), .A2(new_n532), .B1(G190), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n530), .A2(KEYINPUT86), .A3(new_n489), .A4(new_n485), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n524), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(new_n370), .A3(new_n485), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n368), .ZN(new_n540));
  INV_X1    g0340(.A(new_n517), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n248), .B1(new_n541), .B2(new_n515), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n540), .C1(new_n542), .C2(new_n522), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT79), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  OAI211_X1 g0347(.A(G250), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n548));
  OAI21_X1  g0348(.A(G244), .B1(new_n274), .B2(new_n275), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n279), .A2(KEYINPUT4), .A3(new_n280), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n552));
  INV_X1    g0352(.A(G244), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n304), .B2(new_n305), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n552), .B1(new_n554), .B2(new_n360), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n546), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g0356(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n557));
  NAND2_X1  g0357(.A1(new_n279), .A2(new_n280), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n549), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n554), .A2(KEYINPUT4), .A3(new_n360), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n528), .A2(new_n278), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n306), .A2(new_n561), .B1(G33), .B2(G283), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n559), .A2(new_n560), .A3(new_n562), .A4(KEYINPUT79), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n273), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(G257), .A2(new_n525), .B1(new_n479), .B2(new_n484), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n370), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  NOR2_X1   g0367(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G97), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(KEYINPUT6), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(G20), .C1(new_n567), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n255), .A2(G77), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n512), .B1(new_n335), .B2(new_n336), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n247), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n265), .A2(G97), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n248), .A2(new_n265), .A3(new_n462), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n302), .B(G257), .C1(new_n481), .C2(new_n486), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT80), .B1(new_n476), .B2(new_n478), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n481), .A2(new_n483), .A3(new_n480), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n302), .B1(new_n586), .B2(new_n546), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n587), .B2(new_n563), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n566), .B(new_n581), .C1(new_n588), .C2(G169), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n564), .A2(G190), .A3(new_n565), .ZN(new_n590));
  INV_X1    g0390(.A(new_n578), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n463), .B2(new_n571), .ZN(new_n592));
  OAI21_X1  g0392(.A(G107), .B1(new_n344), .B2(new_n345), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n573), .A3(new_n574), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n247), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n590), .B(new_n595), .C1(new_n588), .C2(new_n439), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n250), .B2(new_n571), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT83), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n306), .A2(new_n249), .A3(G68), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT83), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n597), .C1(new_n250), .C2(new_n571), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(G20), .B1(new_n287), .B2(KEYINPUT19), .ZN(new_n604));
  OR4_X1    g0404(.A1(KEYINPUT82), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n395), .A2(new_n571), .A3(new_n512), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT82), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n247), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n404), .A2(new_n267), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n609), .B(new_n610), .C1(new_n395), .C2(new_n463), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n244), .A2(new_n455), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n554), .B2(G1698), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n306), .A2(new_n360), .A3(G238), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n302), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n471), .A2(new_n473), .A3(G45), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n528), .ZN(new_n617));
  INV_X1    g0417(.A(G274), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n260), .A2(G45), .A3(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n617), .A2(new_n619), .A3(new_n302), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n615), .A2(new_n620), .A3(new_n489), .ZN(new_n621));
  INV_X1    g0421(.A(G238), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n363), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n612), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n549), .B2(new_n278), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n273), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n617), .A2(new_n619), .A3(new_n302), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n439), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OR3_X1    g0428(.A1(new_n611), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(G169), .B1(new_n626), .B2(new_n627), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT81), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n370), .A3(new_n627), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n609), .B(new_n610), .C1(new_n404), .C2(new_n463), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n615), .A2(new_n620), .A3(G179), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT81), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n589), .A2(new_n596), .A3(new_n629), .A4(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n454), .A2(new_n502), .A3(new_n545), .A4(new_n638), .ZN(G372));
  AND2_X1   g0439(.A1(new_n373), .A2(new_n382), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n327), .B1(new_n330), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n378), .A2(new_n380), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n442), .A2(new_n443), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n432), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n404), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n579), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n651), .A2(new_n610), .A3(new_n609), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT87), .B1(new_n635), .B2(new_n630), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n368), .B1(new_n615), .B2(new_n620), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT87), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n632), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n564), .A2(new_n370), .A3(new_n565), .ZN(new_n658));
  AOI21_X1  g0458(.A(G169), .B1(new_n564), .B2(new_n565), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n658), .A2(new_n659), .A3(new_n595), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n629), .A3(new_n637), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n611), .A2(new_n621), .A3(new_n628), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n657), .A2(new_n589), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n596), .A2(new_n589), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n497), .A2(new_n500), .A3(new_n543), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n657), .A2(new_n663), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n532), .B1(new_n535), .B2(new_n439), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n535), .A2(G190), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n537), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n524), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n668), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n662), .B(new_n666), .C1(new_n667), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n454), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n649), .A2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(G213), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT27), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n249), .A2(G13), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n260), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT88), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n680), .B1(new_n260), .B2(new_n681), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n464), .ZN(new_n692));
  MUX2_X1   g0492(.A(new_n501), .B(new_n502), .S(new_n692), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n524), .A2(new_n691), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n545), .A2(new_n696), .B1(new_n544), .B2(new_n691), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n691), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n545), .A2(new_n501), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n543), .B2(new_n691), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT91), .Z(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  NAND3_X1  g0504(.A1(new_n605), .A2(new_n455), .A3(new_n607), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n216), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(new_n709), .A3(G1), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n223), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n676), .A2(new_n713), .A3(new_n700), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n660), .A2(new_n665), .A3(new_n629), .A4(new_n637), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n654), .A2(new_n655), .A3(new_n632), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n655), .B1(new_n654), .B2(new_n632), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n634), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n715), .B(new_n718), .C1(new_n664), .C2(new_n665), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n629), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n538), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n667), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n596), .A2(new_n589), .A3(KEYINPUT92), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n721), .A2(new_n668), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n725), .B2(KEYINPUT93), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n596), .A2(new_n589), .A3(KEYINPUT92), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT92), .B1(new_n596), .B2(new_n589), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT93), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n729), .A2(new_n730), .A3(new_n668), .A4(new_n721), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n691), .B1(new_n726), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n714), .B1(new_n732), .B2(new_n713), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT30), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n564), .A2(new_n565), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n615), .A2(new_n620), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n530), .ZN(new_n738));
  OR4_X1    g0538(.A1(new_n735), .A2(new_n736), .A3(new_n738), .A4(new_n495), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(G179), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n736), .A2(new_n740), .A3(new_n488), .A4(new_n535), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n588), .A2(new_n530), .A3(new_n737), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n735), .B1(new_n742), .B2(new_n495), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT31), .B1(new_n744), .B2(new_n691), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n502), .A2(new_n545), .A3(new_n638), .A4(new_n700), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n734), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n733), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n712), .B1(new_n751), .B2(G1), .ZN(G364));
  AOI21_X1  g0552(.A(new_n293), .B1(new_n681), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n695), .B1(G330), .B2(new_n693), .C1(new_n708), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n708), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n306), .A2(new_n216), .ZN(new_n757));
  INV_X1    g0557(.A(G355), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n216), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n239), .A2(new_n291), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n707), .A2(new_n306), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n223), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(new_n291), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n219), .B1(G20), .B2(new_n368), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n756), .B1(new_n765), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n370), .A2(new_n439), .A3(KEYINPUT95), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT95), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G179), .B2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n249), .A2(G190), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT96), .B(KEYINPUT32), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n489), .B1(new_n773), .B2(new_n775), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n249), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n781), .A2(new_n782), .B1(G97), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n249), .A2(new_n370), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G200), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT94), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n489), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n786), .B1(new_n792), .B2(new_n202), .C1(new_n781), .C2(new_n782), .ZN(new_n793));
  INV_X1    g0593(.A(new_n787), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n794), .A2(G190), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n306), .B1(new_n796), .B2(new_n406), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n794), .A2(new_n489), .A3(G200), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(G58), .B2(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n249), .A2(new_n489), .A3(new_n439), .A4(G179), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n395), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n249), .A2(new_n439), .A3(G179), .A4(G190), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(G107), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n790), .A2(G190), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n799), .B(new_n804), .C1(new_n256), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n276), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G311), .B2(new_n795), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n778), .A2(G329), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n800), .A2(G303), .B1(new_n803), .B2(G283), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n791), .A2(G326), .B1(G294), .B2(new_n785), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT33), .B(G317), .Z(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n806), .B2(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n793), .A2(new_n807), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n772), .B1(new_n818), .B2(new_n769), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n768), .B(KEYINPUT97), .Z(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n693), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n755), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G396));
  NAND2_X1  g0623(.A1(new_n676), .A2(new_n700), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n691), .A2(new_n413), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n641), .B1(new_n825), .B2(new_n410), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n416), .A2(new_n691), .ZN(new_n827));
  OR3_X1    g0627(.A1(new_n826), .A2(KEYINPUT101), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT101), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n676), .A2(new_n830), .A3(new_n700), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n750), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n756), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n750), .A2(new_n832), .A3(new_n833), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n769), .A2(new_n766), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n756), .B1(new_n839), .B2(G77), .ZN(new_n840));
  INV_X1    g0640(.A(new_n803), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n801), .A2(new_n512), .B1(new_n841), .B2(new_n395), .ZN(new_n842));
  INV_X1    g0642(.A(G294), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n276), .B1(new_n796), .B2(new_n455), .C1(new_n843), .C2(new_n808), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n842), .B(new_n844), .C1(G311), .C2(new_n778), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n805), .A2(G283), .B1(G97), .B2(new_n785), .ZN(new_n846));
  INV_X1    g0646(.A(G303), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(new_n846), .C1(new_n847), .C2(new_n792), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT99), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G143), .A2(new_n798), .B1(new_n795), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n806), .B2(new_n851), .C1(new_n852), .C2(new_n792), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT34), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n801), .A2(new_n202), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n841), .A2(new_n256), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n338), .B2(new_n784), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT100), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n306), .B1(new_n779), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n863), .B1(new_n860), .B2(new_n862), .C1(new_n853), .C2(new_n854), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n849), .B1(new_n855), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n840), .B1(new_n865), .B2(new_n769), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n767), .B2(new_n830), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n837), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G384));
  INV_X1    g0669(.A(new_n222), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT35), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n570), .B1(new_n567), .B2(new_n572), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n870), .B(G116), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n871), .B2(new_n872), .ZN(new_n874));
  XNOR2_X1  g0674(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(G77), .B1(new_n338), .B2(new_n256), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n877), .A2(new_n223), .B1(G50), .B2(new_n256), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n260), .A2(G13), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n827), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n833), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n450), .A2(new_n691), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n451), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  INV_X1    g0687(.A(new_n689), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n383), .A2(new_n355), .A3(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n372), .B(new_n376), .C1(new_n379), .C2(new_n689), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n890), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n887), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n890), .B(KEYINPUT37), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n383), .A2(new_n355), .A3(new_n888), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n886), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n894), .B2(new_n895), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n327), .A2(new_n700), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n640), .A2(new_n888), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n898), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT103), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n723), .A2(new_n724), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT93), .B1(new_n911), .B2(new_n675), .ZN(new_n912));
  INV_X1    g0712(.A(new_n719), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n731), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n713), .B1(new_n914), .B2(new_n700), .ZN(new_n915));
  INV_X1    g0715(.A(new_n714), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n454), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n454), .B(KEYINPUT103), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n648), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n909), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n744), .A2(new_n691), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT31), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n749), .A3(new_n745), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n884), .A2(new_n926), .A3(new_n830), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n884), .A2(KEYINPUT104), .A3(new_n926), .A4(new_n830), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n897), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT40), .B1(new_n900), .B2(new_n901), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT105), .B1(new_n934), .B2(new_n927), .ZN(new_n935));
  INV_X1    g0735(.A(new_n926), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n831), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n932), .B1(new_n893), .B2(new_n896), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT105), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n884), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(G330), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n454), .A2(new_n750), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT106), .Z(new_n945));
  AOI22_X1  g0745(.A1(new_n931), .A2(new_n932), .B1(new_n935), .B2(new_n940), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n946), .A2(new_n454), .A3(new_n926), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n922), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n260), .B2(new_n681), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n945), .A2(new_n922), .A3(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n880), .B1(new_n949), .B2(new_n950), .ZN(G367));
  AND2_X1   g0751(.A1(new_n691), .A2(new_n611), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n720), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n657), .A2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT107), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n955), .B2(new_n954), .ZN(new_n958));
  INV_X1    g0758(.A(new_n820), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n806), .A2(new_n780), .B1(new_n202), .B2(new_n796), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n841), .A2(new_n406), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n306), .B1(new_n338), .B2(new_n801), .C1(new_n808), .C2(new_n851), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(G137), .C2(new_n778), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(KEYINPUT112), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n791), .A2(G143), .B1(G68), .B2(new_n785), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n962), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(G283), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n276), .B1(new_n796), .B2(new_n969), .C1(new_n847), .C2(new_n808), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G97), .B2(new_n803), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n778), .A2(G317), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT46), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n800), .A2(G116), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n973), .B2(new_n974), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n785), .A2(G107), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G294), .A2(new_n805), .B1(new_n791), .B2(G311), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n971), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n968), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n769), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n770), .B1(new_n404), .B2(new_n216), .C1(new_n232), .C2(new_n762), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n960), .A2(new_n756), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n729), .B1(new_n595), .B2(new_n700), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n660), .A2(new_n691), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n985), .A2(KEYINPUT108), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT108), .B1(new_n985), .B2(new_n986), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n701), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT109), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(KEYINPUT42), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n660), .B1(new_n989), .B2(new_n544), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(new_n691), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT43), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n993), .A2(new_n996), .B1(new_n997), .B2(new_n958), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n958), .A2(new_n997), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n989), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n699), .A2(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT110), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n708), .B(KEYINPUT41), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n703), .A2(new_n989), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT45), .Z(new_n1007));
  NOR2_X1   g0807(.A1(new_n703), .A2(new_n989), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT44), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(new_n699), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n501), .A2(new_n700), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n697), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT111), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT111), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n701), .A3(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n695), .B(new_n1016), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n751), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1011), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1005), .B1(new_n1020), .B2(new_n751), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1021), .A2(new_n754), .B1(new_n1002), .B2(new_n1000), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n984), .B1(new_n1004), .B2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n697), .A2(new_n959), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n761), .B1(new_n229), .B2(new_n291), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n706), .B2(new_n757), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n350), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT50), .B1(new_n350), .B2(G50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n706), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1026), .A2(new_n1030), .B1(new_n512), .B2(new_n707), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n756), .B1(new_n1031), .B2(new_n771), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n800), .A2(G77), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n571), .B2(new_n841), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n306), .B1(new_n796), .B2(new_n256), .C1(new_n202), .C2(new_n808), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G150), .C2(new_n778), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n791), .A2(G159), .B1(new_n650), .B2(new_n785), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n350), .C2(new_n806), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n778), .A2(G326), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n306), .B1(new_n803), .B2(G116), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n784), .A2(new_n969), .B1(new_n801), .B2(new_n843), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n805), .A2(G311), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G303), .A2(new_n795), .B1(new_n798), .B2(G317), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n792), .C2(new_n809), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1039), .B(new_n1040), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1038), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1032), .B1(new_n1051), .B2(new_n769), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1017), .A2(new_n754), .B1(new_n1024), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1018), .A2(new_n708), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1017), .A2(new_n751), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(G393));
  NAND2_X1  g0856(.A1(new_n236), .A2(new_n761), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n770), .C1(new_n571), .C2(new_n216), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT113), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n708), .B(new_n754), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n779), .A2(new_n809), .B1(new_n969), .B2(new_n801), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT115), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n276), .B1(new_n512), .B2(new_n841), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1061), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT116), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n796), .A2(new_n843), .B1(new_n784), .B2(new_n455), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n791), .A2(G317), .B1(G311), .B2(new_n798), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(G303), .C2(new_n805), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n785), .A2(G77), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n350), .B2(new_n796), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n791), .A2(G150), .B1(G159), .B2(new_n798), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G50), .C2(new_n805), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n306), .B1(new_n841), .B2(new_n395), .C1(new_n801), .C2(new_n256), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G143), .B2(new_n778), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT114), .Z(new_n1077));
  AOI22_X1  g0877(.A1(new_n1065), .A2(new_n1069), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n769), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1001), .B2(new_n768), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1011), .B2(new_n754), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1020), .A2(new_n708), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1011), .A2(new_n1019), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(G390));
  NAND3_X1  g0885(.A1(new_n750), .A2(new_n830), .A3(new_n884), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n884), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n914), .A2(new_n700), .A3(new_n830), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n881), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n904), .B1(new_n893), .B2(new_n896), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT117), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT117), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n827), .B1(new_n732), .B2(new_n830), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1090), .C1(new_n1094), .C2(new_n1087), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n885), .A2(new_n903), .B1(new_n902), .B2(new_n905), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1086), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n926), .A2(G330), .A3(new_n830), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1087), .A2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n1097), .C1(new_n1092), .C2(new_n1095), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT118), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n920), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT103), .B1(new_n733), .B2(new_n454), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n649), .B(new_n943), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n882), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1087), .A2(new_n1100), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1086), .B2(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1086), .A2(new_n1109), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n1094), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1104), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1094), .A2(new_n1086), .A3(new_n1109), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1111), .B2(new_n1108), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n921), .A2(new_n1115), .A3(KEYINPUT118), .A4(new_n943), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1117), .A2(KEYINPUT119), .A3(new_n1103), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT119), .B1(new_n1117), .B2(new_n1103), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n708), .B1(new_n1103), .B2(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n276), .B1(new_n796), .B2(new_n571), .C1(new_n455), .C2(new_n808), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n779), .A2(new_n843), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1121), .A2(new_n802), .A3(new_n857), .A4(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1070), .B1(new_n806), .B2(new_n512), .C1(new_n969), .C2(new_n792), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n800), .A2(G150), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT53), .Z(new_n1127));
  AOI22_X1  g0927(.A1(G128), .A2(new_n791), .B1(new_n805), .B2(G137), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n778), .A2(G125), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n795), .B1(new_n798), .B2(G132), .ZN(new_n1132));
  AND4_X1   g0932(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n306), .B1(new_n841), .B2(new_n202), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(KEYINPUT120), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(KEYINPUT120), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n780), .C2(new_n784), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1123), .A2(new_n1125), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n756), .B1(new_n351), .B2(new_n839), .C1(new_n1139), .C2(new_n1079), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n902), .A2(new_n905), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n766), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1103), .B2(new_n754), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1120), .A2(new_n1143), .ZN(G378));
  NAND2_X1  g0944(.A1(new_n646), .A2(new_n432), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n888), .A2(new_n431), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT55), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1145), .B(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  AND4_X1   g0950(.A1(G330), .A2(new_n933), .A3(new_n941), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1150), .B1(new_n946), .B2(G330), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n909), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT122), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1150), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n942), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n946), .A2(G330), .A3(new_n1150), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n908), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n908), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT122), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1155), .A2(new_n767), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G128), .A2(new_n798), .B1(new_n795), .B2(G137), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n801), .B2(new_n1130), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n806), .A2(new_n861), .B1(new_n784), .B2(new_n851), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G125), .C2(new_n791), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n244), .B(new_n290), .C1(new_n841), .C2(new_n780), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G124), .B2(new_n778), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n805), .A2(G97), .B1(G68), .B2(new_n785), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n455), .B2(new_n792), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n306), .A2(G41), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G107), .B2(new_n798), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n1033), .C1(new_n338), .C2(new_n841), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n779), .A2(new_n969), .B1(new_n796), .B2(new_n404), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1175), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1177), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1184));
  AND4_X1   g0984(.A1(new_n1173), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n756), .B1(G50), .B2(new_n839), .C1(new_n1185), .C2(new_n1079), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n1162), .A2(new_n753), .B1(new_n1163), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1117), .A2(new_n1103), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT119), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1117), .A2(new_n1103), .A3(KEYINPUT119), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1107), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1188), .B1(new_n1193), .B2(new_n1162), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1107), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1188), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n709), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1187), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n1087), .A2(new_n766), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n756), .B1(new_n839), .B2(G68), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n276), .B1(new_n808), .B2(new_n969), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G107), .B2(new_n795), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n963), .B1(G97), .B2(new_n800), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n847), .C2(new_n779), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n805), .A2(G116), .B1(new_n650), .B2(new_n785), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n843), .B2(new_n792), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n805), .A2(new_n1131), .B1(G50), .B2(new_n785), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n861), .B2(new_n792), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n306), .B1(new_n808), .B2(new_n852), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G150), .B2(new_n795), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n778), .A2(G128), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n800), .A2(G159), .B1(new_n803), .B2(G58), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1206), .A2(new_n1208), .B1(new_n1210), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1202), .B1(new_n1216), .B2(new_n769), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1115), .A2(new_n754), .B1(new_n1201), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1113), .A2(new_n1116), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1220), .B2(new_n1005), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT123), .Z(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(G387), .ZN(new_n1224));
  INV_X1    g1024(.A(G378), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n1199), .A3(new_n1222), .ZN(G407));
  NOR2_X1   g1028(.A1(new_n679), .A2(G343), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1199), .A2(new_n1225), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G407), .A2(G213), .A3(new_n1230), .ZN(G409));
  AOI21_X1  g1031(.A(new_n753), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1163), .A2(new_n1186), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT125), .Z(new_n1235));
  NOR3_X1   g1035(.A1(new_n1193), .A2(new_n1005), .A3(new_n1162), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1225), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1187), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1238), .A2(KEYINPUT124), .A3(G378), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT124), .B1(new_n1199), .B2(G378), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1237), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1229), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1220), .A2(KEYINPUT60), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1195), .A2(new_n1115), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1246), .B(new_n708), .C1(KEYINPUT60), .C2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G384), .B1(new_n1248), .B2(new_n1218), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(G384), .A3(new_n1218), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(KEYINPUT126), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G2897), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1244), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1251), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(new_n1249), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1258), .A2(KEYINPUT126), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1254), .B1(new_n1258), .B2(KEYINPUT126), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1256), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1245), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1243), .A2(new_n1244), .A3(new_n1258), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G393), .B(G396), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G390), .B(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1224), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1268), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(G387), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1197), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n708), .B1(new_n1193), .B2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1239), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT124), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1240), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1229), .B1(new_n1281), .B2(new_n1237), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(KEYINPUT63), .A3(new_n1258), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1263), .A2(new_n1266), .A3(new_n1273), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1282), .B2(new_n1261), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1264), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1282), .A2(KEYINPUT62), .A3(new_n1258), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1272), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1269), .A2(KEYINPUT127), .A3(new_n1271), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1284), .B1(new_n1290), .B2(new_n1294), .ZN(G405));
  OAI21_X1  g1095(.A(new_n1281), .B1(G378), .B2(new_n1199), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1296), .A2(new_n1258), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1258), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1272), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1272), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(G402));
endmodule


