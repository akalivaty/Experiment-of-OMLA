

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n879) );
  AND2_X1 U553 ( .A1(n532), .A2(n531), .ZN(G160) );
  AND2_X2 U554 ( .A1(n696), .A2(G1996), .ZN(n684) );
  NOR2_X2 U555 ( .A1(n991), .A2(n687), .ZN(n693) );
  NOR2_X2 U556 ( .A1(n527), .A2(G2105), .ZN(n875) );
  BUF_X2 U557 ( .A(n875), .Z(n518) );
  NOR2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  NOR2_X2 U559 ( .A1(n550), .A2(n549), .ZN(n681) );
  NOR2_X4 U560 ( .A1(n794), .A2(n683), .ZN(n696) );
  AND2_X1 U561 ( .A1(G125), .A2(n535), .ZN(n519) );
  NAND2_X1 U562 ( .A1(G8), .A2(n749), .ZN(n520) );
  NOR2_X1 U563 ( .A1(n771), .A2(n738), .ZN(n521) );
  INV_X1 U564 ( .A(KEYINPUT90), .ZN(n700) );
  XNOR2_X1 U565 ( .A(n701), .B(n700), .ZN(n704) );
  INV_X1 U566 ( .A(KEYINPUT28), .ZN(n705) );
  XNOR2_X1 U567 ( .A(KEYINPUT94), .B(KEYINPUT30), .ZN(n717) );
  XNOR2_X1 U568 ( .A(n718), .B(n717), .ZN(n719) );
  AND2_X1 U569 ( .A1(n735), .A2(n734), .ZN(n737) );
  XNOR2_X1 U570 ( .A(KEYINPUT17), .B(n539), .ZN(n526) );
  NOR2_X1 U571 ( .A1(G651), .A2(n627), .ZN(n654) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n646) );
  NOR2_X1 U573 ( .A1(n525), .A2(n519), .ZN(n532) );
  INV_X2 U574 ( .A(G2104), .ZN(n527) );
  NAND2_X1 U575 ( .A1(n875), .A2(G101), .ZN(n522) );
  XNOR2_X1 U576 ( .A(n522), .B(KEYINPUT23), .ZN(n523) );
  XNOR2_X1 U577 ( .A(n523), .B(KEYINPUT66), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n527), .A2(G2105), .ZN(n524) );
  XNOR2_X1 U579 ( .A(n524), .B(KEYINPUT65), .ZN(n546) );
  BUF_X1 U580 ( .A(n546), .Z(n535) );
  INV_X1 U581 ( .A(n526), .ZN(n543) );
  NAND2_X1 U582 ( .A1(G137), .A2(n543), .ZN(n529) );
  NAND2_X1 U583 ( .A1(G113), .A2(n879), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U585 ( .A(n530), .B(KEYINPUT67), .ZN(n531) );
  AND2_X1 U586 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U587 ( .A1(G99), .A2(n518), .ZN(n534) );
  NAND2_X1 U588 ( .A1(G111), .A2(n879), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n535), .A2(G123), .ZN(n536) );
  XOR2_X1 U591 ( .A(KEYINPUT18), .B(n536), .Z(n537) );
  NOR2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT17), .B(n539), .Z(n876) );
  NAND2_X1 U594 ( .A1(n876), .A2(G135), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n947) );
  XNOR2_X1 U596 ( .A(G2096), .B(n947), .ZN(n542) );
  OR2_X1 U597 ( .A1(G2100), .A2(n542), .ZN(G156) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  NAND2_X1 U601 ( .A1(G138), .A2(n543), .ZN(n545) );
  NAND2_X1 U602 ( .A1(G102), .A2(n518), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n545), .A2(n544), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G114), .A2(n879), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G126), .A2(n546), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  BUF_X1 U607 ( .A(n681), .Z(G164) );
  INV_X1 U608 ( .A(G651), .ZN(n555) );
  NOR2_X1 U609 ( .A1(G543), .A2(n555), .ZN(n551) );
  XOR2_X1 U610 ( .A(KEYINPUT1), .B(n551), .Z(n647) );
  NAND2_X1 U611 ( .A1(n647), .A2(G64), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT70), .ZN(n554) );
  XOR2_X1 U613 ( .A(G543), .B(KEYINPUT0), .Z(n627) );
  NAND2_X1 U614 ( .A1(G52), .A2(n654), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n562) );
  NOR2_X1 U616 ( .A1(n627), .A2(n555), .ZN(n650) );
  NAND2_X1 U617 ( .A1(n650), .A2(G77), .ZN(n556) );
  XOR2_X1 U618 ( .A(KEYINPUT71), .B(n556), .Z(n558) );
  NAND2_X1 U619 ( .A1(n646), .A2(G90), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT72), .B(n559), .Z(n560) );
  XNOR2_X1 U622 ( .A(KEYINPUT9), .B(n560), .ZN(n561) );
  NOR2_X1 U623 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U624 ( .A1(n647), .A2(G63), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT77), .B(n563), .Z(n565) );
  NAND2_X1 U626 ( .A1(n654), .A2(G51), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U628 ( .A(KEYINPUT6), .B(n566), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n646), .A2(G89), .ZN(n567) );
  XNOR2_X1 U630 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U631 ( .A1(G76), .A2(n650), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT5), .B(n570), .Z(n571) );
  XNOR2_X1 U634 ( .A(KEYINPUT76), .B(n571), .ZN(n572) );
  NOR2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT7), .B(n574), .Z(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT78), .B(n575), .ZN(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U641 ( .A(G223), .B(KEYINPUT73), .ZN(n830) );
  NAND2_X1 U642 ( .A1(n830), .A2(G567), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  XOR2_X1 U644 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n579) );
  NAND2_X1 U645 ( .A1(G56), .A2(n647), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(n586) );
  XNOR2_X1 U647 ( .A(KEYINPUT75), .B(KEYINPUT13), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n646), .A2(G81), .ZN(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT12), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G68), .A2(n650), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n654), .A2(G43), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n991) );
  INV_X1 U656 ( .A(G860), .ZN(n614) );
  OR2_X1 U657 ( .A1(n991), .A2(n614), .ZN(G153) );
  INV_X1 U658 ( .A(G171), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U660 ( .A1(G92), .A2(n646), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G66), .A2(n647), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G79), .A2(n650), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G54), .A2(n654), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U667 ( .A(KEYINPUT15), .B(n595), .Z(n990) );
  OR2_X1 U668 ( .A1(n990), .A2(G868), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(G284) );
  NAND2_X1 U670 ( .A1(G53), .A2(n654), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G65), .A2(n647), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G91), .A2(n646), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G78), .A2(n650), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n982) );
  INV_X1 U677 ( .A(n982), .ZN(G299) );
  XNOR2_X1 U678 ( .A(KEYINPUT79), .B(G868), .ZN(n604) );
  NOR2_X1 U679 ( .A1(G286), .A2(n604), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n614), .A2(G559), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n607), .A2(n990), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n991), .ZN(n609) );
  XNOR2_X1 U686 ( .A(KEYINPUT80), .B(n609), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G868), .A2(n990), .ZN(n610) );
  NOR2_X1 U688 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G559), .A2(n990), .ZN(n613) );
  XOR2_X1 U691 ( .A(n991), .B(n613), .Z(n662) );
  NAND2_X1 U692 ( .A1(n614), .A2(n662), .ZN(n623) );
  NAND2_X1 U693 ( .A1(G67), .A2(n647), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n615), .B(KEYINPUT82), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G93), .A2(n646), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G55), .A2(n654), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G80), .A2(n650), .ZN(n618) );
  XNOR2_X1 U699 ( .A(KEYINPUT81), .B(n618), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n664) );
  XNOR2_X1 U702 ( .A(n623), .B(n664), .ZN(G145) );
  NAND2_X1 U703 ( .A1(G49), .A2(n654), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n647), .A2(n626), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G75), .A2(n650), .ZN(n630) );
  XOR2_X1 U710 ( .A(KEYINPUT84), .B(n630), .Z(n635) );
  NAND2_X1 U711 ( .A1(G50), .A2(n654), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G62), .A2(n647), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U714 ( .A(KEYINPUT83), .B(n633), .Z(n634) );
  NOR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n646), .A2(G88), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(G303) );
  INV_X1 U718 ( .A(G303), .ZN(G166) );
  NAND2_X1 U719 ( .A1(n647), .A2(G60), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n638), .B(KEYINPUT68), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G85), .A2(n646), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G72), .A2(n650), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G47), .A2(n654), .ZN(n641) );
  XNOR2_X1 U725 ( .A(KEYINPUT69), .B(n641), .ZN(n642) );
  NOR2_X1 U726 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U728 ( .A1(G86), .A2(n646), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G61), .A2(n647), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n650), .A2(G73), .ZN(n651) );
  XOR2_X1 U732 ( .A(KEYINPUT2), .B(n651), .Z(n652) );
  NOR2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n654), .A2(G48), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(G305) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(G288), .ZN(n661) );
  XNOR2_X1 U737 ( .A(G166), .B(G290), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n657), .B(n664), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n982), .B(n658), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n659), .B(G305), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n661), .B(n660), .ZN(n898) );
  XNOR2_X1 U742 ( .A(n662), .B(n898), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n663), .A2(G868), .ZN(n667) );
  INV_X1 U744 ( .A(G868), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n668) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n671), .A2(G2072), .ZN(n672) );
  XOR2_X1 U752 ( .A(KEYINPUT85), .B(n672), .Z(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U756 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U757 ( .A1(G96), .A2(n675), .ZN(n836) );
  NAND2_X1 U758 ( .A1(n836), .A2(G2106), .ZN(n679) );
  NAND2_X1 U759 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U760 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G108), .A2(n677), .ZN(n837) );
  NAND2_X1 U762 ( .A1(n837), .A2(G567), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n679), .A2(n678), .ZN(n856) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n856), .A2(n680), .ZN(n835) );
  NAND2_X1 U766 ( .A1(n835), .A2(G36), .ZN(G176) );
  XNOR2_X1 U767 ( .A(G1981), .B(G305), .ZN(n978) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n794) );
  NOR2_X1 U769 ( .A1(G1384), .A2(n681), .ZN(n682) );
  XNOR2_X1 U770 ( .A(n682), .B(KEYINPUT64), .ZN(n795) );
  INV_X1 U771 ( .A(n795), .ZN(n683) );
  XOR2_X1 U772 ( .A(n684), .B(KEYINPUT26), .Z(n686) );
  INV_X1 U773 ( .A(n696), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n727), .A2(G1341), .ZN(n685) );
  NAND2_X1 U775 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U776 ( .A1(n990), .A2(n693), .ZN(n692) );
  AND2_X1 U777 ( .A1(n727), .A2(G1348), .ZN(n688) );
  XNOR2_X1 U778 ( .A(n688), .B(KEYINPUT91), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n696), .A2(G2067), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n695) );
  OR2_X1 U782 ( .A1(n990), .A2(n693), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n703) );
  NAND2_X1 U784 ( .A1(n696), .A2(G2072), .ZN(n697) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(n697), .Z(n699) );
  NAND2_X1 U786 ( .A1(G1956), .A2(n727), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n982), .A2(n704), .ZN(n702) );
  NAND2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U790 ( .A1(n982), .A2(n704), .ZN(n706) );
  XNOR2_X1 U791 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U792 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U793 ( .A(KEYINPUT29), .B(KEYINPUT92), .ZN(n709) );
  XNOR2_X1 U794 ( .A(n710), .B(n709), .ZN(n714) );
  XNOR2_X1 U795 ( .A(KEYINPUT25), .B(G2078), .ZN(n1008) );
  NOR2_X1 U796 ( .A1(n727), .A2(n1008), .ZN(n712) );
  AND2_X1 U797 ( .A1(n727), .A2(G1961), .ZN(n711) );
  NOR2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n720) );
  AND2_X1 U799 ( .A1(G171), .A2(n720), .ZN(n713) );
  NOR2_X2 U800 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U801 ( .A(n715), .B(KEYINPUT93), .ZN(n725) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n727), .ZN(n749) );
  NAND2_X1 U803 ( .A1(G8), .A2(n727), .ZN(n771) );
  NOR2_X1 U804 ( .A1(G1966), .A2(n771), .ZN(n746) );
  NOR2_X1 U805 ( .A1(n749), .A2(n746), .ZN(n716) );
  NAND2_X1 U806 ( .A1(G8), .A2(n716), .ZN(n718) );
  NOR2_X1 U807 ( .A1(G168), .A2(n719), .ZN(n722) );
  NOR2_X1 U808 ( .A1(G171), .A2(n720), .ZN(n721) );
  NOR2_X1 U809 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U810 ( .A(KEYINPUT31), .B(n723), .Z(n724) );
  NAND2_X1 U811 ( .A1(n725), .A2(n724), .ZN(n744) );
  AND2_X1 U812 ( .A1(G286), .A2(G8), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n744), .A2(n726), .ZN(n735) );
  INV_X1 U814 ( .A(G8), .ZN(n733) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n771), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U818 ( .A(n730), .B(KEYINPUT96), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n731), .A2(G303), .ZN(n732) );
  OR2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U821 ( .A(KEYINPUT97), .B(KEYINPUT32), .Z(n736) );
  XNOR2_X1 U822 ( .A(n737), .B(n736), .ZN(n764) );
  NAND2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n985) );
  INV_X1 U824 ( .A(n985), .ZN(n738) );
  OR2_X1 U825 ( .A1(KEYINPUT33), .A2(n521), .ZN(n742) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NAND2_X1 U827 ( .A1(KEYINPUT33), .A2(n753), .ZN(n739) );
  NOR2_X1 U828 ( .A1(n771), .A2(n739), .ZN(n740) );
  XOR2_X1 U829 ( .A(n740), .B(KEYINPUT98), .Z(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n756) );
  INV_X1 U831 ( .A(n756), .ZN(n743) );
  AND2_X1 U832 ( .A1(n764), .A2(n743), .ZN(n751) );
  INV_X1 U833 ( .A(n744), .ZN(n745) );
  NOR2_X1 U834 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U835 ( .A(KEYINPUT95), .B(n747), .ZN(n748) );
  INV_X1 U836 ( .A(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n750), .A2(n520), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n751), .A2(n765), .ZN(n758) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n986) );
  INV_X1 U841 ( .A(KEYINPUT33), .ZN(n754) );
  AND2_X1 U842 ( .A1(n986), .A2(n754), .ZN(n755) );
  OR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U845 ( .A(n759), .B(KEYINPUT99), .ZN(n760) );
  NOR2_X1 U846 ( .A1(n978), .A2(n760), .ZN(n761) );
  XNOR2_X1 U847 ( .A(n761), .B(KEYINPUT100), .ZN(n775) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n762) );
  XOR2_X1 U849 ( .A(KEYINPUT101), .B(n762), .Z(n763) );
  NAND2_X1 U850 ( .A1(G8), .A2(n763), .ZN(n767) );
  NAND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n768), .A2(n771), .ZN(n773) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U855 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  OR2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U858 ( .A1(n775), .A2(n774), .ZN(n808) );
  NAND2_X1 U859 ( .A1(G117), .A2(n879), .ZN(n777) );
  NAND2_X1 U860 ( .A1(G129), .A2(n535), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U862 ( .A1(n518), .A2(G105), .ZN(n778) );
  XOR2_X1 U863 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U865 ( .A1(n876), .A2(G141), .ZN(n781) );
  NAND2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n887) );
  NAND2_X1 U867 ( .A1(G1996), .A2(n887), .ZN(n792) );
  NAND2_X1 U868 ( .A1(G131), .A2(n876), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT88), .ZN(n790) );
  NAND2_X1 U870 ( .A1(G95), .A2(n518), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G119), .A2(n535), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G107), .A2(n879), .ZN(n786) );
  XNOR2_X1 U874 ( .A(KEYINPUT87), .B(n786), .ZN(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n864) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n864), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U879 ( .A(KEYINPUT89), .B(n793), .ZN(n953) );
  INV_X1 U880 ( .A(n953), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n824) );
  NAND2_X1 U882 ( .A1(n796), .A2(n824), .ZN(n812) );
  NAND2_X1 U883 ( .A1(n876), .A2(G140), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT86), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G104), .A2(n518), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U887 ( .A(KEYINPUT34), .B(n800), .ZN(n805) );
  NAND2_X1 U888 ( .A1(G116), .A2(n879), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G128), .A2(n535), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U891 ( .A(KEYINPUT35), .B(n803), .Z(n804) );
  NOR2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n806), .ZN(n894) );
  XNOR2_X1 U894 ( .A(G2067), .B(KEYINPUT37), .ZN(n821) );
  NOR2_X1 U895 ( .A1(n894), .A2(n821), .ZN(n955) );
  NAND2_X1 U896 ( .A1(n824), .A2(n955), .ZN(n819) );
  NAND2_X1 U897 ( .A1(n812), .A2(n819), .ZN(n807) );
  NOR2_X2 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U899 ( .A(n809), .B(KEYINPUT102), .ZN(n811) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U901 ( .A1(n824), .A2(n993), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n827) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n887), .ZN(n957) );
  INV_X1 U904 ( .A(n812), .ZN(n816) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n864), .ZN(n949) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n813) );
  XOR2_X1 U907 ( .A(n813), .B(KEYINPUT103), .Z(n814) );
  NOR2_X1 U908 ( .A1(n949), .A2(n814), .ZN(n815) );
  NOR2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n957), .A2(n817), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n894), .A2(n821), .ZN(n963) );
  NAND2_X1 U914 ( .A1(n822), .A2(n963), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U916 ( .A(n825), .B(KEYINPUT104), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n827), .A2(n826), .ZN(n829) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n828) );
  XNOR2_X1 U919 ( .A(n829), .B(n828), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n830), .ZN(G217) );
  INV_X1 U921 ( .A(G661), .ZN(n832) );
  NAND2_X1 U922 ( .A1(G2), .A2(G15), .ZN(n831) );
  NOR2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U924 ( .A(KEYINPUT108), .B(n833), .Z(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XOR2_X1 U933 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U934 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U939 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U940 ( .A(G2084), .B(G2078), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(G227) );
  XNOR2_X1 U942 ( .A(G1991), .B(KEYINPUT110), .ZN(n855) );
  XOR2_X1 U943 ( .A(G1981), .B(G1996), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1961), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1956), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(G229) );
  INV_X1 U953 ( .A(n856), .ZN(G319) );
  NAND2_X1 U954 ( .A1(G100), .A2(n518), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G112), .A2(n879), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U957 ( .A1(G124), .A2(n535), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n876), .A2(G136), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U961 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U962 ( .A(G162), .B(n864), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n865), .B(n947), .ZN(n874) );
  NAND2_X1 U964 ( .A1(G118), .A2(n879), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G130), .A2(n535), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U967 ( .A1(G106), .A2(n518), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G142), .A2(n876), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(KEYINPUT45), .B(n870), .Z(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n886) );
  NAND2_X1 U973 ( .A1(G103), .A2(n518), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G139), .A2(n876), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U976 ( .A1(G115), .A2(n879), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G127), .A2(n535), .ZN(n880) );
  NAND2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n966) );
  XNOR2_X1 U981 ( .A(G164), .B(n966), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n896) );
  XNOR2_X1 U983 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n887), .B(KEYINPUT111), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U986 ( .A(n890), .B(KEYINPUT48), .Z(n892) );
  XNOR2_X1 U987 ( .A(G160), .B(KEYINPUT46), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U989 ( .A(n894), .B(n893), .Z(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U991 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n991), .B(n898), .ZN(n900) );
  XNOR2_X1 U993 ( .A(G171), .B(n990), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(G286), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G397) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n917) );
  XNOR2_X1 U1000 ( .A(G2443), .B(G2427), .ZN(n914) );
  XOR2_X1 U1001 ( .A(G2430), .B(KEYINPUT107), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2454), .B(G2435), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1004 ( .A(G2438), .B(KEYINPUT106), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2446), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n915), .A2(G14), .ZN(n920) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n920), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G19), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(G6), .B(G1981), .ZN(n921) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1022 ( .A(KEYINPUT125), .B(n923), .Z(n927) );
  XNOR2_X1 U1023 ( .A(KEYINPUT59), .B(KEYINPUT126), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n924), .B(G4), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G1348), .B(n925), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(G20), .B(G1956), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(KEYINPUT60), .B(n930), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(G1966), .B(G21), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(G5), .B(G1961), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(G1986), .B(G24), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(G1971), .B(G22), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G1976), .B(KEYINPUT127), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(n937), .B(G23), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT58), .B(n940), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT61), .B(n943), .ZN(n945) );
  INV_X1 U1043 ( .A(G16), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n946), .A2(G11), .ZN(n1005) );
  XNOR2_X1 U1046 ( .A(G160), .B(G2084), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1049 ( .A(KEYINPUT115), .B(n951), .Z(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n961) );
  XOR2_X1 U1052 ( .A(G2090), .B(G162), .Z(n956) );
  XNOR2_X1 U1053 ( .A(KEYINPUT116), .B(n956), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(KEYINPUT51), .B(n959), .Z(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(KEYINPUT117), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT118), .B(n965), .ZN(n971) );
  XOR2_X1 U1060 ( .A(G2072), .B(n966), .Z(n968) );
  XOR2_X1 U1061 ( .A(G164), .B(G2078), .Z(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT50), .B(n969), .Z(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT52), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n1023) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n1023), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n974), .B(KEYINPUT120), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(G29), .ZN(n1003) );
  XOR2_X1 U1070 ( .A(G16), .B(KEYINPUT56), .Z(n976) );
  XNOR2_X1 U1071 ( .A(KEYINPUT123), .B(n976), .ZN(n1001) );
  XNOR2_X1 U1072 ( .A(G301), .B(G1961), .ZN(n981) );
  XOR2_X1 U1073 ( .A(G1966), .B(G168), .Z(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(KEYINPUT57), .B(n979), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n999) );
  XNOR2_X1 U1077 ( .A(n982), .B(G1956), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(G1971), .A2(G303), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1082 ( .A(KEYINPUT124), .B(n989), .Z(n997) );
  XNOR2_X1 U1083 ( .A(G1348), .B(n990), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(G1341), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1028) );
  XNOR2_X1 U1092 ( .A(KEYINPUT121), .B(G2067), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1006), .B(G26), .ZN(n1016) );
  XOR2_X1 U1094 ( .A(G2072), .B(G33), .Z(n1007) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(G28), .ZN(n1014) );
  XNOR2_X1 U1096 ( .A(G27), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1996), .B(G32), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1991), .B(G25), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1017), .B(KEYINPUT53), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(G2084), .B(G34), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT54), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G35), .B(G2090), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(n1023), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT122), .B(n1026), .Z(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

