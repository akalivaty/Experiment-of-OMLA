//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT73), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(G110), .B(G140), .Z(new_n196));
  XNOR2_X1  g010(.A(new_n195), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G104), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G107), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  OAI22_X1  g017(.A1(new_n201), .A2(G107), .B1(KEYINPUT86), .B2(KEYINPUT3), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT87), .B1(new_n199), .B2(G104), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT87), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n201), .A3(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n200), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n203), .B1(new_n212), .B2(new_n198), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT66), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT66), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G143), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT66), .A2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT66), .A2(G146), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n218), .B1(new_n225), .B2(G143), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n220), .B1(new_n229), .B2(KEYINPUT1), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n222), .B(KEYINPUT90), .C1(new_n226), .C2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT90), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n216), .A2(new_n232), .A3(new_n219), .A4(new_n221), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n213), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT68), .A2(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT68), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n214), .A2(new_n215), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n228), .B1(new_n241), .B2(new_n227), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n222), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n213), .A2(KEYINPUT10), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n201), .A2(G107), .ZN(new_n246));
  INV_X1    g060(.A(new_n210), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(new_n205), .A3(new_n207), .A4(new_n204), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(G101), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT0), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n220), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT0), .A3(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT67), .B1(new_n242), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n226), .A2(KEYINPUT0), .A3(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n227), .B1(new_n223), .B2(new_n224), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n229), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n257), .A4(new_n262), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n252), .A2(new_n264), .A3(new_n265), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n251), .B1(new_n212), .B2(new_n198), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n250), .A2(G101), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n272), .A2(KEYINPUT88), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT88), .B1(new_n272), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT89), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n212), .A2(new_n198), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n273), .A3(KEYINPUT4), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n272), .A2(KEYINPUT88), .A3(new_n273), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT89), .A3(new_n271), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n245), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT11), .ZN(new_n287));
  INV_X1    g101(.A(G134), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(G137), .ZN(new_n289));
  INV_X1    g103(.A(G137), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT11), .A3(G134), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(G137), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G131), .ZN(new_n294));
  AOI21_X1  g108(.A(G131), .B1(new_n288), .B2(G137), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n289), .A2(new_n295), .A3(new_n291), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n197), .B1(new_n286), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n298), .B2(new_n286), .ZN(new_n300));
  INV_X1    g114(.A(new_n245), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT89), .B1(new_n284), .B2(new_n271), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n277), .B(new_n270), .C1(new_n282), .C2(new_n283), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n298), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n231), .ZN(new_n306));
  INV_X1    g120(.A(new_n203), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n233), .B(new_n307), .C1(new_n250), .C2(G101), .ZN(new_n308));
  OAI22_X1  g122(.A1(new_n306), .A2(new_n308), .B1(new_n213), .B2(new_n243), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n309), .A2(KEYINPUT91), .A3(KEYINPUT12), .A4(new_n297), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n279), .A2(new_n307), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n237), .A2(new_n238), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n223), .A2(new_n224), .A3(new_n227), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n315), .A2(new_n267), .B1(new_n226), .B2(new_n221), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n298), .B1(new_n317), .B2(new_n234), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n310), .B1(KEYINPUT12), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT91), .B1(new_n318), .B2(KEYINPUT12), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n197), .B1(new_n305), .B2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n300), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G469), .B1(new_n323), .B2(G902), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT92), .B1(new_n319), .B2(new_n320), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n318), .A2(KEYINPUT12), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n309), .A2(KEYINPUT12), .A3(new_n297), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n327), .A3(new_n330), .A4(new_n310), .ZN(new_n331));
  INV_X1    g145(.A(new_n197), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n325), .A2(new_n331), .A3(new_n304), .A4(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n299), .A2(KEYINPUT93), .A3(new_n331), .A4(new_n325), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n286), .A2(new_n298), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n197), .B1(new_n337), .B2(new_n305), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G469), .ZN(new_n340));
  INV_X1    g154(.A(G902), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n189), .B1(new_n324), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n201), .ZN(new_n345));
  INV_X1    g159(.A(G237), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n194), .A2(G143), .A3(G214), .A4(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n191), .A2(new_n193), .A3(G214), .A4(new_n346), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n227), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT95), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT18), .A3(G131), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n225), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n355), .A2(KEYINPUT79), .A3(G140), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n353), .B2(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G146), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n350), .A2(new_n352), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G131), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n347), .B2(new_n349), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n351), .A3(KEYINPUT18), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT16), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n366));
  INV_X1    g180(.A(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G125), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n365), .A2(new_n366), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT80), .B1(new_n357), .B2(new_n364), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n217), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n365), .A2(new_n366), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n364), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n374), .A2(G146), .A3(new_n371), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n370), .A2(KEYINPUT81), .A3(G146), .A4(new_n371), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n361), .A2(KEYINPUT17), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n347), .A2(new_n349), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G131), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n347), .A2(new_n360), .A3(new_n349), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n381), .B1(new_n385), .B2(KEYINPUT17), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n345), .B(new_n363), .C1(new_n380), .C2(new_n386), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n353), .A2(KEYINPUT19), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT19), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n357), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n383), .A2(new_n384), .B1(new_n225), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n376), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n363), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT96), .ZN(new_n394));
  INV_X1    g208(.A(new_n345), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n391), .A2(new_n376), .B1(new_n359), .B2(new_n362), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT96), .B1(new_n397), .B2(new_n345), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n387), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(G475), .A2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT20), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  INV_X1    g218(.A(new_n386), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n405), .A2(new_n379), .A3(new_n373), .A4(new_n378), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n345), .B1(new_n406), .B2(new_n363), .ZN(new_n407));
  INV_X1    g221(.A(new_n387), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n341), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n402), .A2(new_n404), .B1(G475), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n239), .A2(G143), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n227), .A2(G128), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(G134), .ZN(new_n414));
  XNOR2_X1  g228(.A(G116), .B(G122), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n199), .ZN(new_n416));
  INV_X1    g230(.A(G122), .ZN(new_n417));
  OR3_X1    g231(.A1(new_n417), .A2(KEYINPUT14), .A3(G116), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(G116), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n417), .B2(G116), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n418), .A2(KEYINPUT97), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(G107), .C1(KEYINPUT97), .C2(new_n418), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n414), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n412), .B(KEYINPUT13), .Z(new_n424));
  INV_X1    g238(.A(new_n411), .ZN(new_n425));
  OAI21_X1  g239(.A(G134), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n415), .B(new_n199), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(G134), .C2(new_n413), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n187), .A2(new_n429), .A3(G953), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n423), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n430), .B1(new_n423), .B2(new_n428), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n341), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n410), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n341), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(G898), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n190), .A2(G952), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(G234), .B2(G237), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G116), .B(G119), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT5), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n449));
  INV_X1    g263(.A(G119), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(G116), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n451), .A2(G113), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT2), .B(G113), .Z(new_n453));
  AOI22_X1  g267(.A1(new_n448), .A2(new_n452), .B1(new_n453), .B2(new_n447), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n213), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(G116), .B(G119), .Z(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT2), .B(G113), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n447), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n252), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n455), .B1(new_n284), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n461), .B1(new_n282), .B2(new_n283), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n455), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n469));
  OR3_X1    g283(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n464), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n264), .A2(new_n265), .A3(new_n269), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n316), .A2(new_n355), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n190), .A2(G224), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n464), .B(KEYINPUT8), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n213), .A2(new_n454), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n455), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n475), .B1(KEYINPUT94), .B2(KEYINPUT7), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(KEYINPUT94), .B2(KEYINPUT7), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  AND4_X1   g297(.A1(KEYINPUT7), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n485), .B2(new_n465), .ZN(new_n486));
  OAI21_X1  g300(.A(G210), .B1(G237), .B2(G902), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n477), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n477), .B2(new_n486), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n439), .B(new_n446), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n343), .A2(new_n438), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n450), .A2(G128), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n312), .B2(new_n450), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT24), .B(G110), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n239), .A2(KEYINPUT23), .A3(G119), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n450), .A2(G128), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n500), .B(new_n496), .C1(KEYINPUT23), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n499), .B1(new_n502), .B2(G110), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n380), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n498), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n502), .B2(G110), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n376), .A3(new_n354), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n504), .A2(new_n509), .A3(new_n515), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(G234), .ZN(new_n520));
  OAI21_X1  g334(.A(G217), .B1(new_n520), .B2(G902), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n341), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n526), .A3(new_n341), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n517), .A2(new_n341), .A3(new_n518), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n521), .B1(new_n528), .B2(KEYINPUT25), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n194), .A2(G210), .A3(new_n346), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT27), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT26), .B(G101), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n289), .A2(new_n295), .A3(new_n291), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n290), .A2(G134), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n360), .B1(new_n543), .B2(new_n292), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT69), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT69), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n296), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n541), .B1(new_n549), .B2(new_n316), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n545), .A4(new_n548), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n460), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT72), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n264), .A2(new_n297), .A3(new_n269), .A4(new_n265), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n550), .A2(new_n551), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n243), .A2(new_n296), .A3(new_n546), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n460), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n540), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n549), .A2(new_n316), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n553), .A2(new_n554), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT28), .B1(new_n564), .B2(new_n556), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n539), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(KEYINPUT74), .B(new_n539), .C1(new_n561), .C2(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n550), .A2(KEYINPUT30), .A3(new_n551), .A4(new_n556), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT30), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n559), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n460), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT71), .A4(new_n460), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n557), .A2(new_n538), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT31), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT31), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n582), .B(new_n579), .C1(new_n576), .C2(new_n577), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n570), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n570), .B(KEYINPUT75), .C1(new_n581), .C2(new_n583), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n534), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n588), .A2(KEYINPUT78), .A3(KEYINPUT32), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT78), .B1(new_n588), .B2(KEYINPUT32), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n578), .A2(new_n557), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT76), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n539), .ZN(new_n595));
  INV_X1    g409(.A(new_n557), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n576), .B2(new_n577), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT76), .B1(new_n597), .B2(new_n538), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n561), .A2(new_n565), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT29), .B1(new_n599), .B2(new_n538), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n565), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n538), .A2(KEYINPUT29), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n563), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n557), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT77), .B1(new_n606), .B2(KEYINPUT28), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT77), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n608), .B(new_n540), .C1(new_n605), .C2(new_n557), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n602), .B(new_n603), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n610), .A2(new_n341), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n592), .B1(new_n601), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n578), .A2(new_n580), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n582), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n578), .A2(KEYINPUT31), .A3(new_n580), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT75), .B1(new_n616), .B2(new_n570), .ZN(new_n617));
  INV_X1    g431(.A(new_n587), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n533), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT32), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n612), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n532), .B1(new_n591), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n495), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  AOI21_X1  g438(.A(G902), .B1(new_n586), .B2(new_n587), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n592), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n588), .ZN(new_n627));
  INV_X1    g441(.A(new_n532), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n627), .A2(new_n628), .A3(new_n343), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n409), .A2(G475), .ZN(new_n630));
  INV_X1    g444(.A(new_n404), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n403), .B1(new_n399), .B2(new_n400), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n431), .A2(new_n432), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  OAI22_X1  g451(.A1(new_n431), .A2(new_n432), .B1(KEYINPUT99), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n434), .A2(G902), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT100), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n433), .A2(new_n434), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n636), .A2(new_n643), .A3(new_n638), .A4(new_n639), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n633), .A2(KEYINPUT101), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT101), .B1(new_n633), .B2(new_n645), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n629), .A2(new_n492), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G104), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  NAND2_X1  g467(.A1(new_n477), .A2(new_n486), .ZN(new_n654));
  INV_X1    g468(.A(new_n487), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n488), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n446), .B(KEYINPUT103), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n439), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n436), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n410), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n629), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR3_X1   g480(.A1(new_n510), .A2(KEYINPUT36), .A3(new_n516), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT36), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n504), .A2(new_n509), .B1(new_n668), .B2(new_n515), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n523), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n530), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n626), .A2(new_n588), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n495), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT104), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n675), .B(new_n677), .ZN(G12));
  OAI211_X1 g492(.A(KEYINPUT32), .B(new_n533), .C1(new_n617), .C2(new_n618), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT78), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n619), .A2(new_n620), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n588), .A2(KEYINPUT78), .A3(KEYINPUT32), .ZN(new_n683));
  INV_X1    g497(.A(new_n612), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n682), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n439), .B1(new_n489), .B2(new_n490), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n673), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n444), .B1(new_n440), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n633), .A2(new_n436), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT105), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n685), .A2(new_n343), .A3(new_n687), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XOR2_X1   g507(.A(new_n689), .B(KEYINPUT39), .Z(new_n694));
  AND2_X1   g508(.A1(new_n343), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT40), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n593), .A2(new_n538), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n605), .A2(new_n539), .A3(new_n557), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT106), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI211_X1 g514(.A(KEYINPUT106), .B(new_n699), .C1(new_n597), .C2(new_n539), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n341), .ZN(new_n702));
  OAI21_X1  g516(.A(G472), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(KEYINPUT107), .B(G472), .C1(new_n700), .C2(new_n702), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n705), .B(new_n706), .C1(KEYINPUT32), .C2(new_n588), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n591), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n657), .B(KEYINPUT38), .Z(new_n710));
  INV_X1    g524(.A(new_n439), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n633), .A2(new_n660), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n710), .A2(new_n711), .A3(new_n672), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n695), .A2(new_n696), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n697), .A2(new_n709), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  NAND2_X1  g530(.A1(new_n633), .A2(new_n645), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n689), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n343), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n685), .A2(new_n719), .A3(new_n687), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  OAI21_X1  g535(.A(new_n492), .B1(new_n646), .B2(new_n647), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n339), .A2(new_n341), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n188), .A3(new_n342), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n685), .A2(new_n726), .A3(new_n628), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NOR2_X1   g543(.A1(new_n662), .A2(new_n725), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n685), .A2(new_n730), .A3(new_n628), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT108), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n685), .A2(new_n730), .A3(new_n733), .A4(new_n628), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AOI21_X1  g550(.A(new_n711), .B1(new_n656), .B2(new_n488), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n724), .A2(new_n188), .A3(new_n342), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n438), .A2(new_n672), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n445), .B2(new_n442), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n685), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  OAI21_X1  g557(.A(new_n602), .B1(new_n607), .B2(new_n609), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(new_n539), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n581), .A2(new_n583), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n533), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT109), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n749), .B(new_n533), .C1(new_n745), .C2(new_n746), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n748), .B(new_n750), .C1(new_n625), .C2(new_n592), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n532), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n725), .A2(new_n659), .A3(new_n712), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  OR2_X1    g569(.A1(new_n717), .A2(new_n689), .ZN(new_n756));
  NOR4_X1   g570(.A1(new_n751), .A2(new_n738), .A3(new_n756), .A4(new_n673), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n355), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n657), .A2(new_n711), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n343), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n761), .A2(new_n762), .A3(new_n756), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n619), .A2(KEYINPUT110), .A3(new_n620), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n588), .B2(KEYINPUT32), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n612), .B1(new_n588), .B2(KEYINPUT32), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n628), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT111), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n772), .A3(new_n628), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n764), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n761), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n685), .A2(new_n775), .A3(new_n628), .A4(new_n718), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n762), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n759), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n773), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n772), .B1(new_n769), .B2(new_n628), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n763), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n762), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(KEYINPUT112), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n360), .ZN(G33));
  AND4_X1   g599(.A1(new_n685), .A2(new_n775), .A3(new_n628), .A4(new_n691), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n288), .ZN(G36));
  NAND2_X1  g601(.A1(new_n410), .A2(new_n645), .ZN(new_n788));
  OR2_X1    g602(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n789));
  NAND2_X1  g603(.A1(KEYINPUT113), .A2(KEYINPUT43), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n788), .B2(new_n790), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n627), .A2(new_n673), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n300), .A2(new_n322), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n340), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  NAND2_X1  g620(.A1(G469), .A2(G902), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(KEYINPUT46), .A3(new_n807), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n342), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n188), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n814), .A2(new_n694), .A3(new_n760), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n801), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT115), .B(G137), .Z(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(G39));
  NAND3_X1  g632(.A1(new_n718), .A2(new_n532), .A3(new_n760), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n685), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n814), .A2(KEYINPUT47), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n367), .ZN(G42));
  NOR4_X1   g639(.A1(new_n532), .A2(new_n189), .A3(new_n788), .A4(new_n711), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n710), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n724), .A2(new_n342), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT49), .ZN(new_n832));
  OR4_X1    g646(.A1(new_n709), .A2(new_n828), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n834));
  INV_X1    g648(.A(new_n687), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n591), .B2(new_n621), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n691), .A2(new_n343), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n757), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n672), .A2(new_n689), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n712), .A2(new_n686), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n343), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n681), .A2(new_n683), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(new_n843), .B2(new_n707), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n838), .A2(new_n839), .A3(new_n720), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n751), .A2(new_n673), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n718), .A3(new_n739), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n692), .A2(new_n720), .A3(new_n847), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n692), .A2(new_n847), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n740), .A2(new_n689), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n685), .A2(new_n856), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n751), .A2(new_n673), .A3(new_n756), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n761), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n786), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n659), .B1(new_n717), .B2(new_n661), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n627), .A2(new_n628), .A3(new_n343), .A4(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n727), .A2(new_n742), .A3(new_n754), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n495), .B1(new_n622), .B2(new_n674), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n860), .A2(new_n863), .A3(new_n735), .A4(new_n864), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n784), .A2(new_n850), .A3(new_n855), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n850), .A2(new_n865), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n778), .A2(new_n783), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n834), .B(KEYINPUT54), .C1(new_n866), .C2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n863), .A2(new_n735), .A3(new_n864), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n860), .A3(new_n849), .A4(new_n845), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n853), .B1(new_n872), .B2(new_n784), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n852), .B(KEYINPUT53), .C1(new_n774), .C2(new_n777), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n850), .A2(new_n865), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n867), .A2(new_n868), .A3(new_n854), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n834), .B1(new_n881), .B2(KEYINPUT54), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n792), .A2(new_n445), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n752), .ZN(new_n884));
  INV_X1    g698(.A(new_n725), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n710), .A3(new_n711), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT50), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(KEYINPUT50), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n821), .B(new_n823), .C1(new_n188), .C2(new_n831), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n884), .A2(new_n711), .A3(new_n657), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n888), .A2(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n725), .A2(new_n711), .A3(new_n657), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n532), .A2(new_n445), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n708), .A2(new_n591), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT119), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n633), .A2(new_n645), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n883), .A2(new_n893), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT118), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n846), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n892), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n892), .A2(new_n899), .A3(KEYINPUT51), .A4(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n771), .A2(new_n773), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(KEYINPUT121), .A2(KEYINPUT48), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(new_n649), .B2(new_n896), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n884), .A2(new_n738), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n443), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g728(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n901), .A2(new_n907), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n905), .A2(new_n906), .A3(new_n910), .A4(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n879), .A2(new_n882), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(G952), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n190), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT122), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n833), .B1(new_n919), .B2(new_n922), .ZN(G75));
  INV_X1    g737(.A(new_n194), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n920), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT123), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n873), .A2(new_n876), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(G902), .ZN(new_n930));
  INV_X1    g744(.A(G210), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n469), .A2(new_n470), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n476), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n935), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n928), .B(new_n937), .C1(new_n930), .C2(new_n931), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n927), .B1(new_n936), .B2(new_n938), .ZN(G51));
  XOR2_X1   g753(.A(new_n807), .B(KEYINPUT57), .Z(new_n940));
  NOR3_X1   g754(.A1(new_n869), .A2(KEYINPUT54), .A3(new_n875), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n877), .B1(new_n873), .B2(new_n876), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n339), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n930), .A2(new_n806), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n927), .B1(new_n944), .B2(new_n945), .ZN(G54));
  INV_X1    g760(.A(new_n399), .ZN(new_n947));
  NAND2_X1  g761(.A1(KEYINPUT58), .A2(G475), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n930), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n926), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n930), .A2(new_n947), .A3(new_n948), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(G60));
  NAND2_X1  g766(.A1(new_n636), .A2(new_n638), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n941), .B2(new_n942), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n926), .ZN(new_n958));
  INV_X1    g772(.A(new_n955), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n879), .B2(new_n882), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n960), .B2(new_n953), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n929), .A2(new_n670), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n873), .B2(new_n876), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n965), .B(new_n926), .C1(new_n519), .C2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n966), .A2(new_n519), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n970), .A2(KEYINPUT61), .A3(new_n926), .A4(new_n965), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(G66));
  INV_X1    g786(.A(G224), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n441), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n871), .B2(new_n924), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n194), .A2(G898), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n469), .B2(new_n470), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(G69));
  NAND2_X1  g797(.A1(new_n571), .A2(new_n573), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(new_n390), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(G900), .B2(new_n924), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n907), .A2(new_n694), .A3(new_n814), .A4(new_n841), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n838), .A2(new_n720), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n824), .A2(new_n786), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n816), .A2(new_n868), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n990), .B2(new_n924), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n992));
  INV_X1    g806(.A(new_n985), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n838), .A2(new_n715), .A3(new_n720), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n661), .A2(new_n717), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n695), .A2(new_n760), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n824), .B1(new_n622), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n996), .A2(new_n816), .A3(new_n997), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n993), .B1(new_n1001), .B2(new_n194), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1003));
  OR3_X1    g817(.A1(new_n992), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n992), .B2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  INV_X1    g822(.A(new_n871), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1001), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(new_n538), .A3(new_n593), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1008), .B1(new_n990), .B2(new_n1009), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n593), .A2(new_n538), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n927), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n595), .A2(new_n613), .A3(new_n598), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n881), .A2(new_n1008), .A3(new_n1015), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1011), .A2(new_n1014), .A3(new_n1016), .ZN(G57));
endmodule


