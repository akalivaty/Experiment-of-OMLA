//Secret key is'1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_c1355" written by ABC on Thu Dec 14 03:36:57 2023

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138, new_n139, new_n140, new_n141, new_n142, new_n143, new_n144,
    new_n145, new_n146, new_n147, new_n148, new_n149, new_n150, new_n151,
    new_n152, new_n153, new_n154, new_n155, new_n156, new_n157, new_n158,
    new_n159, new_n160, new_n161, new_n162, new_n163, new_n164, new_n165,
    new_n166, new_n167, new_n168, new_n169, new_n170, new_n171, new_n172,
    new_n173, new_n174, new_n175, new_n176, new_n177, new_n178, new_n179,
    new_n180, new_n181, new_n182, new_n183, new_n184, new_n185, new_n186,
    new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n461,
    new_n462, new_n463, new_n465, new_n466, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n475, new_n476, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n503, new_n504,
    new_n505, new_n507, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n515, new_n516, new_n517, new_n518, new_n520, new_n521, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n625,
    new_n626, new_n628, new_n629, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654;
  OR2_X1    g000(.A1(KEYINPUT8), .A2(G85gat), .ZN(new_n138));
  INV_X1    g001(.A(G92gat), .ZN(new_n139));
  NAND2_X1  g002(.A1(KEYINPUT8), .A2(G85gat), .ZN(new_n140));
  NAND3_X1  g003(.A1(new_n138), .A2(new_n139), .A3(new_n140), .ZN(new_n141));
  NOR2_X1   g004(.A1(KEYINPUT8), .A2(G85gat), .ZN(new_n142));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n143));
  AOI22_X1  g006(.A1(new_n142), .A2(G92gat), .B1(new_n143), .B2(KEYINPUT9), .ZN(new_n144));
  XNOR2_X1  g007(.A(G99gat), .B(G106gat), .ZN(new_n145));
  NAND3_X1  g008(.A1(new_n141), .A2(new_n144), .A3(new_n145), .ZN(new_n146));
  INV_X1    g009(.A(new_n146), .ZN(new_n147));
  AOI21_X1  g010(.A(new_n145), .B1(new_n141), .B2(new_n144), .ZN(new_n148));
  NOR2_X1   g011(.A1(new_n147), .A2(new_n148), .ZN(new_n149));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n150));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n151));
  OR2_X1    g014(.A1(new_n150), .A2(new_n151), .ZN(new_n152));
  NAND2_X1  g015(.A1(new_n150), .A2(new_n151), .ZN(new_n153));
  NAND2_X1  g016(.A1(new_n152), .A2(new_n153), .ZN(new_n154));
  INV_X1    g017(.A(new_n154), .ZN(new_n155));
  NAND2_X1  g018(.A1(new_n149), .A2(new_n155), .ZN(new_n156));
  INV_X1    g019(.A(new_n148), .ZN(new_n157));
  NAND2_X1  g020(.A1(new_n157), .A2(new_n146), .ZN(new_n158));
  NAND2_X1  g021(.A1(new_n158), .A2(new_n154), .ZN(new_n159));
  NAND2_X1  g022(.A1(new_n156), .A2(new_n159), .ZN(new_n160));
  INV_X1    g023(.A(G232gat), .ZN(new_n161));
  INV_X1    g024(.A(G233gat), .ZN(new_n162));
  NOR2_X1   g025(.A1(new_n161), .A2(new_n162), .ZN(new_n163));
  NAND2_X1  g026(.A1(new_n160), .A2(new_n163), .ZN(new_n164));
  INV_X1    g027(.A(new_n164), .ZN(new_n165));
  XOR2_X1   g028(.A(G134gat), .B(G162gat), .Z(new_n166));
  XNOR2_X1  g029(.A(G190gat), .B(G218gat), .ZN(new_n167));
  XNOR2_X1  g030(.A(new_n166), .B(new_n167), .ZN(new_n168));
  XOR2_X1   g031(.A(KEYINPUT34), .B(KEYINPUT35), .Z(new_n169));
  XNOR2_X1  g032(.A(new_n168), .B(new_n169), .ZN(new_n170));
  NOR2_X1   g033(.A1(new_n160), .A2(new_n163), .ZN(new_n171));
  NOR3_X1   g034(.A1(new_n165), .A2(new_n170), .A3(new_n171), .ZN(new_n172));
  INV_X1    g035(.A(KEYINPUT36), .ZN(new_n173));
  OAI21_X1  g036(.A(new_n173), .B1(new_n160), .B2(new_n163), .ZN(new_n174));
  INV_X1    g037(.A(new_n163), .ZN(new_n175));
  NAND4_X1  g038(.A1(new_n156), .A2(new_n159), .A3(KEYINPUT36), .A4(new_n175), .ZN(new_n176));
  NAND3_X1  g039(.A1(new_n174), .A2(new_n164), .A3(new_n176), .ZN(new_n177));
  NAND2_X1  g040(.A1(new_n177), .A2(new_n170), .ZN(new_n178));
  NAND2_X1  g041(.A1(new_n178), .A2(KEYINPUT37), .ZN(new_n179));
  INV_X1    g042(.A(KEYINPUT37), .ZN(new_n180));
  NAND3_X1  g043(.A1(new_n177), .A2(new_n180), .A3(new_n170), .ZN(new_n181));
  AOI21_X1  g044(.A(new_n172), .B1(new_n179), .B2(new_n181), .ZN(new_n182));
  XNOR2_X1  g045(.A(G1gat), .B(G8gat), .ZN(new_n183));
  INV_X1    g046(.A(G15gat), .ZN(new_n184));
  INV_X1    g047(.A(G22gat), .ZN(new_n185));
  NAND2_X1  g048(.A1(new_n184), .A2(new_n185), .ZN(new_n186));
  AOI21_X1  g049(.A(KEYINPUT14), .B1(G15gat), .B2(G22gat), .ZN(new_n187));
  AND3_X1   g050(.A1(KEYINPUT14), .A2(G15gat), .A3(G22gat), .ZN(new_n188));
  OAI211_X1 g051(.A(new_n183), .B(new_n186), .C1(new_n187), .C2(new_n188), .ZN(new_n189));
  INV_X1    g052(.A(KEYINPUT15), .ZN(new_n190));
  OAI21_X1  g053(.A(new_n190), .B1(new_n188), .B2(new_n187), .ZN(new_n191));
  NAND2_X1  g054(.A1(G15gat), .A2(G22gat), .ZN(new_n192));
  INV_X1    g055(.A(KEYINPUT14), .ZN(new_n193));
  NAND2_X1  g056(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g057(.A1(KEYINPUT14), .A2(G15gat), .A3(G22gat), .ZN(new_n195));
  NAND3_X1  g058(.A1(new_n194), .A2(KEYINPUT15), .A3(new_n195), .ZN(new_n196));
  NAND3_X1  g059(.A1(new_n191), .A2(new_n196), .A3(new_n186), .ZN(new_n197));
  INV_X1    g060(.A(new_n183), .ZN(new_n198));
  AND3_X1   g061(.A1(new_n197), .A2(KEYINPUT16), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g062(.A(KEYINPUT16), .B1(new_n197), .B2(new_n198), .ZN(new_n200));
  OAI21_X1  g063(.A(new_n189), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  XOR2_X1   g064(.A(G57gat), .B(G64gat), .Z(new_n202));
  XOR2_X1   g065(.A(G71gat), .B(G78gat), .Z(new_n203));
  XNOR2_X1  g066(.A(new_n202), .B(new_n203), .ZN(new_n204));
  OR2_X1    g067(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g068(.A1(new_n201), .A2(new_n204), .ZN(new_n206));
  NAND3_X1  g069(.A1(new_n205), .A2(KEYINPUT20), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g070(.A(G127gat), .B(G155gat), .ZN(new_n208));
  XNOR2_X1  g071(.A(new_n208), .B(KEYINPUT19), .ZN(new_n209));
  INV_X1    g072(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g073(.A1(G231gat), .A2(G233gat), .ZN(new_n211));
  AND3_X1   g074(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g075(.A(new_n210), .B1(new_n207), .B2(new_n211), .ZN(new_n213));
  NOR2_X1   g076(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g077(.A(G183gat), .B(G211gat), .ZN(new_n215));
  INV_X1    g078(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g079(.A1(new_n205), .A2(new_n206), .ZN(new_n217));
  INV_X1    g080(.A(KEYINPUT20), .ZN(new_n218));
  AOI21_X1  g081(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g082(.A(KEYINPUT20), .B(new_n215), .C1(new_n205), .C2(new_n206), .ZN(new_n220));
  NOR2_X1   g083(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g084(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  OAI22_X1  g085(.A1(new_n212), .A2(new_n213), .B1(new_n220), .B2(new_n219), .ZN(new_n223));
  NAND2_X1  g086(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g087(.A1(G230gat), .A2(G233gat), .ZN(new_n225));
  XOR2_X1   g088(.A(new_n202), .B(new_n203), .Z(new_n226));
  NAND2_X1  g089(.A1(new_n226), .A2(new_n149), .ZN(new_n227));
  NAND2_X1  g090(.A1(new_n158), .A2(new_n204), .ZN(new_n228));
  AOI21_X1  g091(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g092(.A1(new_n229), .A2(KEYINPUT10), .ZN(new_n230));
  NAND3_X1  g093(.A1(new_n227), .A2(new_n228), .A3(new_n225), .ZN(new_n231));
  NAND2_X1  g094(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g095(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT10), .A4(new_n225), .ZN(new_n233));
  NAND2_X1  g096(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g097(.A(G120gat), .B(G148gat), .ZN(new_n235));
  XNOR2_X1  g098(.A(G176gat), .B(G204gat), .ZN(new_n236));
  XOR2_X1   g099(.A(new_n235), .B(new_n236), .Z(new_n237));
  INV_X1    g100(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g101(.A(new_n234), .B(new_n238), .ZN(new_n239));
  INV_X1    g102(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g103(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g104(.A(G169gat), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g105(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g106(.A(new_n243), .B(KEYINPUT11), .ZN(new_n244));
  NAND2_X1  g107(.A1(new_n201), .A2(new_n155), .ZN(new_n245));
  OAI211_X1 g108(.A(new_n154), .B(new_n189), .C1(new_n199), .C2(new_n200), .ZN(new_n246));
  NAND3_X1  g109(.A1(new_n245), .A2(KEYINPUT17), .A3(new_n246), .ZN(new_n247));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n248));
  NAND3_X1  g111(.A1(new_n201), .A2(new_n248), .A3(new_n155), .ZN(new_n249));
  NAND2_X1  g112(.A1(G229gat), .A2(G233gat), .ZN(new_n250));
  XOR2_X1   g113(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  XNOR2_X1  g114(.A(new_n251), .B(KEYINPUT13), .ZN(new_n252));
  NAND3_X1  g115(.A1(new_n247), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g116(.A1(new_n245), .A2(new_n246), .A3(new_n251), .ZN(new_n254));
  AOI21_X1  g117(.A(new_n244), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g118(.A(KEYINPUT18), .ZN(new_n256));
  AND3_X1   g119(.A1(new_n247), .A2(new_n249), .A3(new_n252), .ZN(new_n257));
  NAND2_X1  g120(.A1(new_n254), .A2(new_n244), .ZN(new_n258));
  OAI21_X1  g121(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g122(.A1(new_n254), .A2(new_n244), .ZN(new_n260));
  NAND3_X1  g123(.A1(new_n260), .A2(KEYINPUT18), .A3(new_n253), .ZN(new_n261));
  AOI21_X1  g124(.A(new_n255), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR3_X1   g125(.A1(new_n224), .A2(new_n240), .A3(new_n262), .ZN(new_n263));
  INV_X1    g126(.A(G141gat), .ZN(new_n264));
  INV_X1    g127(.A(G148gat), .ZN(new_n265));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g130(.A1(new_n267), .A2(G141gat), .A3(G148gat), .ZN(new_n268));
  OAI211_X1 g131(.A(new_n266), .B(new_n268), .C1(G141gat), .C2(G148gat), .ZN(new_n269));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n270));
  XNOR2_X1  g133(.A(KEYINPUT4), .B(G155gat), .ZN(new_n271));
  OAI211_X1 g134(.A(new_n269), .B(new_n270), .C1(G162gat), .C2(new_n271), .ZN(new_n272));
  INV_X1    g135(.A(G155gat), .ZN(new_n273));
  INV_X1    g136(.A(G162gat), .ZN(new_n274));
  NAND2_X1  g137(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g138(.A1(new_n275), .A2(new_n270), .B1(G141gat), .B2(G148gat), .ZN(new_n276));
  XNOR2_X1  g139(.A(KEYINPUT2), .B(G148gat), .ZN(new_n277));
  OAI21_X1  g140(.A(new_n276), .B1(G141gat), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g141(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g142(.A(KEYINPUT7), .ZN(new_n280));
  XNOR2_X1  g143(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g144(.A1(KEYINPUT0), .A2(G113gat), .ZN(new_n282));
  NAND3_X1  g145(.A1(new_n282), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n283));
  NAND2_X1  g146(.A1(KEYINPUT1), .A2(G127gat), .ZN(new_n284));
  NAND3_X1  g147(.A1(new_n284), .A2(KEYINPUT0), .A3(G113gat), .ZN(new_n285));
  NAND2_X1  g148(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g149(.A(G120gat), .B1(KEYINPUT0), .B2(G113gat), .ZN(new_n287));
  XNOR2_X1  g150(.A(new_n286), .B(new_n287), .ZN(new_n288));
  OAI21_X1  g151(.A(G134gat), .B1(KEYINPUT1), .B2(G127gat), .ZN(new_n289));
  INV_X1    g152(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g153(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g154(.A(new_n287), .ZN(new_n292));
  XNOR2_X1  g155(.A(new_n286), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g156(.A1(new_n293), .A2(new_n289), .ZN(new_n294));
  NAND2_X1  g157(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n296));
  NAND2_X1  g159(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g160(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g161(.A1(new_n281), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  INV_X1    g163(.A(new_n279), .ZN(new_n301));
  NAND2_X1  g164(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g165(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n304));
  NAND3_X1  g167(.A1(new_n291), .A2(new_n294), .A3(new_n279), .ZN(new_n305));
  NAND3_X1  g168(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g169(.A(new_n300), .ZN(new_n307));
  NAND3_X1  g170(.A1(new_n295), .A2(KEYINPUT5), .A3(new_n301), .ZN(new_n308));
  NAND3_X1  g171(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g172(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n311));
  XNOR2_X1  g174(.A(G57gat), .B(G85gat), .ZN(new_n312));
  XOR2_X1   g175(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g176(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g177(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g178(.A1(new_n303), .A2(new_n309), .A3(new_n313), .ZN(new_n316));
  NAND2_X1  g179(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g180(.A1(G211gat), .A2(G218gat), .ZN(new_n318));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n319));
  NAND2_X1  g182(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g183(.A1(G211gat), .A2(G218gat), .ZN(new_n321));
  NAND3_X1  g184(.A1(KEYINPUT22), .A2(G211gat), .A3(G218gat), .ZN(new_n322));
  NAND3_X1  g185(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g186(.A1(G197gat), .A2(G204gat), .ZN(new_n324));
  XOR2_X1   g187(.A(KEYINPUT21), .B(G204gat), .Z(new_n325));
  INV_X1    g188(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g189(.A(new_n323), .B(new_n324), .C1(new_n326), .C2(G197gat), .ZN(new_n327));
  AND2_X1   g190(.A1(G197gat), .A2(G204gat), .ZN(new_n328));
  NOR2_X1   g191(.A1(G197gat), .A2(G204gat), .ZN(new_n329));
  OAI211_X1 g192(.A(new_n321), .B(new_n318), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g193(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n332));
  XNOR2_X1  g195(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XOR2_X1   g196(.A(G64gat), .B(G92gat), .Z(new_n334));
  INV_X1    g197(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g198(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g199(.A(new_n331), .ZN(new_n337));
  NOR2_X1   g200(.A1(new_n337), .A2(new_n332), .ZN(new_n338));
  AOI21_X1  g201(.A(new_n331), .B1(G226gat), .B2(G233gat), .ZN(new_n339));
  OAI21_X1  g202(.A(new_n334), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g203(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g204(.A(G183gat), .B(G190gat), .Z(new_n342));
  AND2_X1   g205(.A1(new_n342), .A2(KEYINPUT23), .ZN(new_n343));
  XNOR2_X1  g206(.A(G169gat), .B(G176gat), .ZN(new_n344));
  NOR3_X1   g207(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  OR3_X1    g208(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g209(.A1(new_n342), .A2(new_n344), .ZN(new_n347));
  INV_X1    g210(.A(KEYINPUT24), .ZN(new_n348));
  XNOR2_X1  g211(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g212(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n351));
  XNOR2_X1  g214(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g215(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  INV_X1    g216(.A(new_n351), .ZN(new_n354));
  XNOR2_X1  g217(.A(new_n350), .B(new_n354), .ZN(new_n355));
  NAND3_X1  g218(.A1(new_n355), .A2(new_n340), .A3(new_n336), .ZN(new_n356));
  NAND2_X1  g219(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g220(.A1(new_n317), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g221(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  XNOR2_X1  g222(.A(new_n359), .B(KEYINPUT27), .ZN(new_n360));
  INV_X1    g223(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g224(.A1(new_n281), .A2(new_n331), .ZN(new_n362));
  NOR2_X1   g225(.A1(new_n279), .A2(new_n331), .ZN(new_n363));
  INV_X1    g226(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g227(.A(new_n361), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g228(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g229(.A1(new_n362), .A2(new_n361), .A3(new_n364), .ZN(new_n367));
  NAND2_X1  g230(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g231(.A(KEYINPUT26), .B(G78gat), .ZN(new_n369));
  XNOR2_X1  g232(.A(new_n369), .B(G106gat), .ZN(new_n370));
  XOR2_X1   g233(.A(G22gat), .B(G50gat), .Z(new_n371));
  XNOR2_X1  g234(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n373));
  OAI21_X1  g236(.A(new_n372), .B1(new_n365), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g237(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g238(.A1(new_n366), .A2(new_n367), .A3(new_n373), .A4(new_n372), .ZN(new_n376));
  NAND2_X1  g239(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g240(.A1(new_n358), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g241(.A1(new_n316), .A2(new_n356), .A3(new_n353), .ZN(new_n379));
  AOI21_X1  g242(.A(new_n300), .B1(new_n299), .B2(new_n302), .ZN(new_n380));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n381));
  NOR2_X1   g244(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g245(.A1(new_n306), .A2(new_n308), .ZN(new_n383));
  OAI21_X1  g246(.A(new_n382), .B1(new_n307), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g247(.A(new_n313), .B1(new_n380), .B2(new_n381), .ZN(new_n385));
  AOI21_X1  g248(.A(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g249(.A1(new_n353), .A2(KEYINPUT25), .A3(new_n356), .ZN(new_n387));
  AOI21_X1  g250(.A(KEYINPUT25), .B1(new_n353), .B2(new_n356), .ZN(new_n388));
  NOR2_X1   g251(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g252(.A1(new_n389), .A2(new_n317), .ZN(new_n390));
  OAI22_X1  g253(.A1(new_n378), .A2(new_n386), .B1(new_n390), .B2(new_n377), .ZN(new_n391));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g255(.A1(new_n297), .A2(new_n298), .ZN(new_n393));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n394));
  XOR2_X1   g257(.A(new_n394), .B(KEYINPUT31), .Z(new_n395));
  INV_X1    g258(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g259(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g260(.A(new_n350), .ZN(new_n398));
  NAND3_X1  g261(.A1(new_n297), .A2(new_n298), .A3(new_n395), .ZN(new_n399));
  NAND3_X1  g262(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g263(.A1(new_n400), .A2(KEYINPUT30), .ZN(new_n401));
  AOI21_X1  g264(.A(new_n398), .B1(new_n397), .B2(new_n399), .ZN(new_n402));
  OAI21_X1  g265(.A(G99gat), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g267(.A(new_n404), .B(KEYINPUT29), .ZN(new_n405));
  XNOR2_X1  g268(.A(new_n405), .B(G71gat), .ZN(new_n406));
  NAND2_X1  g269(.A1(new_n397), .A2(new_n399), .ZN(new_n407));
  NAND2_X1  g270(.A1(new_n407), .A2(new_n350), .ZN(new_n408));
  INV_X1    g271(.A(G99gat), .ZN(new_n409));
  NAND4_X1  g272(.A1(new_n408), .A2(KEYINPUT30), .A3(new_n400), .A4(new_n409), .ZN(new_n410));
  NAND3_X1  g273(.A1(new_n403), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  INV_X1    g274(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g275(.A(new_n406), .B1(new_n403), .B2(new_n410), .ZN(new_n413));
  OAI21_X1  g276(.A(new_n392), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g277(.A1(new_n403), .A2(new_n410), .ZN(new_n415));
  INV_X1    g278(.A(new_n406), .ZN(new_n416));
  NAND2_X1  g279(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g280(.A1(new_n417), .A2(KEYINPUT32), .A3(new_n411), .ZN(new_n418));
  AOI21_X1  g281(.A(new_n391), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  INV_X1    g282(.A(new_n377), .ZN(new_n420));
  AOI21_X1  g283(.A(new_n420), .B1(new_n417), .B2(new_n411), .ZN(new_n421));
  NAND2_X1  g284(.A1(new_n421), .A2(new_n390), .ZN(new_n422));
  INV_X1    g285(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g286(.A(new_n182), .B(new_n263), .C1(new_n419), .C2(new_n423), .ZN(new_n424));
  INV_X1    g287(.A(new_n317), .ZN(new_n425));
  OAI21_X1  g288(.A(G1gat), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g289(.A(new_n426), .B(KEYINPUT38), .ZN(new_n427));
  INV_X1    g290(.A(KEYINPUT39), .ZN(new_n428));
  NOR2_X1   g291(.A1(new_n419), .A2(new_n423), .ZN(new_n429));
  INV_X1    g292(.A(new_n172), .ZN(new_n430));
  AND3_X1   g293(.A1(new_n177), .A2(new_n180), .A3(new_n170), .ZN(new_n431));
  AOI21_X1  g294(.A(new_n180), .B1(new_n177), .B2(new_n170), .ZN(new_n432));
  OAI21_X1  g295(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g296(.A1(new_n224), .A2(new_n433), .A3(new_n262), .ZN(new_n434));
  INV_X1    g297(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g298(.A(new_n428), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g299(.A1(new_n414), .A2(new_n418), .ZN(new_n437));
  OR2_X1    g300(.A1(new_n387), .A2(new_n388), .ZN(new_n438));
  NAND2_X1  g301(.A1(new_n438), .A2(new_n425), .ZN(new_n439));
  INV_X1    g302(.A(new_n386), .ZN(new_n440));
  AOI22_X1  g303(.A1(new_n317), .A2(new_n357), .B1(new_n375), .B2(new_n376), .ZN(new_n441));
  AOI22_X1  g304(.A1(new_n439), .A2(new_n420), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g305(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g306(.A1(new_n443), .A2(new_n422), .ZN(new_n444));
  NAND3_X1  g307(.A1(new_n444), .A2(KEYINPUT39), .A3(new_n434), .ZN(new_n445));
  NAND3_X1  g308(.A1(new_n436), .A2(new_n239), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g309(.A1(new_n425), .A2(G1gat), .ZN(new_n447));
  OAI21_X1  g310(.A(new_n427), .B1(new_n446), .B2(new_n447), .ZN(G1324gat));
  NOR2_X1   g311(.A1(new_n438), .A2(G8gat), .ZN(new_n449));
  NAND4_X1  g312(.A1(new_n436), .A2(new_n239), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  INV_X1    g313(.A(KEYINPUT40), .ZN(new_n451));
  OAI211_X1 g314(.A(new_n451), .B(G8gat), .C1(new_n424), .C2(new_n438), .ZN(new_n452));
  INV_X1    g315(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g316(.A1(new_n444), .A2(new_n389), .A3(new_n182), .A4(new_n263), .ZN(new_n454));
  AOI21_X1  g317(.A(new_n451), .B1(new_n454), .B2(G8gat), .ZN(new_n455));
  OAI21_X1  g318(.A(new_n450), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g319(.A(KEYINPUT41), .ZN(new_n457));
  NAND2_X1  g320(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g321(.A(KEYINPUT41), .B(new_n450), .C1(new_n453), .C2(new_n455), .ZN(new_n459));
  NAND2_X1  g322(.A1(new_n458), .A2(new_n459), .ZN(G1325gat));
  NOR3_X1   g323(.A1(new_n424), .A2(new_n184), .A3(new_n437), .ZN(new_n461));
  NAND2_X1  g324(.A1(new_n417), .A2(new_n411), .ZN(new_n462));
  NAND4_X1  g325(.A1(new_n436), .A2(new_n462), .A3(new_n239), .A4(new_n445), .ZN(new_n463));
  AOI21_X1  g326(.A(new_n461), .B1(new_n463), .B2(new_n184), .ZN(G1326gat));
  NOR3_X1   g327(.A1(new_n424), .A2(new_n185), .A3(new_n377), .ZN(new_n465));
  OR2_X1    g328(.A1(new_n446), .A2(new_n377), .ZN(new_n466));
  AOI21_X1  g329(.A(new_n465), .B1(new_n466), .B2(new_n185), .ZN(G1327gat));
  INV_X1    g330(.A(new_n224), .ZN(new_n468));
  NOR2_X1   g331(.A1(new_n468), .A2(new_n182), .ZN(new_n469));
  NOR2_X1   g332(.A1(new_n240), .A2(new_n262), .ZN(new_n470));
  NAND3_X1  g333(.A1(new_n444), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g334(.A1(new_n471), .A2(new_n425), .ZN(new_n472));
  XNOR2_X1  g335(.A(KEYINPUT42), .B(G29gat), .ZN(new_n473));
  XNOR2_X1  g336(.A(new_n472), .B(new_n473), .ZN(G1328gat));
  NOR2_X1   g337(.A1(new_n471), .A2(new_n438), .ZN(new_n475));
  XOR2_X1   g338(.A(KEYINPUT43), .B(G36gat), .Z(new_n476));
  XNOR2_X1  g339(.A(new_n475), .B(new_n476), .ZN(G1329gat));
  OAI21_X1  g340(.A(G43gat), .B1(new_n471), .B2(new_n437), .ZN(new_n478));
  INV_X1    g341(.A(G43gat), .ZN(new_n479));
  NAND2_X1  g342(.A1(new_n462), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g343(.A(new_n478), .B1(new_n471), .B2(new_n480), .ZN(new_n481));
  INV_X1    g344(.A(KEYINPUT44), .ZN(new_n482));
  XNOR2_X1  g345(.A(new_n481), .B(new_n482), .ZN(G1330gat));
  NOR2_X1   g346(.A1(new_n471), .A2(new_n377), .ZN(new_n484));
  XOR2_X1   g347(.A(new_n484), .B(G50gat), .Z(G1331gat));
  NOR2_X1   g348(.A1(new_n429), .A2(new_n433), .ZN(new_n486));
  INV_X1    g349(.A(new_n255), .ZN(new_n487));
  AND3_X1   g350(.A1(new_n260), .A2(KEYINPUT18), .A3(new_n253), .ZN(new_n488));
  AOI21_X1  g351(.A(KEYINPUT18), .B1(new_n260), .B2(new_n253), .ZN(new_n489));
  OAI21_X1  g352(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g353(.A1(new_n224), .A2(new_n490), .A3(new_n239), .ZN(new_n491));
  NAND2_X1  g354(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g355(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g356(.A1(new_n493), .A2(new_n317), .ZN(new_n494));
  XNOR2_X1  g357(.A(new_n494), .B(G57gat), .ZN(G1332gat));
  INV_X1    g358(.A(G64gat), .ZN(new_n496));
  NAND3_X1  g359(.A1(new_n493), .A2(new_n496), .A3(new_n389), .ZN(new_n497));
  INV_X1    g360(.A(KEYINPUT45), .ZN(new_n498));
  NAND2_X1  g361(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g362(.A1(new_n493), .A2(KEYINPUT45), .A3(new_n496), .A4(new_n389), .ZN(new_n500));
  OAI21_X1  g363(.A(G64gat), .B1(new_n492), .B2(new_n438), .ZN(new_n501));
  NAND3_X1  g364(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(G1333gat));
  INV_X1    g365(.A(G71gat), .ZN(new_n503));
  NOR3_X1   g366(.A1(new_n492), .A2(new_n503), .A3(new_n437), .ZN(new_n504));
  NAND2_X1  g367(.A1(new_n493), .A2(new_n462), .ZN(new_n505));
  AOI21_X1  g368(.A(new_n504), .B1(new_n503), .B2(new_n505), .ZN(G1334gat));
  NAND2_X1  g369(.A1(new_n493), .A2(new_n420), .ZN(new_n507));
  XNOR2_X1  g370(.A(new_n507), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g371(.A1(new_n444), .A2(new_n469), .ZN(new_n509));
  NOR2_X1   g372(.A1(new_n490), .A2(new_n239), .ZN(new_n510));
  NAND2_X1  g373(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g374(.A1(new_n511), .A2(new_n425), .ZN(new_n512));
  INV_X1    g375(.A(G85gat), .ZN(new_n513));
  XNOR2_X1  g376(.A(new_n512), .B(new_n513), .ZN(G1336gat));
  NOR2_X1   g377(.A1(new_n511), .A2(new_n438), .ZN(new_n515));
  AND2_X1   g378(.A1(KEYINPUT46), .A2(G92gat), .ZN(new_n516));
  NOR2_X1   g379(.A1(KEYINPUT46), .A2(G92gat), .ZN(new_n517));
  OAI21_X1  g380(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g381(.A(new_n518), .B1(new_n515), .B2(new_n517), .ZN(G1337gat));
  NOR3_X1   g382(.A1(new_n511), .A2(new_n409), .A3(new_n437), .ZN(new_n520));
  NAND3_X1  g383(.A1(new_n509), .A2(new_n462), .A3(new_n510), .ZN(new_n521));
  AOI21_X1  g384(.A(new_n520), .B1(new_n409), .B2(new_n521), .ZN(G1338gat));
  NAND3_X1  g385(.A1(new_n509), .A2(new_n420), .A3(new_n510), .ZN(new_n523));
  XNOR2_X1  g386(.A(new_n523), .B(G106gat), .ZN(G1339gat));
  NAND4_X1  g387(.A1(new_n468), .A2(new_n182), .A3(new_n262), .A4(new_n239), .ZN(new_n525));
  INV_X1    g388(.A(KEYINPUT50), .ZN(new_n526));
  INV_X1    g389(.A(KEYINPUT47), .ZN(new_n527));
  OAI21_X1  g390(.A(new_n238), .B1(new_n229), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g391(.A1(new_n232), .A2(new_n528), .A3(new_n233), .ZN(new_n529));
  AOI21_X1  g392(.A(new_n528), .B1(new_n232), .B2(new_n233), .ZN(new_n530));
  NOR2_X1   g393(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g394(.A(KEYINPUT48), .B1(new_n262), .B2(new_n531), .ZN(new_n532));
  INV_X1    g395(.A(KEYINPUT48), .ZN(new_n533));
  OR2_X1    g396(.A1(new_n529), .A2(new_n530), .ZN(new_n534));
  NAND3_X1  g397(.A1(new_n490), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g398(.A1(new_n532), .A2(new_n535), .A3(new_n182), .ZN(new_n536));
  NOR2_X1   g399(.A1(new_n257), .A2(new_n258), .ZN(new_n537));
  NOR2_X1   g400(.A1(new_n537), .A2(KEYINPUT49), .ZN(new_n538));
  AOI21_X1  g401(.A(new_n538), .B1(new_n433), .B2(new_n531), .ZN(new_n539));
  NAND2_X1  g402(.A1(new_n239), .A2(new_n182), .ZN(new_n540));
  AOI21_X1  g403(.A(new_n252), .B1(new_n247), .B2(new_n249), .ZN(new_n541));
  AOI21_X1  g404(.A(new_n251), .B1(new_n245), .B2(new_n246), .ZN(new_n542));
  OR2_X1    g405(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI22_X1  g406(.A1(new_n243), .A2(new_n543), .B1(new_n537), .B2(KEYINPUT49), .ZN(new_n544));
  NAND3_X1  g407(.A1(new_n539), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g408(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g409(.A(new_n526), .B1(new_n546), .B2(new_n224), .ZN(new_n547));
  AOI211_X1 g410(.A(KEYINPUT50), .B(new_n468), .C1(new_n536), .C2(new_n545), .ZN(new_n548));
  OAI21_X1  g411(.A(new_n525), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g412(.A1(new_n549), .A2(new_n377), .ZN(new_n550));
  AOI211_X1 g413(.A(new_n425), .B(new_n389), .C1(new_n417), .C2(new_n411), .ZN(new_n551));
  NAND2_X1  g414(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g415(.A(G113gat), .B1(new_n552), .B2(new_n262), .ZN(new_n553));
  NAND2_X1  g416(.A1(new_n421), .A2(new_n317), .ZN(new_n554));
  INV_X1    g417(.A(new_n554), .ZN(new_n555));
  AND2_X1   g418(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g419(.A1(new_n556), .A2(new_n438), .ZN(new_n557));
  OAI21_X1  g420(.A(KEYINPUT51), .B1(new_n262), .B2(G113gat), .ZN(new_n558));
  OAI21_X1  g421(.A(new_n558), .B1(KEYINPUT51), .B2(G113gat), .ZN(new_n559));
  OAI21_X1  g422(.A(new_n553), .B1(new_n557), .B2(new_n559), .ZN(G1340gat));
  NOR2_X1   g423(.A1(new_n239), .A2(G120gat), .ZN(new_n561));
  NAND3_X1  g424(.A1(new_n556), .A2(new_n438), .A3(new_n561), .ZN(new_n562));
  INV_X1    g425(.A(KEYINPUT52), .ZN(new_n563));
  OR2_X1    g426(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g427(.A(G120gat), .B1(new_n552), .B2(new_n239), .ZN(new_n565));
  NAND2_X1  g428(.A1(new_n562), .A2(new_n563), .ZN(new_n566));
  NAND3_X1  g429(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G1341gat));
  NAND4_X1  g430(.A1(new_n549), .A2(new_n551), .A3(new_n377), .A4(new_n468), .ZN(new_n568));
  NAND2_X1  g431(.A1(new_n568), .A2(G127gat), .ZN(new_n569));
  NOR3_X1   g432(.A1(new_n224), .A2(G127gat), .A3(new_n389), .ZN(new_n570));
  NAND3_X1  g433(.A1(new_n549), .A2(new_n555), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g434(.A1(new_n571), .A2(KEYINPUT53), .ZN(new_n572));
  INV_X1    g435(.A(KEYINPUT53), .ZN(new_n573));
  NAND4_X1  g436(.A1(new_n549), .A2(new_n573), .A3(new_n555), .A4(new_n570), .ZN(new_n574));
  NAND3_X1  g437(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g438(.A(KEYINPUT54), .ZN(new_n576));
  NAND2_X1  g439(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g440(.A1(new_n569), .A2(new_n572), .A3(KEYINPUT54), .A4(new_n574), .ZN(new_n578));
  NAND2_X1  g441(.A1(new_n577), .A2(new_n578), .ZN(G1342gat));
  INV_X1    g442(.A(G134gat), .ZN(new_n580));
  NOR2_X1   g443(.A1(new_n389), .A2(new_n182), .ZN(new_n581));
  NAND3_X1  g444(.A1(new_n556), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g445(.A(KEYINPUT55), .ZN(new_n583));
  OR2_X1    g446(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g447(.A(G134gat), .B1(new_n552), .B2(new_n182), .ZN(new_n585));
  NAND2_X1  g448(.A1(new_n582), .A2(new_n583), .ZN(new_n586));
  NAND3_X1  g449(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G1343gat));
  AOI21_X1  g450(.A(new_n377), .B1(new_n414), .B2(new_n418), .ZN(new_n588));
  NAND4_X1  g451(.A1(new_n549), .A2(new_n317), .A3(new_n438), .A4(new_n588), .ZN(new_n589));
  NOR2_X1   g452(.A1(new_n589), .A2(new_n262), .ZN(new_n590));
  XNOR2_X1  g453(.A(new_n590), .B(new_n264), .ZN(G1344gat));
  INV_X1    g454(.A(KEYINPUT56), .ZN(new_n592));
  AND4_X1   g455(.A1(new_n317), .A2(new_n549), .A3(new_n438), .A4(new_n588), .ZN(new_n593));
  NAND2_X1  g456(.A1(new_n593), .A2(new_n240), .ZN(new_n594));
  OAI21_X1  g457(.A(new_n592), .B1(new_n594), .B2(new_n277), .ZN(new_n595));
  OR4_X1    g458(.A1(new_n592), .A2(new_n589), .A3(new_n277), .A4(new_n239), .ZN(new_n596));
  NAND2_X1  g459(.A1(new_n594), .A2(G148gat), .ZN(new_n597));
  NAND3_X1  g460(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G1345gat));
  AOI21_X1  g461(.A(G155gat), .B1(new_n593), .B2(new_n468), .ZN(new_n599));
  INV_X1    g462(.A(new_n271), .ZN(new_n600));
  NOR3_X1   g463(.A1(new_n589), .A2(new_n600), .A3(new_n224), .ZN(new_n601));
  OAI21_X1  g464(.A(KEYINPUT57), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g465(.A1(new_n593), .A2(new_n271), .A3(new_n468), .ZN(new_n603));
  INV_X1    g466(.A(KEYINPUT57), .ZN(new_n604));
  OAI21_X1  g467(.A(new_n273), .B1(new_n589), .B2(new_n224), .ZN(new_n605));
  NAND3_X1  g468(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g469(.A1(new_n602), .A2(new_n606), .ZN(G1346gat));
  NAND2_X1  g470(.A1(new_n549), .A2(new_n588), .ZN(new_n608));
  NOR2_X1   g471(.A1(new_n608), .A2(new_n425), .ZN(new_n609));
  NAND2_X1  g472(.A1(new_n609), .A2(new_n581), .ZN(new_n610));
  OAI21_X1  g473(.A(KEYINPUT58), .B1(new_n610), .B2(G162gat), .ZN(new_n611));
  NAND2_X1  g474(.A1(new_n610), .A2(G162gat), .ZN(new_n612));
  INV_X1    g475(.A(KEYINPUT58), .ZN(new_n613));
  NAND4_X1  g476(.A1(new_n609), .A2(new_n613), .A3(new_n274), .A4(new_n581), .ZN(new_n614));
  NAND3_X1  g477(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(G1347gat));
  NOR2_X1   g478(.A1(new_n438), .A2(new_n317), .ZN(new_n616));
  NAND3_X1  g479(.A1(new_n550), .A2(new_n462), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g480(.A(G169gat), .B1(new_n617), .B2(new_n262), .ZN(new_n618));
  NAND3_X1  g481(.A1(new_n549), .A2(new_n421), .A3(new_n616), .ZN(new_n619));
  OR2_X1    g482(.A1(new_n262), .A2(G169gat), .ZN(new_n620));
  OAI21_X1  g483(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(G1348gat));
  OAI21_X1  g484(.A(G176gat), .B1(new_n617), .B2(new_n239), .ZN(new_n622));
  OR2_X1    g485(.A1(new_n239), .A2(G176gat), .ZN(new_n623));
  OAI21_X1  g486(.A(new_n622), .B1(new_n619), .B2(new_n623), .ZN(G1349gat));
  OAI21_X1  g487(.A(G183gat), .B1(new_n617), .B2(new_n224), .ZN(new_n625));
  OR2_X1    g488(.A1(new_n224), .A2(G183gat), .ZN(new_n626));
  OAI21_X1  g489(.A(new_n625), .B1(new_n619), .B2(new_n626), .ZN(G1350gat));
  OAI21_X1  g490(.A(G190gat), .B1(new_n617), .B2(new_n182), .ZN(new_n628));
  OR2_X1    g491(.A1(new_n182), .A2(G190gat), .ZN(new_n629));
  OAI21_X1  g492(.A(new_n628), .B1(new_n619), .B2(new_n629), .ZN(G1351gat));
  AOI21_X1  g493(.A(new_n262), .B1(KEYINPUT59), .B2(G197gat), .ZN(new_n631));
  NAND4_X1  g494(.A1(new_n549), .A2(new_n588), .A3(new_n616), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g495(.A1(KEYINPUT59), .A2(G197gat), .ZN(new_n633));
  XOR2_X1   g496(.A(new_n632), .B(new_n633), .Z(G1352gat));
  NAND4_X1  g497(.A1(new_n549), .A2(new_n240), .A3(new_n588), .A4(new_n616), .ZN(new_n635));
  NOR2_X1   g498(.A1(new_n635), .A2(new_n326), .ZN(new_n636));
  AND2_X1   g499(.A1(new_n636), .A2(KEYINPUT60), .ZN(new_n637));
  NOR2_X1   g500(.A1(new_n636), .A2(KEYINPUT60), .ZN(new_n638));
  NAND2_X1  g501(.A1(new_n635), .A2(G204gat), .ZN(new_n639));
  AOI21_X1  g502(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(G1353gat));
  NAND4_X1  g503(.A1(new_n549), .A2(new_n468), .A3(new_n588), .A4(new_n616), .ZN(new_n641));
  INV_X1    g504(.A(KEYINPUT62), .ZN(new_n642));
  INV_X1    g505(.A(G211gat), .ZN(new_n643));
  NAND2_X1  g506(.A1(new_n643), .A2(KEYINPUT61), .ZN(new_n644));
  NAND3_X1  g507(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g508(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g509(.A(new_n642), .B1(new_n641), .B2(new_n644), .ZN(new_n647));
  OAI22_X1  g510(.A1(new_n646), .A2(new_n647), .B1(KEYINPUT61), .B2(new_n643), .ZN(new_n648));
  INV_X1    g511(.A(new_n647), .ZN(new_n649));
  NOR2_X1   g512(.A1(new_n643), .A2(KEYINPUT61), .ZN(new_n650));
  NAND3_X1  g513(.A1(new_n649), .A2(new_n650), .A3(new_n645), .ZN(new_n651));
  NAND2_X1  g514(.A1(new_n648), .A2(new_n651), .ZN(G1354gat));
  NAND4_X1  g515(.A1(new_n549), .A2(new_n433), .A3(new_n588), .A4(new_n616), .ZN(new_n653));
  XOR2_X1   g516(.A(KEYINPUT63), .B(G218gat), .Z(new_n654));
  XNOR2_X1  g517(.A(new_n653), .B(new_n654), .ZN(G1355gat));
endmodule


