//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G97), .A2(G257), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G87), .A2(G250), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G77), .A2(G244), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G116), .ZN(new_n217));
  INV_X1    g0017(.A(G270), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n206), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NAND2_X1  g0021(.A1(new_n203), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(G20), .A3(new_n225), .ZN(new_n226));
  OR3_X1    g0026(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n227));
  OAI21_X1  g0027(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n221), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n218), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n217), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  INV_X1    g0049(.A(G20), .ZN(new_n250));
  NOR3_X1   g0050(.A1(new_n249), .A2(new_n250), .A3(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n224), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(KEYINPUT68), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(new_n250), .B2(G1), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G58), .A2(G68), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n250), .B1(new_n263), .B2(new_n261), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n250), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT8), .B(G58), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI211_X1 g0073(.A(new_n264), .B(new_n268), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n253), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n260), .B(new_n262), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(KEYINPUT72), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n278), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G222), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G223), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n290), .B1(new_n291), .B2(new_n288), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n225), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n283), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n296), .A2(new_n281), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n279), .A2(new_n280), .B1(G200), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n277), .A2(KEYINPUT72), .ZN(new_n303));
  INV_X1    g0103(.A(G190), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT73), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT73), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n298), .A2(new_n306), .A3(G190), .A4(new_n300), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n302), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n302), .A2(KEYINPUT10), .A3(new_n303), .A4(new_n308), .ZN(new_n312));
  INV_X1    g0112(.A(new_n301), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n276), .B1(new_n313), .B2(G169), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT69), .B(new_n276), .C1(new_n313), .C2(G169), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(G179), .C2(new_n301), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n311), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G20), .A2(G77), .ZN(new_n321));
  XOR2_X1   g0121(.A(KEYINPUT15), .B(G87), .Z(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT70), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n272), .B(new_n324), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n321), .B1(new_n269), .B2(new_n323), .C1(new_n325), .C2(new_n266), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n253), .B1(new_n291), .B2(new_n251), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n259), .A2(G77), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n288), .A2(G232), .A3(new_n289), .ZN(new_n330));
  INV_X1    g0130(.A(G107), .ZN(new_n331));
  INV_X1    g0131(.A(G238), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n330), .B1(new_n331), .B2(new_n288), .C1(new_n292), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n297), .ZN(new_n334));
  INV_X1    g0134(.A(new_n283), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n299), .A2(G244), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n329), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(G200), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n334), .A2(G190), .A3(new_n335), .A4(new_n336), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n344), .A2(new_n327), .A3(new_n345), .A4(new_n328), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n319), .B1(new_n320), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT80), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n265), .A2(G159), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G58), .A2(G68), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n203), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n357), .A2(KEYINPUT76), .A3(G20), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT76), .B1(new_n357), .B2(G20), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n352), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n286), .A2(new_n250), .A3(new_n287), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n250), .A4(new_n287), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n202), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n351), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n359), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n357), .A2(KEYINPUT76), .A3(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(KEYINPUT3), .A2(G33), .ZN(new_n370));
  NOR2_X1   g0170(.A1(KEYINPUT3), .A2(G33), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT7), .B1(new_n372), .B2(new_n250), .ZN(new_n373));
  INV_X1    g0173(.A(new_n364), .ZN(new_n374));
  OAI21_X1  g0174(.A(G68), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n375), .A4(new_n352), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(new_n376), .A3(new_n253), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n259), .A2(new_n273), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n272), .A2(new_n251), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(G223), .B(new_n289), .C1(new_n370), .C2(new_n371), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n288), .A2(KEYINPUT77), .A3(G223), .A4(new_n289), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n288), .A2(G226), .A3(G1698), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n297), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n283), .B1(new_n299), .B2(G232), .ZN(new_n389));
  AOI21_X1  g0189(.A(G200), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT78), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(KEYINPUT78), .A3(new_n297), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n389), .A2(new_n304), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n350), .B1(new_n380), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n399), .A2(new_n396), .A3(KEYINPUT17), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n349), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n380), .A2(new_n350), .A3(new_n397), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT17), .B1(new_n399), .B2(new_n396), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(KEYINPUT80), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n394), .A2(new_n338), .A3(new_n389), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n388), .A2(new_n389), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n341), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n405), .A4(new_n407), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(KEYINPUT79), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n401), .B(new_n404), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n271), .A2(G77), .B1(G50), .B2(new_n265), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n202), .A2(G20), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n275), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(KEYINPUT11), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n249), .A2(G1), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT74), .B1(new_n421), .B2(new_n417), .ZN(new_n422));
  XOR2_X1   g0222(.A(new_n422), .B(KEYINPUT12), .Z(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(KEYINPUT11), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n259), .A2(G68), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n419), .A2(new_n423), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n288), .A2(G226), .A3(new_n289), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n283), .B1(new_n430), .B2(new_n297), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n299), .A2(G238), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n435), .A3(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n426), .B1(new_n437), .B2(G200), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n304), .B2(new_n437), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n431), .A2(new_n435), .A3(new_n432), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n441));
  OAI21_X1  g0241(.A(G169), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT14), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(new_n444), .A3(G169), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n434), .A2(G179), .A3(new_n436), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n426), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n343), .A2(KEYINPUT71), .A3(new_n346), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n439), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n348), .A2(new_n415), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n348), .A2(new_n415), .A3(new_n453), .A4(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n456), .A2(new_n458), .B1(new_n225), .B2(new_n295), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n255), .A2(G45), .ZN(new_n460));
  OR2_X1    g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n459), .A2(G270), .B1(G274), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(G257), .B(new_n289), .C1(new_n370), .C2(new_n371), .ZN(new_n465));
  OAI211_X1 g0265(.A(G264), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n286), .A2(G303), .A3(new_n287), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n297), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n420), .A2(G20), .A3(new_n217), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n420), .A2(G20), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n255), .A2(G33), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n275), .A2(new_n472), .A3(G116), .A4(new_n473), .ZN(new_n474));
  AOI22_X1  g0274(.A1(new_n252), .A2(new_n224), .B1(G20), .B2(new_n217), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n250), .C1(G33), .C2(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n475), .A2(KEYINPUT20), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT20), .B1(new_n475), .B2(new_n478), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n471), .B(new_n474), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n470), .A2(G169), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT85), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT85), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n470), .A2(new_n481), .A3(new_n485), .A4(G169), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n484), .B(new_n341), .C1(new_n464), .C2(new_n469), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n470), .A2(new_n338), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n481), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n470), .A2(G200), .ZN(new_n491));
  INV_X1    g0291(.A(new_n481), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n491), .B(new_n492), .C1(new_n304), .C2(new_n470), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n487), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT83), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n472), .A2(G97), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n254), .A2(new_n473), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(new_n477), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n331), .B1(new_n363), .B2(new_n364), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n266), .A2(new_n291), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT6), .ZN(new_n503));
  AND2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G97), .A2(G107), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n331), .A2(KEYINPUT6), .A3(G97), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n250), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n501), .A2(new_n502), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n500), .B1(new_n509), .B2(new_n275), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(new_n289), .C1(new_n370), .C2(new_n371), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n289), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n476), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n297), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n462), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n458), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n296), .A3(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n463), .A2(G274), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT82), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT82), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n518), .B(new_n338), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n510), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n523), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT82), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n513), .A2(new_n514), .A3(new_n516), .A4(new_n476), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n530), .A2(new_n531), .B1(new_n297), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G169), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n495), .B1(new_n527), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n518), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n341), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(KEYINPUT83), .A3(new_n526), .A4(new_n510), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n525), .A2(new_n524), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n513), .A2(new_n514), .ZN(new_n542));
  INV_X1    g0342(.A(new_n517), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n296), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(G200), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(G190), .A3(new_n518), .ZN(new_n546));
  OAI21_X1  g0346(.A(G107), .B1(new_n373), .B2(new_n374), .ZN(new_n547));
  INV_X1    g0347(.A(new_n502), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n506), .A2(new_n507), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n547), .B(new_n548), .C1(new_n250), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n499), .B1(new_n550), .B2(new_n253), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n494), .A2(new_n540), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(G33), .A2(G41), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n460), .B(G250), .C1(new_n555), .C2(new_n224), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G244), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n558));
  OAI211_X1 g0358(.A(G238), .B(new_n289), .C1(new_n370), .C2(new_n371), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n557), .B1(new_n561), .B2(new_n297), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n460), .A2(new_n282), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(G190), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT84), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n563), .B(new_n557), .C1(new_n561), .C2(new_n297), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT84), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(G190), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n250), .B1(new_n429), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n505), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n250), .B(G68), .C1(new_n370), .C2(new_n371), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n571), .B1(new_n429), .B2(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n253), .B1(new_n251), .B2(new_n323), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n254), .A2(G87), .A3(new_n473), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n562), .A2(new_n564), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(G200), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n341), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n254), .A2(new_n322), .A3(new_n473), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n567), .A2(new_n338), .B1(new_n585), .B2(new_n579), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n570), .A2(new_n583), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n250), .B(G87), .C1(new_n370), .C2(new_n371), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n288), .A2(new_n590), .A3(new_n250), .A4(G87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n560), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n250), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n250), .A2(G107), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT23), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n592), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(KEYINPUT24), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n589), .A2(new_n591), .B1(new_n250), .B2(new_n593), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n596), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n253), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G257), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n603));
  OAI211_X1 g0403(.A(G250), .B(new_n289), .C1(new_n370), .C2(new_n371), .ZN(new_n604));
  OR2_X1    g0404(.A1(KEYINPUT86), .A2(G294), .ZN(new_n605));
  NAND2_X1  g0405(.A1(KEYINPUT86), .A2(G294), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(G33), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT87), .A4(new_n607), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n297), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n459), .A2(G264), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n523), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n251), .A2(new_n331), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT25), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n498), .A2(new_n331), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n612), .A2(G190), .A3(new_n523), .A4(new_n613), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n602), .A2(new_n615), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n614), .A2(new_n341), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n612), .A2(new_n338), .A3(new_n523), .A4(new_n613), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n597), .A2(KEYINPUT24), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n600), .A2(new_n599), .A3(new_n596), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n275), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n619), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n622), .B(new_n623), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n587), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n455), .A2(new_n554), .A3(new_n629), .ZN(G372));
  AND2_X1   g0430(.A1(new_n487), .A2(new_n490), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n628), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n552), .B1(new_n535), .B2(new_n539), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n584), .A2(KEYINPUT88), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT88), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n582), .B2(new_n341), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n586), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n570), .A2(new_n583), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n632), .A2(new_n633), .A3(new_n621), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT89), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n527), .A2(new_n534), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n637), .A2(new_n638), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n645), .B1(new_n631), .B2(new_n628), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT89), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n633), .A4(new_n621), .ZN(new_n648));
  INV_X1    g0448(.A(new_n637), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n535), .A2(new_n587), .A3(new_n539), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n641), .A2(new_n644), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n455), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n318), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n448), .A2(new_n343), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n655), .A2(new_n401), .A3(new_n404), .A4(new_n439), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n410), .A2(new_n411), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n311), .A2(new_n312), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n654), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n255), .A2(new_n250), .A3(G13), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT27), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(KEYINPUT91), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(KEYINPUT91), .ZN(new_n670));
  OAI211_X1 g0470(.A(G213), .B(new_n667), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n481), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n631), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n494), .A2(new_n674), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n631), .A2(new_n673), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n628), .A2(new_n673), .ZN(new_n682));
  INV_X1    g0482(.A(new_n628), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n673), .B1(new_n626), .B2(new_n627), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n621), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n681), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n681), .A2(new_n685), .B1(new_n628), .B2(new_n673), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n688), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  INV_X1    g0491(.A(new_n673), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n652), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT94), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n652), .B2(new_n692), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n691), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n640), .A3(new_n637), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .A3(new_n692), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT95), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT95), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n697), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n554), .A2(new_n705), .A3(new_n629), .A4(new_n692), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n629), .A2(new_n633), .A3(new_n494), .A4(new_n692), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n489), .A2(new_n533), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n567), .A2(new_n612), .A3(new_n613), .ZN(new_n711));
  OR3_X1    g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n537), .A2(new_n338), .A3(new_n582), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n614), .A2(new_n470), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n712), .B(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n533), .A2(G179), .A3(new_n567), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT92), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n470), .A4(new_n614), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT92), .B1(new_n714), .B2(new_n715), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n712), .A2(new_n720), .A3(new_n721), .A4(new_n713), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n673), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n706), .A2(new_n708), .A3(new_n717), .A4(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n704), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT96), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT96), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n704), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n255), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n229), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G41), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n574), .A2(G116), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n735), .A2(new_n255), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n223), .B2(new_n735), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT28), .Z(new_n740));
  NAND2_X1  g0540(.A1(new_n733), .A2(new_n740), .ZN(G364));
  AOI21_X1  g0541(.A(new_n224), .B1(G20), .B2(new_n341), .ZN(new_n742));
  OR3_X1    g0542(.A1(new_n304), .A2(G179), .A3(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n250), .A2(new_n338), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(new_n304), .A3(G200), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n745), .A2(new_n477), .B1(new_n747), .B2(new_n202), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G200), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n372), .B1(new_n751), .B2(G58), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT32), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n250), .A2(G179), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G190), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n754), .A2(new_n304), .A3(G200), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n752), .B1(new_n753), .B2(new_n758), .C1(new_n331), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n746), .A2(new_n755), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n291), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n758), .A2(new_n753), .B1(new_n764), .B2(G87), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n261), .B2(new_n766), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n749), .A2(new_n760), .A3(new_n762), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n759), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n764), .A2(G303), .B1(new_n769), .B2(G283), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n605), .A2(new_n606), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(new_n745), .ZN(new_n772));
  INV_X1    g0572(.A(new_n766), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G326), .ZN(new_n774));
  INV_X1    g0574(.A(new_n751), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n761), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G329), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI221_X1 g0581(.A(new_n372), .B1(new_n756), .B2(new_n780), .C1(new_n747), .C2(new_n781), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n772), .A2(new_n777), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n742), .B1(new_n768), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n244), .A2(G45), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n734), .A2(new_n288), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n785), .B(new_n786), .C1(G45), .C2(new_n222), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n229), .A2(G355), .A3(new_n288), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(G116), .C2(new_n229), .ZN(new_n789));
  INV_X1    g0589(.A(new_n742), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n250), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n677), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n784), .B(new_n795), .C1(new_n796), .C2(new_n792), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n249), .A2(G20), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n255), .B1(new_n798), .B2(G45), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n735), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n801), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n796), .A2(G330), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n679), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT98), .Z(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n343), .A2(new_n692), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n343), .A2(KEYINPUT102), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT102), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n329), .A2(new_n339), .A3(new_n342), .A4(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n329), .A2(new_n673), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n346), .ZN(new_n816));
  OAI211_X1 g0616(.A(KEYINPUT103), .B(new_n810), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT103), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n816), .B1(new_n811), .B2(new_n813), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n809), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n694), .B2(new_n696), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n652), .A2(new_n692), .A3(new_n821), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(new_n727), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n727), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n803), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G137), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n747), .A2(new_n267), .B1(new_n766), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT100), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n832), .B2(new_n775), .C1(new_n757), .C2(new_n761), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT34), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n745), .A2(new_n201), .B1(new_n759), .B2(new_n202), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n372), .B(new_n835), .C1(G50), .C2(new_n764), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(new_n836), .C1(new_n837), .C2(new_n756), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n763), .A2(new_n331), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n759), .A2(new_n573), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n839), .B(new_n840), .C1(G303), .C2(new_n773), .ZN(new_n841));
  INV_X1    g0641(.A(new_n747), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(G283), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n751), .A2(G294), .B1(new_n744), .B2(G97), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n372), .B1(new_n756), .B2(new_n778), .ZN(new_n845));
  INV_X1    g0645(.A(new_n761), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(G116), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n841), .A2(new_n843), .A3(new_n844), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n790), .B1(new_n838), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n742), .A2(new_n791), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n803), .B(new_n849), .C1(new_n291), .C2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT101), .Z(new_n854));
  INV_X1    g0654(.A(new_n791), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n821), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n828), .A2(new_n856), .ZN(G384));
  INV_X1    g0657(.A(new_n671), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n658), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n399), .A2(new_n858), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n414), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n380), .A2(new_n397), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n408), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n408), .A3(new_n866), .A4(new_n860), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n862), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n447), .A2(new_n426), .A3(new_n673), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT104), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n447), .A2(KEYINPUT104), .A3(new_n426), .A4(new_n673), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n426), .A2(new_n673), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n439), .A2(new_n448), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n814), .A2(new_n692), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n824), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  AOI221_X4 g0684(.A(new_n884), .B1(new_n865), .B2(new_n867), .C1(new_n414), .C2(new_n861), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n885), .B2(new_n869), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT106), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n868), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n398), .A2(new_n400), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n861), .B1(new_n657), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n865), .A2(KEYINPUT106), .A3(new_n867), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n871), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n448), .A2(new_n673), .ZN(new_n898));
  AOI221_X4 g0698(.A(new_n859), .B1(new_n872), .B2(new_n883), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n697), .A2(new_n455), .A3(new_n703), .A4(new_n702), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n661), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n899), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n706), .A2(new_n708), .A3(new_n725), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n880), .A3(new_n821), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n880), .A3(new_n821), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n894), .A2(new_n871), .B1(new_n907), .B2(KEYINPUT107), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n904), .A2(new_n821), .A3(new_n880), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n885), .B2(new_n869), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n906), .A2(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n455), .A2(new_n904), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(G330), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n902), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n255), .B2(new_n798), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT35), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n250), .B(new_n224), .C1(new_n549), .C2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(G116), .C1(new_n918), .C2(new_n549), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  AND4_X1   g0721(.A1(G77), .A2(new_n223), .A3(new_n355), .A4(new_n356), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n202), .A2(G50), .ZN(new_n923));
  OAI211_X1 g0723(.A(G1), .B(new_n249), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n921), .A3(new_n924), .ZN(G367));
  OAI22_X1  g0725(.A1(new_n747), .A2(new_n757), .B1(new_n761), .B2(new_n261), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n744), .A2(G68), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n927), .B1(new_n201), .B2(new_n763), .C1(new_n775), .C2(new_n267), .ZN(new_n928));
  INV_X1    g0728(.A(new_n756), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n926), .B(new_n928), .C1(G137), .C2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n288), .B1(new_n759), .B2(new_n291), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT113), .Z(new_n932));
  OAI211_X1 g0732(.A(new_n930), .B(new_n932), .C1(new_n832), .C2(new_n766), .ZN(new_n933));
  INV_X1    g0733(.A(G303), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n775), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n372), .B1(new_n759), .B2(new_n477), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G317), .B2(new_n929), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT112), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n764), .A2(KEYINPUT46), .A3(G116), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT46), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n763), .B2(new_n217), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n939), .B(new_n941), .C1(new_n771), .C2(new_n747), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT111), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(G283), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n766), .A2(new_n778), .B1(new_n761), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G107), .B2(new_n744), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n938), .A2(new_n944), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n933), .B1(new_n935), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT47), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n803), .B1(new_n951), .B2(new_n742), .ZN(new_n952));
  INV_X1    g0752(.A(new_n786), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n794), .B1(new_n229), .B2(new_n323), .C1(new_n240), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n673), .A2(new_n581), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n639), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n637), .B2(new_n955), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(new_n792), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n952), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n633), .B1(new_n551), .B2(new_n692), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n642), .A2(new_n673), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n962), .A2(new_n689), .A3(KEYINPUT44), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT44), .B1(new_n962), .B2(new_n689), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT109), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n962), .A2(new_n689), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n962), .B2(new_n689), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n967), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(new_n688), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n679), .B(new_n686), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n685), .A2(new_n682), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n680), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n973), .B(new_n976), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n704), .A2(new_n731), .A3(new_n728), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n731), .B1(new_n704), .B2(new_n728), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n972), .A2(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n735), .B(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n800), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n975), .A2(new_n962), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT42), .Z(new_n985));
  INV_X1    g0785(.A(new_n962), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n683), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n673), .B1(new_n987), .B2(new_n540), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n983), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n687), .A2(new_n962), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n990), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n992), .B1(new_n991), .B2(new_n993), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n959), .B1(new_n982), .B2(new_n996), .ZN(G387));
  INV_X1    g0797(.A(new_n977), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n978), .B2(new_n979), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n730), .A2(new_n732), .A3(new_n977), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n735), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n744), .A2(G283), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n751), .A2(G317), .B1(new_n846), .B2(G303), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n778), .B2(new_n747), .C1(new_n776), .C2(new_n766), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1002), .B1(new_n771), .B2(new_n763), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT114), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n929), .A2(G326), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(KEYINPUT49), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n288), .B1(new_n769), .B2(G116), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n751), .A2(G50), .B1(new_n744), .B2(new_n322), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n757), .B2(new_n766), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n291), .A2(new_n763), .B1(new_n759), .B2(new_n477), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n288), .B1(new_n756), .B2(new_n267), .C1(new_n747), .C2(new_n272), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n202), .B2(new_n761), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n790), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n974), .A2(new_n792), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n325), .A2(G50), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n737), .B1(G68), .B2(G77), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n457), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n953), .B1(new_n237), .B2(G45), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n734), .A2(new_n372), .A3(new_n736), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n734), .A2(new_n331), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n793), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1021), .A2(new_n803), .A3(new_n1022), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n998), .B2(new_n800), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1001), .A2(new_n1035), .ZN(G393));
  INV_X1    g0836(.A(new_n735), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n999), .B2(new_n972), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n971), .B(new_n687), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n998), .C1(new_n978), .C2(new_n979), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n800), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n794), .B1(new_n477), .B2(new_n229), .C1(new_n247), .C2(new_n953), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n331), .A2(new_n759), .B1(new_n763), .B2(new_n946), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n288), .B1(new_n846), .B2(G294), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n776), .B2(new_n756), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1044), .B(new_n1046), .C1(G303), .C2(new_n842), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n751), .B1(new_n773), .B2(G317), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1047), .B(new_n1050), .C1(new_n217), .C2(new_n745), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n775), .A2(new_n757), .B1(new_n766), .B2(new_n267), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n745), .A2(new_n291), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n840), .B(new_n1054), .C1(G68), .C2(new_n764), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n325), .A2(new_n761), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n372), .B1(new_n842), .B2(G50), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n756), .A2(new_n832), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1051), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n803), .B1(new_n1060), .B2(new_n742), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1043), .B(new_n1061), .C1(new_n986), .C2(new_n792), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1042), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1041), .A2(new_n1064), .ZN(G390));
  NAND3_X1  g0865(.A1(new_n726), .A2(G330), .A3(new_n821), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n881), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n821), .A2(new_n692), .A3(new_n700), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1069), .A2(new_n882), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n904), .A2(G330), .A3(new_n821), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n881), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT118), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT117), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1066), .A2(new_n1076), .A3(new_n881), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n1066), .B2(new_n881), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n907), .A2(new_n678), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n824), .A2(new_n882), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1075), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1066), .A2(new_n881), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT117), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1079), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1066), .A2(new_n1076), .A3(new_n881), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(KEYINPUT118), .A3(new_n1081), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1074), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n455), .A2(G330), .A3(new_n904), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n900), .A2(new_n661), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n886), .B(new_n896), .C1(new_n898), .C2(new_n883), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n894), .A2(new_n871), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n898), .B(KEYINPUT116), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n1070), .C2(new_n881), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1094), .A2(new_n1097), .A3(new_n1067), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1079), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1037), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1101), .B2(new_n1093), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n800), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n775), .A2(new_n837), .B1(new_n759), .B2(new_n261), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G159), .B2(new_n744), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n372), .B1(new_n929), .B2(G125), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n829), .B2(new_n747), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n846), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n773), .A2(G128), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n763), .A2(new_n267), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n766), .A2(new_n946), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1115), .B(new_n1054), .C1(G116), .C2(new_n751), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n764), .A2(G87), .B1(new_n769), .B2(G68), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n372), .B1(new_n747), .B2(new_n331), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G294), .B2(new_n929), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n761), .A2(new_n477), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1114), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1122), .A2(new_n742), .B1(new_n272), .B2(new_n852), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n801), .B(new_n1123), .C1(new_n897), .C2(new_n855), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1103), .A2(new_n1104), .A3(new_n1124), .ZN(G378));
  INV_X1    g0925(.A(new_n1092), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1100), .B2(new_n1090), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n319), .A2(KEYINPUT120), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT120), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n311), .A2(new_n1131), .A3(new_n312), .A4(new_n318), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n858), .A2(new_n276), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1129), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1133), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1128), .A3(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n912), .B2(G330), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n910), .A2(new_n911), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n907), .A2(KEYINPUT107), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1095), .A2(new_n906), .A3(new_n1145), .ZN(new_n1146));
  AND4_X1   g0946(.A1(G330), .A2(new_n1144), .A3(new_n1142), .A4(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n899), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT121), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n912), .A2(G330), .A3(new_n1142), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1144), .A2(new_n1146), .A3(G330), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1142), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n897), .A2(new_n898), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n859), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n872), .A2(new_n883), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1148), .A2(new_n1149), .A3(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(KEYINPUT121), .B(new_n899), .C1(new_n1143), .C2(new_n1147), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1127), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1127), .A2(KEYINPUT57), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n735), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1159), .A2(new_n800), .A3(new_n1160), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1142), .A2(new_n791), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n852), .A2(new_n261), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n747), .A2(new_n477), .B1(new_n756), .B2(new_n946), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n927), .B1(new_n217), .B2(new_n766), .C1(new_n775), .C2(new_n331), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n322), .C2(new_n846), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G41), .B(new_n288), .C1(new_n764), .C2(G77), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT119), .Z(new_n1174));
  OAI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(new_n201), .C2(new_n759), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT58), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n261), .B1(new_n370), .B2(G41), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n751), .A2(G128), .B1(new_n764), .B2(new_n1109), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n773), .A2(G125), .B1(new_n846), .B2(G137), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n744), .A2(G150), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n842), .A2(G132), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G33), .B1(new_n929), .B2(G124), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G41), .B1(new_n769), .B2(G159), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1176), .A2(new_n1177), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n803), .B1(new_n1188), .B2(new_n742), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1168), .A2(new_n1169), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1166), .A2(new_n1167), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT122), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT122), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1166), .A2(new_n1193), .A3(new_n1167), .A4(new_n1190), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(G375));
  AOI22_X1  g0995(.A1(G283), .A2(new_n751), .B1(new_n773), .B2(G294), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n477), .B2(new_n763), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n745), .A2(new_n323), .B1(new_n291), .B2(new_n759), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n372), .B1(new_n756), .B2(new_n934), .C1(new_n747), .C2(new_n217), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n331), .B2(new_n761), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n775), .A2(new_n829), .B1(new_n745), .B2(new_n261), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G159), .B2(new_n764), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n929), .A2(G128), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G132), .A2(new_n773), .B1(new_n769), .B2(G58), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n372), .B1(new_n842), .B2(new_n1109), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n267), .B2(new_n761), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1201), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT123), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n801), .B1(new_n790), .B2(new_n1211), .C1(new_n880), .C2(new_n855), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n202), .B2(new_n852), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1080), .A2(new_n1075), .A3(new_n1082), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT118), .B1(new_n1088), .B2(new_n1081), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1073), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1213), .B1(new_n1216), .B2(new_n800), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1092), .B(new_n1073), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n981), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1217), .B1(new_n1219), .B2(new_n1093), .ZN(G381));
  INV_X1    g1020(.A(G375), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1103), .A2(new_n1104), .A3(new_n1124), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G390), .A2(G381), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1001), .A2(new_n807), .A3(new_n1035), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G387), .A3(G384), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .A4(new_n1226), .ZN(G407));
  NAND3_X1  g1027(.A1(new_n1221), .A2(new_n672), .A3(new_n1222), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(G407), .A2(G213), .A3(new_n1228), .ZN(G409));
  AOI21_X1  g1029(.A(new_n807), .B1(new_n1001), .B2(new_n1035), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n959), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n730), .A2(new_n732), .B1(new_n1039), .B2(new_n998), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n981), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n799), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n994), .A2(new_n995), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1232), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(G390), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1063), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(G387), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1231), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(G390), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(new_n1239), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1166), .A2(G378), .A3(new_n1167), .A4(new_n1190), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1164), .A2(new_n800), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1190), .B(new_n1248), .C1(new_n1161), .C2(new_n1234), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1222), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n672), .A2(G213), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1216), .B2(new_n1126), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1218), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(KEYINPUT124), .B(new_n1218), .C1(new_n1093), .C2(new_n1254), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1037), .B1(new_n1256), .B2(KEYINPUT60), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1217), .B1(G384), .B2(KEYINPUT125), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1260), .A2(new_n1264), .A3(new_n1262), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1251), .A2(new_n1252), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1247), .A2(new_n1250), .B1(G213), .B2(new_n672), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1268), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n672), .A2(G213), .A3(G2897), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1267), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1264), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1276), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1266), .A2(new_n1267), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1275), .B1(new_n1282), .B2(new_n1271), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1246), .B1(new_n1274), .B2(new_n1283), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1277), .A2(new_n1278), .A3(new_n1276), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1280), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT126), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1271), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT126), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1279), .A2(new_n1289), .A3(new_n1281), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1291), .A2(KEYINPUT63), .B1(new_n1271), .B2(new_n1268), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1246), .A2(KEYINPUT61), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1269), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1284), .B1(new_n1292), .B2(new_n1295), .ZN(G405));
  AND3_X1   g1096(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1244), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1266), .B(new_n1267), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1241), .B(new_n1245), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT127), .B1(G375), .B2(new_n1222), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n1304), .B(G378), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1302), .B1(new_n1306), .B2(new_n1247), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1247), .ZN(new_n1308));
  NOR4_X1   g1108(.A1(new_n1303), .A2(new_n1305), .A3(new_n1301), .A4(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1307), .A2(new_n1309), .ZN(G402));
endmodule


