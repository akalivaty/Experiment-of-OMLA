//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n560, new_n561, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT67), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n461), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n464), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n473), .A2(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n484), .B1(new_n472), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G2105), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(G124), .B2(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(G114), .B2(new_n461), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n472), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n461), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n477), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n494), .B1(new_n496), .B2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n504), .A2(new_n508), .A3(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n510), .B2(new_n511), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n507), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n508), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(new_n508), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT72), .B(G89), .ZN(new_n522));
  OAI221_X1 g097(.A(new_n518), .B1(new_n519), .B2(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G168));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n521), .A2(new_n528), .B1(new_n519), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G171));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n521), .A2(new_n537), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n506), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT75), .ZN(G188));
  XNOR2_X1  g124(.A(KEYINPUT76), .B(G65), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n504), .A2(new_n550), .B1(G78), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n506), .ZN(new_n552));
  INV_X1    g127(.A(new_n521), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(G299));
  OR2_X1    g134(.A1(new_n535), .A2(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n535), .A2(KEYINPUT77), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(G301));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n516), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT78), .B(new_n507), .C1(new_n513), .C2(new_n515), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G303));
  NAND2_X1  g142(.A1(new_n553), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n509), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n521), .A2(new_n572), .B1(new_n519), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n506), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n553), .A2(G85), .B1(new_n509), .B2(G47), .ZN(new_n579));
  XOR2_X1   g154(.A(new_n579), .B(KEYINPUT80), .Z(new_n580));
  AOI22_X1  g155(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n506), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n580), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n553), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  AOI22_X1  g162(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n506), .B1(new_n589), .B2(new_n519), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT81), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n585), .B1(G868), .B2(new_n593), .ZN(G284));
  OAI21_X1  g169(.A(new_n585), .B1(G868), .B2(new_n593), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G868), .B2(new_n558), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(G868), .B2(new_n558), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n593), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n593), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n463), .A2(new_n501), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT13), .B(G2100), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n612), .B(new_n613), .C1(G111), .C2(new_n461), .ZN(new_n614));
  INV_X1    g189(.A(G135), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n472), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n488), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n609), .A2(new_n619), .ZN(G156));
  XOR2_X1   g195(.A(G1341), .B(G1348), .Z(new_n621));
  XOR2_X1   g196(.A(G2427), .B(G2430), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT85), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT84), .B(G2438), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n628), .B(new_n629), .Z(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n630), .A2(new_n633), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n621), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(KEYINPUT87), .ZN(new_n637));
  NOR3_X1   g212(.A1(new_n634), .A2(new_n635), .A3(new_n621), .ZN(new_n638));
  INV_X1    g213(.A(G14), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(KEYINPUT87), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT18), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n651), .B(new_n654), .Z(G227));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n657), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n666), .B(new_n667), .C1(new_n665), .C2(new_n664), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  INV_X1    g246(.A(G1981), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(new_n674), .ZN(G229));
  OAI21_X1  g250(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n676));
  INV_X1    g251(.A(G116), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(G2105), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n488), .B2(G128), .ZN(new_n679));
  INV_X1    g254(.A(G140), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n472), .A2(KEYINPUT90), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(KEYINPUT90), .B1(new_n472), .B2(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G29), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G26), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2067), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G1971), .Z(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(G6), .A2(G16), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n577), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n694), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT34), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n691), .A2(G24), .ZN(new_n706));
  INV_X1    g281(.A(G290), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n691), .ZN(new_n708));
  INV_X1    g283(.A(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n711));
  INV_X1    g286(.A(G107), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(new_n472), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G131), .ZN(new_n715));
  INV_X1    g290(.A(G119), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n487), .A2(KEYINPUT89), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT89), .B1(new_n487), .B2(new_n716), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G25), .B(new_n719), .S(G29), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  NAND3_X1  g297(.A1(new_n705), .A2(new_n710), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT36), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT24), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n686), .B1(new_n725), .B2(G34), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(KEYINPUT93), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G160), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n686), .ZN(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT94), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n593), .A2(new_n691), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G4), .B2(new_n691), .ZN(new_n737));
  INV_X1    g312(.A(G1348), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n542), .A2(new_n691), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n691), .B2(G19), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n743), .A2(G1341), .B1(new_n733), .B2(new_n732), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n739), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n743), .A2(G1341), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n691), .A2(KEYINPUT23), .A3(G20), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n748));
  INV_X1    g323(.A(G20), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G16), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n750), .C1(new_n558), .C2(new_n691), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1956), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n745), .A2(new_n746), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT29), .B(G2090), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G21), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G168), .B2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n757), .B1(G1966), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G5), .B2(G16), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n761), .A2(G5), .A3(G16), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n762), .B(new_n763), .C1(new_n535), .C2(new_n691), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n616), .A2(new_n617), .A3(new_n686), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G11), .Z(new_n768));
  AOI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n759), .C2(G1966), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  NOR2_X1   g345(.A1(G164), .A2(new_n686), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G27), .B2(new_n686), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n766), .B(new_n769), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n760), .B(new_n773), .C1(new_n770), .C2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n488), .A2(G129), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n714), .A2(G141), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n463), .A2(G105), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND4_X1  g354(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT95), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n686), .A2(G32), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT27), .B(G1996), .Z(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(KEYINPUT96), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(KEYINPUT96), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n786), .B(new_n787), .Z(new_n788));
  AND2_X1   g363(.A1(new_n686), .A2(G33), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT92), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT25), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n714), .A2(G139), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n501), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n792), .B(new_n793), .C1(new_n461), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(G2072), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n764), .A2(new_n765), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT30), .B(G28), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n798), .B(new_n799), .C1(new_n686), .C2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n753), .A2(new_n774), .A3(new_n788), .A4(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n724), .A2(new_n735), .A3(new_n803), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n690), .B(new_n804), .C1(new_n797), .C2(new_n796), .ZN(G311));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n690), .ZN(new_n806));
  INV_X1    g381(.A(new_n796), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(G2072), .B2(new_n807), .ZN(G150));
  NAND2_X1  g383(.A1(new_n509), .A2(G55), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT98), .B(G93), .Z(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n521), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n504), .A2(G67), .ZN(new_n812));
  NAND2_X1  g387(.A1(G80), .A2(G543), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n506), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n811), .A2(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n817), .A2(G860), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT101), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT100), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n817), .A2(new_n819), .ZN(new_n824));
  INV_X1    g399(.A(new_n542), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n818), .A2(new_n825), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n593), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n823), .B1(G860), .B2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n683), .B(G164), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(new_n607), .ZN(new_n836));
  INV_X1    g411(.A(G142), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n472), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n488), .A2(G130), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n461), .A2(G118), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n719), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n836), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n795), .A2(new_n780), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n781), .B2(new_n795), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(G160), .B(new_n618), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G162), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g429(.A1(G166), .A2(new_n696), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n516), .A2(G288), .ZN(new_n856));
  AOI21_X1  g431(.A(G305), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n855), .A2(new_n856), .A3(G305), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n707), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n861), .A2(new_n857), .A3(G290), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT42), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n829), .B(new_n601), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n593), .A2(G299), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n592), .A2(new_n558), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT103), .B1(new_n866), .B2(new_n867), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n867), .A2(KEYINPUT103), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n870), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n864), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G868), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(G868), .B2(new_n824), .ZN(G295));
  OAI21_X1  g455(.A(new_n879), .B1(G868), .B2(new_n824), .ZN(G331));
  AOI21_X1  g456(.A(G286), .B1(new_n560), .B2(new_n561), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n535), .A2(G168), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n826), .A2(new_n885), .A3(new_n828), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n542), .B1(new_n817), .B2(new_n819), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT104), .B1(new_n887), .B2(new_n827), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n886), .B(new_n888), .C1(new_n882), .C2(new_n883), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n890), .A2(new_n874), .A3(new_n875), .A4(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n868), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n863), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n860), .B2(new_n862), .ZN(new_n897));
  OAI21_X1  g472(.A(G290), .B1(new_n861), .B2(new_n857), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n858), .A2(new_n707), .A3(new_n859), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT105), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n890), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n869), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n872), .A2(new_n873), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n890), .A2(new_n904), .A3(KEYINPUT41), .A4(new_n891), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n895), .A2(new_n906), .A3(new_n907), .A4(new_n852), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT107), .ZN(new_n909));
  INV_X1    g484(.A(new_n894), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n892), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n911), .B2(new_n863), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n907), .A4(new_n906), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n901), .A2(new_n910), .A3(new_n892), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n895), .A2(new_n917), .A3(new_n852), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n918), .B2(KEYINPUT43), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n918), .A2(new_n916), .A3(KEYINPUT43), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n907), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n912), .A2(KEYINPUT43), .A3(new_n906), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  MUX2_X1   g499(.A(new_n921), .B(new_n924), .S(KEYINPUT44), .Z(G397));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(G164), .B2(G1384), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n714), .A2(G137), .B1(new_n463), .B2(G101), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(G40), .A3(new_n480), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n930), .B(KEYINPUT109), .Z(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n934), .B2(new_n781), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n934), .A2(new_n781), .A3(KEYINPUT108), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n683), .B(G2067), .Z(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(G1996), .B2(new_n780), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n935), .B(new_n936), .C1(new_n932), .C2(new_n939), .ZN(new_n940));
  OR3_X1    g515(.A1(new_n940), .A2(new_n721), .A3(new_n719), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n683), .A2(G2067), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n932), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n719), .B(new_n721), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT110), .Z(new_n945));
  NOR2_X1   g520(.A1(new_n932), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n709), .ZN(new_n948));
  INV_X1    g523(.A(new_n930), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT48), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n934), .B(KEYINPUT46), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n938), .A2(new_n780), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(new_n932), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  NOR3_X1   g531(.A1(new_n943), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n496), .A2(new_n502), .ZN(new_n958));
  INV_X1    g533(.A(new_n494), .ZN(new_n959));
  AOI21_X1  g534(.A(G1384), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT112), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n929), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n466), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n475), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(G138), .A3(new_n461), .A4(new_n468), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n967), .A2(KEYINPUT4), .B1(new_n500), .B2(new_n501), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n968), .B2(new_n494), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT50), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(new_n963), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n738), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n969), .A2(new_n929), .A3(G2067), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT118), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(KEYINPUT118), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT122), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n592), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n593), .A2(KEYINPUT122), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n980), .A2(KEYINPUT60), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT118), .B1(new_n973), .B2(new_n975), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n977), .B(new_n974), .C1(new_n972), .C2(new_n738), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT60), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(new_n981), .A3(new_n592), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT60), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1956), .ZN(new_n991));
  INV_X1    g566(.A(new_n929), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(KEYINPUT50), .B2(new_n969), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n960), .A2(new_n961), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n558), .A2(KEYINPUT57), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT57), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n555), .B2(new_n557), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT45), .B(new_n964), .C1(new_n968), .C2(new_n494), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT56), .B(G2072), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n927), .A2(new_n992), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n995), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n999), .B1(new_n995), .B2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(KEYINPUT119), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n1006), .B(new_n999), .C1(new_n995), .C2(new_n1002), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT61), .B(new_n1003), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1009));
  INV_X1    g584(.A(new_n1003), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n1004), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n927), .A2(new_n1000), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(KEYINPUT120), .A3(new_n933), .A4(new_n992), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n927), .A2(new_n992), .A3(new_n1000), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(G1996), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n969), .A2(new_n929), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT58), .B(G1341), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1014), .B(new_n1017), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n542), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT59), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n990), .A2(new_n1012), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n980), .A2(new_n592), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1003), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n972), .A2(G2090), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1016), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n927), .A2(KEYINPUT111), .A3(new_n992), .A4(new_n1000), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1028), .B(new_n1029), .C1(new_n1033), .C2(G1971), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n565), .B2(new_n566), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT55), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1971), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n972), .A2(G2090), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT113), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1034), .A2(new_n1037), .A3(new_n1040), .A4(G8), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1018), .A2(new_n1035), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n577), .A2(new_n672), .ZN(new_n1043));
  OAI21_X1  g618(.A(G1981), .B1(new_n574), .B2(new_n576), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n696), .A2(G1976), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1042), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1042), .A2(new_n1050), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1049), .B(new_n1053), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n993), .A2(new_n994), .A3(G2090), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1038), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1060), .B(new_n1035), .C1(new_n565), .C2(new_n566), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1056), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1041), .A2(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n960), .A2(KEYINPUT112), .A3(new_n961), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n970), .B1(new_n969), .B2(KEYINPUT50), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(KEYINPUT116), .A3(new_n733), .A4(new_n963), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n962), .A2(new_n963), .A3(new_n733), .A4(new_n971), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1966), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1016), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1068), .A2(new_n1071), .A3(G168), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT51), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1068), .A2(new_n1073), .A3(new_n1071), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(G286), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1076), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1031), .A2(new_n770), .A3(new_n1032), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n972), .A2(new_n765), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n473), .A2(KEYINPUT124), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n1088));
  AOI211_X1 g663(.A(new_n1087), .B(new_n481), .C1(new_n928), .C2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1013), .A2(G40), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1090));
  AND4_X1   g665(.A1(G301), .A2(new_n1084), .A3(new_n1085), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1082), .A2(new_n1083), .B1(new_n765), .B2(new_n972), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1016), .A2(new_n1087), .ZN(new_n1093));
  AOI21_X1  g668(.A(G301), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1081), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(G301), .A3(new_n1093), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1084), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1096), .B(KEYINPUT54), .C1(new_n1097), .C2(new_n535), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1064), .A2(new_n1080), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1027), .A2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n1056), .B(KEYINPUT114), .Z(new_n1102));
  INV_X1    g677(.A(new_n1041), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1049), .A2(new_n1051), .A3(new_n696), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1043), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT115), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1042), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G286), .A2(new_n1035), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1078), .A2(KEYINPUT117), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT117), .B1(new_n1078), .B2(new_n1110), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1041), .B(new_n1063), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1034), .A2(G8), .A3(new_n1040), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(new_n1062), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1078), .A2(new_n1110), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n1111), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1118), .A2(new_n1102), .A3(new_n1041), .A4(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1109), .B1(new_n1116), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1079), .A2(new_n1075), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1077), .B1(new_n1074), .B2(G8), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT62), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1076), .B(new_n1128), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(new_n1064), .A3(new_n1129), .A4(new_n1094), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1101), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(G290), .A2(G1986), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n949), .B1(new_n948), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n947), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT125), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1123), .A2(new_n1116), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1130), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1099), .B1(new_n1026), .B2(new_n1023), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT125), .B(new_n1134), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n957), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT126), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1144), .B(new_n957), .C1(new_n1135), .C2(new_n1141), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g721(.A(G227), .ZN(new_n1148));
  AND3_X1   g722(.A1(new_n853), .A2(new_n642), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g723(.A(new_n459), .ZN(new_n1150));
  INV_X1    g724(.A(G229), .ZN(new_n1151));
  NAND4_X1  g725(.A1(new_n921), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(G225));
  NAND2_X1  g726(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n1154), .A2(KEYINPUT106), .ZN(new_n1155));
  NAND3_X1  g729(.A1(new_n918), .A2(new_n916), .A3(KEYINPUT43), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g731(.A(new_n459), .B1(new_n1157), .B2(new_n915), .ZN(new_n1158));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n1159));
  NAND4_X1  g733(.A1(new_n1158), .A2(new_n1159), .A3(new_n1151), .A4(new_n1149), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1153), .A2(new_n1160), .ZN(G308));
endmodule


