//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n205));
  AOI21_X1  g004(.A(G36gat), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n202), .A2(new_n207), .A3(G29gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  OAI22_X1  g008(.A1(new_n206), .A2(new_n208), .B1(KEYINPUT15), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(G1gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n220), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n215), .A2(new_n217), .A3(new_n222), .A4(new_n218), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(KEYINPUT17), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n213), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n221), .A2(new_n223), .ZN(new_n228));
  INV_X1    g027(.A(new_n212), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT18), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT92), .B1(new_n224), .B2(new_n212), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n227), .B(KEYINPUT13), .Z(new_n237));
  NAND3_X1  g036(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT92), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n233), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n226), .A2(new_n227), .A3(new_n230), .A4(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(G197gat), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT11), .B(G169gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT12), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n234), .A2(new_n247), .A3(new_n239), .A4(new_n241), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G227gat), .ZN(new_n253));
  INV_X1    g052(.A(G233gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT23), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G169gat), .ZN(new_n263));
  INV_X1    g062(.A(G176gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n257), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(KEYINPUT68), .B2(KEYINPUT24), .ZN(new_n272));
  AND2_X1   g071(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n267), .B(new_n270), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n266), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n258), .A2(G169gat), .A3(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT23), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n278), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n256), .B1(new_n275), .B2(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n278), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT67), .B1(new_n281), .B2(new_n278), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(KEYINPUT69), .A3(new_n274), .A4(new_n266), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n279), .B1(new_n262), .B2(new_n265), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT64), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G183gat), .B2(G190gat), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n291), .A2(new_n292), .A3(new_n294), .A4(new_n267), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n264), .A2(KEYINPUT65), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n264), .A2(KEYINPUT65), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n296), .A2(KEYINPUT23), .A3(new_n263), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n289), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(new_n257), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n288), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G127gat), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n302), .A2(G134gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(G134gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n306));
  INV_X1    g105(.A(G120gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G113gat), .ZN(new_n308));
  INV_X1    g107(.A(G113gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G120gat), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n305), .B(new_n306), .C1(new_n311), .C2(KEYINPUT1), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT1), .B1(new_n308), .B2(new_n310), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n303), .B(new_n304), .C1(new_n313), .C2(KEYINPUT72), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n269), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n279), .B1(KEYINPUT26), .B2(new_n265), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n265), .A2(KEYINPUT26), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(G183gat), .B2(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n301), .A2(new_n315), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n315), .B1(new_n301), .B2(new_n326), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n255), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G15gat), .B(G43gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(G71gat), .B(G99gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT33), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n329), .A2(KEYINPUT32), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT73), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n329), .A2(new_n337), .A3(KEYINPUT32), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n332), .B1(new_n329), .B2(KEYINPUT32), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n329), .A2(new_n333), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n327), .A2(new_n328), .A3(new_n255), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n346));
  INV_X1    g145(.A(new_n344), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n347), .A3(new_n342), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n346), .ZN(new_n350));
  AOI221_X4 g149(.A(new_n344), .B1(new_n340), .B2(new_n341), .C1(new_n336), .C2(new_n338), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n347), .B1(new_n339), .B2(new_n342), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G148gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G141gat), .ZN(new_n356));
  INV_X1    g155(.A(G141gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G148gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  INV_X1    g159(.A(G155gat), .ZN(new_n361));
  INV_X1    g160(.A(G162gat), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT2), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G155gat), .B(G162gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n359), .A2(new_n365), .A3(new_n360), .A4(new_n363), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(KEYINPUT22), .B2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G211gat), .B(G218gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n369), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n367), .A2(new_n379), .A3(new_n368), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n376), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n380), .B1(KEYINPUT84), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n376), .B(KEYINPUT75), .Z(new_n391));
  NAND2_X1  g190(.A1(new_n381), .A2(new_n377), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n380), .A2(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT85), .B(G22gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n387), .A2(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT83), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n396), .A2(G22gat), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n400), .B2(new_n397), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n402), .A2(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT0), .ZN(new_n412));
  XNOR2_X1  g211(.A(G57gat), .B(G85gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT79), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n367), .A2(new_n368), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n417), .A2(KEYINPUT3), .B1(new_n314), .B2(new_n312), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n381), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n315), .A2(new_n369), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n314), .A2(new_n312), .A3(new_n367), .A4(new_n368), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT4), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n426));
  NAND2_X1  g225(.A1(new_n312), .A2(new_n314), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n417), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n422), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n429), .B2(new_n416), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(new_n423), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n315), .A2(new_n369), .A3(KEYINPUT81), .A4(new_n420), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n433), .A2(new_n419), .A3(new_n434), .A4(new_n426), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n414), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n414), .A3(new_n435), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n441), .A2(new_n438), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n442), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n437), .A2(KEYINPUT82), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n440), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT29), .B1(new_n301), .B2(new_n326), .ZN(new_n447));
  INV_X1    g246(.A(G226gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(new_n254), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT76), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n301), .B2(new_n326), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n301), .A2(new_n326), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n377), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n454), .B2(new_n451), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n376), .B(new_n450), .C1(new_n455), .C2(KEYINPUT76), .ZN(new_n456));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  NOR2_X1   g258(.A1(new_n447), .A2(new_n449), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n391), .B1(new_n460), .B2(new_n452), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT77), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n456), .A2(KEYINPUT77), .A3(new_n459), .A4(new_n461), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n459), .B1(new_n456), .B2(new_n461), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n456), .A2(new_n459), .A3(new_n461), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT30), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n446), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n354), .A2(new_n410), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT35), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n409), .B1(new_n349), .B2(new_n353), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT89), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n467), .A2(new_n470), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n439), .B1(new_n442), .B2(new_n437), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n475), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n446), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n409), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n349), .A2(new_n353), .A3(KEYINPUT36), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT36), .B1(new_n349), .B2(new_n353), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT40), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n418), .A2(new_n381), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n433), .A2(new_n492), .A3(new_n434), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n416), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n429), .A2(new_n416), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n494), .A2(KEYINPUT39), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n414), .B1(new_n494), .B2(KEYINPUT39), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n437), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n496), .A2(new_n497), .A3(new_n491), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n464), .A2(new_n466), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n456), .A2(new_n461), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n459), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n456), .B2(new_n461), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT76), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n460), .B2(new_n452), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n376), .B1(new_n514), .B2(new_n450), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n460), .A2(new_n452), .A3(new_n391), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT37), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n517), .A2(new_n504), .A3(new_n508), .A4(new_n507), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n503), .A2(new_n512), .A3(new_n518), .A4(new_n482), .ZN(new_n519));
  AND4_X1   g318(.A1(KEYINPUT88), .A2(new_n502), .A3(new_n519), .A4(new_n410), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n409), .B1(new_n480), .B2(new_n501), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT88), .B1(new_n521), .B2(new_n519), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n487), .B(new_n490), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n252), .B1(new_n485), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT93), .ZN(new_n526));
  AND2_X1   g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  OAI22_X1  g327(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G57gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G64gat), .ZN(new_n531));
  INV_X1    g330(.A(G64gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G57gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n525), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n529), .B(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT21), .ZN(new_n536));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G127gat), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n228), .B1(KEYINPUT21), .B2(new_n535), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(new_n361), .ZN(new_n543));
  XOR2_X1   g342(.A(G183gat), .B(G211gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n541), .A2(new_n546), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  XOR2_X1   g350(.A(G99gat), .B(G106gat), .Z(new_n552));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  INV_X1    g352(.A(G85gat), .ZN(new_n554));
  INV_X1    g353(.A(G92gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(KEYINPUT8), .A2(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n552), .B1(new_n551), .B2(new_n556), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  OR3_X1    g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n213), .A2(new_n225), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n563), .B(new_n564), .C1(new_n212), .C2(new_n562), .ZN(new_n565));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566));
  OR2_X1    g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n566), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n567), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576));
  INV_X1    g375(.A(G230gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n254), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n535), .A2(KEYINPUT10), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n560), .A3(new_n561), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT96), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n579), .A2(new_n560), .A3(new_n582), .A4(new_n561), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n551), .A2(new_n556), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT95), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n535), .A2(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n557), .A2(new_n558), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n578), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n578), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n576), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n524), .A2(new_n549), .A3(new_n575), .A4(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n486), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G1gat), .ZN(G1324gat));
  INV_X1    g405(.A(KEYINPUT42), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n603), .A2(new_n481), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT16), .B(G8gat), .Z(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(G8gat), .B1(new_n603), .B2(new_n481), .ZN(new_n611));
  NOR2_X1   g410(.A1(KEYINPUT98), .A2(KEYINPUT42), .ZN(new_n612));
  MUX2_X1   g411(.A(KEYINPUT98), .B(new_n612), .S(new_n609), .Z(new_n613));
  AOI22_X1  g412(.A1(new_n610), .A2(new_n611), .B1(new_n608), .B2(new_n613), .ZN(G1325gat));
  INV_X1    g413(.A(G15gat), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n603), .A2(new_n615), .A3(new_n490), .ZN(new_n616));
  INV_X1    g415(.A(new_n354), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n603), .B2(new_n617), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT99), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(KEYINPUT99), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(G1326gat));
  OR3_X1    g420(.A1(new_n603), .A2(KEYINPUT100), .A3(new_n410), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT100), .B1(new_n603), .B2(new_n410), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT43), .B(G22gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(G1327gat));
  INV_X1    g425(.A(new_n602), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n549), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n574), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT101), .Z(new_n630));
  AND2_X1   g429(.A1(new_n524), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(new_n203), .A3(new_n486), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT45), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n251), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n484), .B1(new_n478), .B2(KEYINPUT89), .ZN(new_n635));
  AOI211_X1 g434(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n471), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n523), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT102), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n485), .A2(new_n639), .A3(new_n523), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n574), .B(KEYINPUT103), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT44), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n574), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT44), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n634), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(G29gat), .B1(new_n648), .B2(new_n446), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n649), .ZN(G1328gat));
  NAND3_X1  g449(.A1(new_n631), .A2(new_n207), .A3(new_n480), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT46), .Z(new_n652));
  OAI21_X1  g451(.A(G36gat), .B1(new_n648), .B2(new_n481), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(G1329gat));
  NOR2_X1   g453(.A1(new_n617), .A2(G43gat), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n637), .A2(new_n630), .A3(new_n251), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT104), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n524), .A2(new_n658), .A3(new_n630), .A4(new_n655), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT105), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n657), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(G43gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n490), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n647), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n660), .A2(KEYINPUT47), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n668), .A2(KEYINPUT47), .B1(new_n667), .B2(new_n669), .ZN(G1330gat));
  NAND2_X1  g469(.A1(new_n631), .A2(new_n409), .ZN(new_n671));
  INV_X1    g470(.A(G50gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n409), .A2(G50gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n648), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT48), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n677), .B(new_n673), .C1(new_n648), .C2(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(G1331gat));
  AND2_X1   g478(.A1(new_n638), .A2(new_n640), .ZN(new_n680));
  INV_X1    g479(.A(new_n549), .ZN(new_n681));
  NOR4_X1   g480(.A1(new_n681), .A2(new_n251), .A3(new_n574), .A4(new_n602), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n446), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n530), .ZN(G1332gat));
  NOR2_X1   g485(.A1(new_n684), .A2(new_n481), .ZN(new_n687));
  NOR2_X1   g486(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n688));
  AND2_X1   g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n687), .B2(new_n688), .ZN(G1333gat));
  AND2_X1   g490(.A1(new_n680), .A2(new_n683), .ZN(new_n692));
  INV_X1    g491(.A(G71gat), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n354), .ZN(new_n694));
  OAI21_X1  g493(.A(G71gat), .B1(new_n684), .B2(new_n490), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT50), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n694), .A2(KEYINPUT50), .A3(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1334gat));
  NAND2_X1  g499(.A1(new_n692), .A2(new_n409), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g501(.A(new_n575), .B1(new_n485), .B2(new_n523), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n549), .A2(new_n251), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n703), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n704), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n637), .A2(new_n574), .A3(new_n704), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n707), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n712), .A2(new_n554), .A3(new_n486), .A4(new_n627), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n704), .A2(new_n627), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n644), .B2(new_n646), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(new_n486), .ZN(new_n716));
  OAI21_X1  g515(.A(G85gat), .B1(new_n716), .B2(KEYINPUT107), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n486), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(G1336gat));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n481), .A2(G92gat), .A3(new_n602), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n712), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n715), .A2(new_n480), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n720), .B(new_n722), .C1(new_n723), .C2(new_n555), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n555), .B1(new_n715), .B2(new_n480), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n705), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT110), .B1(new_n728), .B2(new_n721), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n730));
  INV_X1    g529(.A(new_n721), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n730), .B(new_n731), .C1(new_n727), .C2(new_n705), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n725), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n724), .B1(new_n733), .B2(new_n720), .ZN(G1337gat));
  INV_X1    g533(.A(new_n715), .ZN(new_n735));
  OAI21_X1  g534(.A(G99gat), .B1(new_n735), .B2(new_n490), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n617), .A2(G99gat), .A3(new_n602), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n712), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(G1338gat));
  INV_X1    g538(.A(G106gat), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n715), .B2(new_n409), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n410), .A2(new_n602), .A3(G106gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n712), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n728), .A2(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT53), .B1(new_n741), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1339gat));
  AOI21_X1  g548(.A(new_n227), .B1(new_n226), .B2(new_n230), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n237), .B1(new_n236), .B2(new_n238), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n246), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT111), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n754), .B(new_n246), .C1(new_n750), .C2(new_n751), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n753), .A2(new_n250), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n600), .A3(new_n601), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(KEYINPUT112), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n598), .B1(new_n592), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n584), .A2(new_n591), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n593), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n593), .B1(new_n589), .B2(new_n590), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n764), .B2(new_n584), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n592), .A2(new_n594), .A3(new_n599), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n763), .B2(new_n765), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n761), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n251), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n759), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n642), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n641), .A2(new_n756), .A3(new_n772), .A4(new_n769), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n549), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n549), .A2(new_n575), .A3(new_n252), .A4(new_n602), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n481), .A2(new_n486), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n617), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n410), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n780), .A2(KEYINPUT113), .A3(new_n410), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G113gat), .B1(new_n787), .B2(new_n252), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n780), .A2(new_n486), .ZN(new_n789));
  INV_X1    g588(.A(new_n477), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n480), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n251), .A2(new_n309), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT114), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n788), .A2(new_n795), .ZN(G1340gat));
  NOR3_X1   g595(.A1(new_n787), .A2(new_n307), .A3(new_n602), .ZN(new_n797));
  AOI21_X1  g596(.A(G120gat), .B1(new_n792), .B2(new_n627), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(G1341gat));
  NAND3_X1  g598(.A1(new_n785), .A2(new_n549), .A3(new_n786), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G127gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n792), .A2(new_n302), .A3(new_n549), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(new_n802), .A3(KEYINPUT115), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1342gat));
  AOI211_X1 g606(.A(G134gat), .B(new_n575), .C1(KEYINPUT116), .C2(KEYINPUT56), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n789), .A2(new_n791), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G134gat), .B1(new_n787), .B2(new_n575), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1343gat));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n780), .A2(new_n814), .A3(new_n409), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n666), .A2(new_n781), .ZN(new_n816));
  XOR2_X1   g615(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n817));
  NAND2_X1  g616(.A1(new_n767), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n251), .A2(new_n818), .A3(new_n772), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n757), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n776), .B1(new_n574), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n779), .B1(new_n821), .B2(new_n681), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT57), .B1(new_n822), .B2(new_n410), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n815), .A2(new_n816), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G141gat), .B1(new_n824), .B2(new_n252), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n666), .A2(new_n480), .A3(new_n410), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n789), .A2(new_n826), .A3(new_n357), .A4(new_n251), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n828), .B(new_n831), .ZN(G1344gat));
  NOR3_X1   g631(.A1(new_n824), .A2(KEYINPUT59), .A3(new_n602), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n789), .A2(new_n826), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT59), .B1(new_n834), .B2(new_n602), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n355), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT57), .B(new_n409), .C1(new_n777), .C2(new_n779), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n574), .B1(new_n757), .B2(new_n819), .ZN(new_n838));
  AND4_X1   g637(.A1(new_n574), .A2(new_n756), .A3(new_n772), .A4(new_n769), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n681), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n778), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n410), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(KEYINPUT119), .A3(new_n778), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT57), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n837), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g646(.A(KEYINPUT120), .B(KEYINPUT57), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR4_X1   g648(.A1(new_n849), .A2(new_n666), .A3(new_n602), .A4(new_n781), .ZN(new_n850));
  NAND2_X1  g649(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n836), .B1(new_n850), .B2(new_n851), .ZN(G1345gat));
  OAI21_X1  g651(.A(G155gat), .B1(new_n824), .B2(new_n681), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n549), .A2(new_n361), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n834), .B2(new_n854), .ZN(G1346gat));
  NOR3_X1   g654(.A1(new_n824), .A2(new_n362), .A3(new_n642), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n789), .A2(new_n574), .A3(new_n826), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n362), .B2(new_n857), .ZN(G1347gat));
  NOR2_X1   g657(.A1(new_n790), .A2(new_n481), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT121), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n780), .A2(new_n446), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n252), .A2(G169gat), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n861), .A2(KEYINPUT122), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT122), .B1(new_n861), .B2(new_n863), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n481), .A2(new_n486), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n780), .A2(new_n410), .A3(new_n354), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G169gat), .B1(new_n868), .B2(new_n252), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n866), .A2(KEYINPUT123), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1348gat));
  AOI211_X1 g673(.A(new_n602), .B(new_n868), .C1(new_n297), .C2(new_n296), .ZN(new_n875));
  INV_X1    g674(.A(new_n861), .ZN(new_n876));
  AOI21_X1  g675(.A(G176gat), .B1(new_n876), .B2(new_n627), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(G1349gat));
  OAI21_X1  g677(.A(G183gat), .B1(new_n868), .B2(new_n681), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n549), .A2(new_n316), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n861), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n876), .A2(new_n269), .A3(new_n641), .ZN(new_n883));
  OAI21_X1  g682(.A(G190gat), .B1(new_n868), .B2(new_n575), .ZN(new_n884));
  XOR2_X1   g683(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(G1351gat));
  AND2_X1   g687(.A1(new_n780), .A2(new_n446), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n666), .A2(new_n481), .A3(new_n410), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G197gat), .B1(new_n893), .B2(new_n251), .ZN(new_n894));
  INV_X1    g693(.A(new_n849), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n490), .A2(new_n867), .ZN(new_n896));
  XOR2_X1   g695(.A(new_n896), .B(KEYINPUT126), .Z(new_n897));
  AND2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n251), .A2(G197gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n602), .A2(G204gat), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n889), .A2(new_n891), .A3(new_n892), .A4(new_n901), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT62), .Z(new_n903));
  NAND3_X1  g702(.A1(new_n895), .A2(new_n627), .A3(new_n897), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G204gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1353gat));
  NAND3_X1  g705(.A1(new_n893), .A2(new_n371), .A3(new_n549), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n549), .B(new_n897), .C1(new_n847), .C2(new_n848), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G211gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n909), .A2(new_n910), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(G1354gat));
  NAND3_X1  g714(.A1(new_n895), .A2(new_n574), .A3(new_n897), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G218gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n372), .A3(new_n641), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1355gat));
endmodule


