//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n202), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n207), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n219), .A2(new_n220), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n220), .B2(new_n219), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n217), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G68), .Z(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n226), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT74), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G58), .A2(G68), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n227), .B1(new_n223), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G159), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n252), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n253), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n259), .B2(new_n201), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(KEYINPUT74), .A3(new_n256), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT7), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n222), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n251), .B1(new_n273), .B2(KEYINPUT16), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT75), .B1(new_n268), .B2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT75), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(new_n266), .A3(KEYINPUT3), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n278), .A3(new_n269), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n263), .A2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n222), .B1(new_n281), .B2(new_n265), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n275), .B1(new_n282), .B2(new_n262), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n250), .B1(new_n284), .B2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT8), .A2(G58), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT8), .A2(G58), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n284), .A2(G13), .A3(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n274), .A2(new_n283), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n267), .A2(new_n269), .A3(G226), .A4(G1698), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n267), .A2(new_n269), .A3(G223), .A4(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n295), .B(new_n297), .C1(new_n266), .C2(new_n210), .ZN(new_n298));
  AND2_X1   g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(new_n226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  INV_X1    g0102(.A(G45), .ZN(new_n303));
  AOI21_X1  g0103(.A(G1), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n304), .A2(G274), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G1), .A3(G13), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n284), .B1(G41), .B2(G45), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n305), .B1(new_n310), .B2(G232), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n301), .A2(G190), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n301), .B2(new_n311), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n294), .A2(KEYINPUT76), .A3(KEYINPUT17), .A4(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n270), .B2(new_n227), .ZN(new_n317));
  AOI211_X1 g0117(.A(new_n263), .B(G20), .C1(new_n267), .C2(new_n269), .ZN(new_n318));
  OAI21_X1  g0118(.A(G68), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n319), .A2(KEYINPUT16), .A3(new_n258), .A4(new_n261), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n283), .A2(new_n320), .A3(new_n250), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n290), .A2(new_n293), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n315), .A2(new_n321), .A3(KEYINPUT76), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT17), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n301), .A2(new_n311), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G169), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n301), .A2(G179), .A3(new_n311), .ZN(new_n329));
  AOI221_X4 g0129(.A(new_n326), .B1(new_n328), .B2(new_n329), .C1(new_n321), .C2(new_n322), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n321), .A2(new_n322), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n329), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT18), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n316), .B(new_n325), .C1(new_n330), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT77), .ZN(new_n335));
  INV_X1    g0135(.A(new_n332), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n326), .B1(new_n294), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(KEYINPUT18), .A3(new_n332), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT77), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n339), .A2(new_n340), .A3(new_n316), .A4(new_n325), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n305), .B1(new_n310), .B2(G238), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n267), .A2(new_n269), .A3(G232), .A4(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n267), .A2(new_n269), .A3(G226), .A4(new_n296), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G97), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n347), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT71), .B1(new_n347), .B2(new_n300), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n343), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n266), .A2(G20), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(G77), .B1(G20), .B2(new_n222), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n227), .A2(new_n266), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n202), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g0159(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n360));
  AND3_X1   g0160(.A1(new_n359), .A2(new_n250), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n292), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT12), .A3(new_n222), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT12), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n292), .B2(G68), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n363), .B(new_n365), .C1(new_n286), .C2(new_n222), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n360), .B1(new_n359), .B2(new_n250), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n355), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT72), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n351), .A2(new_n371), .A3(new_n353), .ZN(new_n372));
  OR3_X1    g0172(.A1(new_n350), .A2(new_n371), .A3(KEYINPUT13), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n354), .A2(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT14), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT14), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n354), .A2(new_n378), .A3(G169), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n372), .A2(new_n373), .ZN(new_n380));
  INV_X1    g0180(.A(G179), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n377), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n368), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n342), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n304), .A2(G274), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n309), .B2(new_n209), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n268), .A2(G33), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n389));
  OAI21_X1  g0189(.A(G77), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n267), .A2(new_n269), .A3(G222), .A4(new_n296), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n267), .A2(new_n269), .A3(G223), .A4(G1698), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n387), .B1(new_n300), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT69), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(G190), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n300), .ZN(new_n397));
  INV_X1    g0197(.A(new_n387), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(G190), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT69), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n394), .A2(new_n313), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT68), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT67), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT9), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n284), .A2(G20), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(new_n249), .A3(G50), .A4(new_n226), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G50), .B2(new_n292), .ZN(new_n409));
  OAI21_X1  g0209(.A(G20), .B1(new_n223), .B2(G50), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n255), .A2(G150), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n227), .A2(G33), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(new_n291), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n409), .B1(new_n413), .B2(new_n250), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n404), .A2(new_n405), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n406), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n289), .A2(new_n356), .B1(G150), .B2(new_n255), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n251), .B1(new_n417), .B2(new_n410), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n404), .B(new_n405), .C1(new_n418), .C2(new_n409), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n402), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT10), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n403), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n402), .B(new_n420), .C1(KEYINPUT68), .C2(KEYINPUT10), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n394), .A2(G169), .B1(new_n418), .B2(new_n409), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n394), .A2(new_n381), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n289), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n412), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n250), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n285), .A2(G77), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n362), .A2(new_n203), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n264), .A2(G232), .A3(new_n296), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n264), .A2(G238), .A3(G1698), .ZN(new_n437));
  INV_X1    g0237(.A(G107), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(new_n264), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n300), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n305), .B1(new_n310), .B2(G244), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n435), .B1(new_n442), .B2(G200), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(G190), .A3(new_n441), .ZN(new_n444));
  INV_X1    g0244(.A(G169), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n442), .A2(new_n445), .B1(new_n431), .B2(new_n434), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n440), .A2(new_n381), .A3(new_n441), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n443), .A2(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n423), .A2(new_n424), .A3(new_n427), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT70), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n449), .B(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT78), .B1(new_n385), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n449), .B(KEYINPUT70), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT78), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n384), .A4(new_n342), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n267), .A2(new_n269), .A3(G257), .A4(new_n296), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT86), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n264), .A2(KEYINPUT86), .A3(G257), .A4(new_n296), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n264), .A2(G264), .A3(G1698), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n270), .A2(G303), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n300), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT82), .B1(new_n465), .B2(G41), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT82), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(new_n302), .A3(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n284), .B(G45), .C1(new_n302), .C2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n300), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n466), .B2(new_n468), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n472), .A2(G270), .B1(G274), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT84), .A2(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT84), .A2(G116), .ZN(new_n477));
  OAI21_X1  g0277(.A(G20), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  INV_X1    g0279(.A(G97), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n227), .C1(G33), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n250), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT20), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n478), .A2(KEYINPUT20), .A3(new_n250), .A4(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n292), .B1(G1), .B2(new_n266), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n250), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n476), .A2(new_n477), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n488), .A2(G116), .B1(new_n362), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n445), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n475), .A2(new_n492), .A3(KEYINPUT21), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n464), .A2(new_n474), .A3(G179), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n486), .A2(new_n491), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT21), .B1(new_n475), .B2(new_n492), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n494), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n475), .A2(G200), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n497), .C1(new_n370), .C2(new_n475), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT87), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n362), .A2(KEYINPUT25), .A3(new_n438), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT25), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n292), .B2(G107), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n488), .A2(G107), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(KEYINPUT84), .A2(G116), .ZN(new_n508));
  NAND2_X1  g0308(.A1(KEYINPUT84), .A2(G116), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n356), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n227), .B2(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n438), .A2(KEYINPUT23), .A3(G20), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n267), .A2(new_n269), .A3(new_n227), .A4(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n264), .A2(new_n518), .A3(new_n227), .A4(G87), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n515), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n250), .B1(new_n520), .B2(KEYINPUT24), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  AOI211_X1 g0322(.A(new_n522), .B(new_n515), .C1(new_n517), .C2(new_n519), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n507), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n267), .A2(new_n269), .A3(G250), .A4(new_n296), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n267), .A2(new_n269), .A3(G257), .A4(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G294), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n300), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n473), .A2(G274), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n466), .A2(new_n468), .ZN(new_n531));
  OAI211_X1 g0331(.A(G264), .B(new_n307), .C1(new_n531), .C2(new_n470), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G169), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n529), .A2(new_n532), .A3(G179), .A4(new_n530), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n503), .B1(new_n524), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n524), .A2(new_n536), .A3(new_n503), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n500), .B(new_n502), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n533), .A2(G200), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n529), .A2(new_n532), .A3(G190), .A4(new_n530), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n524), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n267), .A2(new_n269), .A3(G244), .A4(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n267), .A2(new_n269), .A3(G238), .A4(new_n296), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n508), .A2(G33), .A3(new_n509), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n300), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n303), .A2(G1), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G274), .ZN(new_n550));
  OAI21_X1  g0350(.A(G250), .B1(new_n303), .B2(G1), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n300), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  INV_X1    g0355(.A(new_n429), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n292), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n412), .B2(new_n480), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT85), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n267), .A2(new_n269), .A3(new_n227), .A4(G68), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT85), .B(new_n558), .C1(new_n412), .C2(new_n480), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n227), .B1(new_n346), .B2(new_n558), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G97), .A2(G107), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n210), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n568), .B2(new_n250), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n552), .B1(new_n547), .B2(new_n300), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G190), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n488), .A2(G87), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n555), .A2(new_n569), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n554), .A2(new_n445), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT19), .B1(new_n356), .B2(G97), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n567), .B1(new_n575), .B2(KEYINPUT85), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n563), .A2(new_n562), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n250), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n488), .A2(new_n556), .ZN(new_n579));
  INV_X1    g0379(.A(new_n557), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n570), .A2(new_n381), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n574), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n573), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n543), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n472), .A2(G257), .B1(G274), .B2(new_n473), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n267), .A2(new_n269), .A3(G244), .A4(new_n296), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n264), .A2(G250), .A3(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n479), .A4(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n592), .A2(KEYINPUT81), .A3(new_n300), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT81), .B1(new_n592), .B2(new_n300), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n292), .A2(G97), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n488), .B2(G97), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(G97), .A2(G107), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n565), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n605), .A3(KEYINPUT80), .ZN(new_n606));
  AND2_X1   g0406(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT80), .B1(new_n607), .B2(new_n600), .ZN(new_n608));
  XNOR2_X1  g0408(.A(G97), .B(G107), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n601), .A2(new_n480), .A3(new_n602), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n606), .A2(new_n610), .A3(G20), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n255), .A2(G77), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n270), .A2(new_n227), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(new_n263), .B1(new_n279), .B2(new_n280), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(new_n613), .C1(new_n615), .C2(new_n438), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n599), .B1(new_n616), .B2(new_n250), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n592), .A2(new_n300), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n586), .A3(KEYINPUT83), .A4(G190), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n586), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n370), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n596), .A2(new_n617), .A3(new_n619), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n616), .A2(new_n250), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n598), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n381), .B(new_n586), .C1(new_n593), .C2(new_n594), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n445), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n585), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n539), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n456), .A2(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n427), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n382), .A2(new_n383), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n446), .A2(new_n447), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT90), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n375), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n316), .B(new_n325), .C1(new_n633), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n339), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n423), .A2(new_n424), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n632), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n456), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n524), .A2(new_n536), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n475), .A2(new_n492), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT21), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n464), .A2(new_n474), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(G179), .A3(new_n496), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n642), .A2(new_n645), .A3(new_n647), .A4(new_n493), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n623), .A2(new_n585), .A3(new_n648), .A4(new_n628), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT88), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n622), .A2(new_n617), .A3(new_n619), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n624), .A2(new_n598), .B1(new_n621), .B2(new_n445), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n651), .A2(new_n596), .B1(new_n626), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT88), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n585), .A4(new_n648), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n628), .B2(new_n584), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n578), .A2(new_n580), .A3(new_n572), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n570), .A2(new_n313), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(G169), .B1(new_n548), .B2(new_n553), .ZN(new_n663));
  AOI211_X1 g0463(.A(G179), .B(new_n552), .C1(new_n547), .C2(new_n300), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n662), .A2(new_n571), .B1(new_n665), .B2(new_n581), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .A3(new_n626), .A4(new_n652), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n657), .B1(new_n668), .B2(new_n583), .ZN(new_n669));
  INV_X1    g0469(.A(new_n583), .ZN(new_n670));
  AOI211_X1 g0470(.A(KEYINPUT89), .B(new_n670), .C1(new_n659), .C2(new_n667), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n656), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n640), .B1(new_n641), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g0473(.A(new_n673), .B(KEYINPUT91), .Z(G369));
  NAND3_X1  g0474(.A1(new_n284), .A2(new_n227), .A3(G13), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT92), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n675), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n681), .A3(G213), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G343), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT94), .B1(new_n688), .B2(new_n497), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n502), .A2(new_n645), .A3(new_n647), .A4(new_n493), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND4_X1   g0493(.A1(G343), .A2(new_n524), .A3(new_n685), .A4(new_n684), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n694), .A2(new_n538), .A3(new_n537), .ZN(new_n695));
  INV_X1    g0495(.A(new_n536), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n543), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT95), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT95), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n695), .A2(new_n700), .A3(new_n697), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n686), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n500), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n699), .B2(new_n701), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n705), .A2(new_n642), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n703), .A2(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n218), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n566), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n224), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n672), .B2(new_n705), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n538), .A2(new_n537), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n500), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n585), .A2(new_n623), .A3(new_n628), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n670), .B1(new_n659), .B2(new_n667), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n705), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n720), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n721), .A2(new_n690), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n724), .A2(new_n732), .A3(new_n688), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n495), .A2(new_n621), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n529), .A2(new_n532), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n570), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT96), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT96), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n570), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND4_X1   g0542(.A1(new_n381), .A2(new_n475), .A3(new_n533), .A4(new_n554), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n740), .A2(new_n741), .B1(new_n595), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n705), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n731), .B1(new_n733), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n688), .B1(new_n742), .B2(new_n744), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(KEYINPUT31), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n692), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n730), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n718), .B1(new_n752), .B2(G1), .ZN(G364));
  AND2_X1   g0553(.A1(new_n227), .A2(G13), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n284), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n713), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OR3_X1    g0560(.A1(new_n760), .A2(KEYINPUT97), .A3(G20), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT97), .B1(new_n760), .B2(G20), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n226), .B1(G20), .B2(new_n445), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT98), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n712), .A2(new_n270), .ZN(new_n767));
  INV_X1    g0567(.A(G116), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n767), .A2(G355), .B1(new_n768), .B2(new_n712), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n247), .A2(new_n303), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n712), .A2(new_n264), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G45), .B2(new_n224), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n758), .B1(new_n766), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT99), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n227), .A2(new_n370), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n381), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n381), .A2(new_n313), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n776), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n227), .A2(G190), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(G179), .A3(new_n313), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n264), .B(new_n782), .C1(G311), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n783), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n787), .A2(G179), .A3(new_n313), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n788), .A2(G283), .B1(G329), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n776), .A2(G179), .A3(new_n313), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n779), .A2(new_n783), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(G322), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n227), .B1(new_n789), .B2(G190), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G294), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n786), .A2(new_n792), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n788), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n438), .ZN(new_n804));
  INV_X1    g0604(.A(new_n777), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n270), .B(new_n804), .C1(G87), .C2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT100), .Z(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n790), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n800), .A2(G97), .ZN(new_n811));
  INV_X1    g0611(.A(new_n780), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n794), .A2(G58), .B1(new_n812), .B2(G50), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n785), .A2(G77), .B1(new_n796), .B2(G68), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n810), .A2(new_n811), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n802), .B1(new_n807), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n816), .A2(new_n764), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n775), .B(new_n817), .C1(new_n691), .C2(new_n763), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n693), .A2(new_n757), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n691), .A2(new_n692), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  INV_X1    g0622(.A(KEYINPUT101), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n705), .A2(new_n435), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n635), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n824), .A2(new_n448), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n672), .B2(new_n705), .ZN(new_n828));
  INV_X1    g0628(.A(new_n827), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n668), .A2(new_n583), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT89), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n726), .A2(new_n657), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n688), .B(new_n829), .C1(new_n833), .C2(new_n656), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n751), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n823), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n757), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n751), .A2(new_n828), .A3(KEYINPUT101), .A4(new_n834), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n764), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n760), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n757), .B1(new_n842), .B2(G77), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n264), .B1(new_n777), .B2(new_n202), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n803), .A2(new_n222), .B1(new_n790), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(G58), .C2(new_n800), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n812), .A2(G137), .B1(new_n785), .B2(G159), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n794), .A2(G143), .B1(new_n796), .B2(G150), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n850), .A2(KEYINPUT34), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n847), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(G311), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n777), .A2(new_n438), .B1(new_n790), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n264), .B(new_n855), .C1(new_n489), .C2(new_n785), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n788), .A2(G87), .B1(new_n812), .B2(G303), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n794), .A2(G294), .B1(new_n796), .B2(G283), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n856), .A2(new_n811), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n843), .B1(new_n860), .B2(new_n764), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n829), .B2(new_n760), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n840), .A2(new_n862), .ZN(G384));
  NAND3_X1  g0663(.A1(new_n606), .A2(new_n610), .A3(new_n611), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(G116), .A3(new_n228), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  NOR3_X1   g0669(.A1(new_n224), .A2(new_n203), .A3(new_n259), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n202), .B2(G68), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n284), .B(G13), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n339), .A2(new_n687), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n687), .A2(new_n331), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n294), .A2(new_n315), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n331), .A2(new_n332), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n273), .B1(new_n882), .B2(KEYINPUT16), .ZN(new_n883));
  OAI211_X1 g0683(.A(KEYINPUT105), .B(new_n275), .C1(new_n262), .C2(new_n272), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n250), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n322), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n886), .A2(new_n687), .B1(new_n294), .B2(new_n315), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n332), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT106), .B(new_n881), .C1(new_n889), .C2(new_n879), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n892));
  INV_X1    g0692(.A(new_n881), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n334), .A2(new_n687), .A3(new_n886), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT38), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT39), .ZN(new_n901));
  INV_X1    g0701(.A(new_n877), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n334), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n903), .A2(KEYINPUT108), .B1(new_n893), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n903), .A2(KEYINPUT108), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n897), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n899), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n901), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n633), .A2(new_n688), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT107), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n876), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n669), .A2(new_n671), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n650), .A2(new_n655), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n705), .B(new_n827), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n705), .A2(new_n634), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT103), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n916), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n921), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n834), .A2(KEYINPUT104), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n705), .A2(new_n383), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n384), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n382), .A2(new_n383), .A3(new_n705), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n929), .A3(new_n900), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n915), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT110), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n456), .A2(new_n720), .A3(new_n728), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n933), .A2(new_n640), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n932), .B(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n829), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(new_n750), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n898), .A2(new_n938), .A3(new_n899), .ZN(new_n939));
  NAND2_X1  g0739(.A1(KEYINPUT109), .A2(KEYINPUT40), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n749), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n748), .B1(new_n630), .B2(new_n688), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n731), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n829), .A3(new_n929), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n945), .A2(KEYINPUT109), .B1(new_n908), .B2(new_n899), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n941), .B1(new_n946), .B2(new_n938), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(G330), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n456), .A2(new_n751), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n641), .A2(new_n750), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n948), .A2(new_n949), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n935), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n284), .B2(new_n754), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n935), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n875), .B1(new_n953), .B2(new_n954), .ZN(G367));
  OAI211_X1 g0755(.A(new_n623), .B(new_n628), .C1(new_n688), .C2(new_n617), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT112), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n705), .A2(new_n626), .A3(new_n652), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n701), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n700), .B1(new_n695), .B2(new_n697), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n706), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n960), .A2(KEYINPUT42), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n628), .B1(new_n957), .B2(new_n722), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n688), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT42), .B1(new_n960), .B2(new_n963), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n705), .A2(new_n660), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n666), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n583), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT111), .Z(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n703), .A2(new_n960), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n973), .A2(new_n975), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n978), .ZN(new_n981));
  INV_X1    g0781(.A(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n981), .B1(new_n982), .B2(new_n976), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n713), .B(KEYINPUT41), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n710), .B2(new_n959), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n960), .B(KEYINPUT44), .C1(new_n708), .C2(new_n709), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n710), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n990));
  INV_X1    g0790(.A(new_n709), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n963), .A2(new_n959), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n703), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n989), .A2(new_n995), .A3(new_n703), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n702), .A2(new_n706), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(new_n693), .A3(new_n963), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1000), .A2(new_n708), .B1(new_n692), .B2(new_n691), .ZN(new_n1003));
  AND4_X1   g0803(.A1(new_n836), .A2(new_n1002), .A3(new_n729), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n999), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n985), .B1(new_n1005), .B2(new_n752), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n980), .B(new_n983), .C1(new_n1006), .C2(new_n756), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n765), .B1(new_n218), .B2(new_n429), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n771), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n239), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n757), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n788), .A2(G77), .ZN(new_n1012));
  INV_X1    g0812(.A(G137), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(new_n790), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n270), .B(new_n1014), .C1(G58), .C2(new_n805), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G150), .A2(new_n794), .B1(new_n785), .B2(G50), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G143), .A2(new_n812), .B1(new_n796), .B2(G159), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n799), .A2(new_n222), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n793), .A2(new_n778), .B1(new_n780), .B2(new_n854), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT113), .Z(new_n1022));
  NOR3_X1   g0822(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n490), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n805), .A2(G116), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1023), .B1(KEYINPUT46), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n796), .A2(G294), .ZN(new_n1026));
  INV_X1    g0826(.A(G317), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n790), .C1(new_n803), .C2(new_n480), .ZN(new_n1028));
  INV_X1    g0828(.A(G283), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n270), .B1(new_n799), .B2(new_n438), .C1(new_n784), .C2(new_n1029), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n1022), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT47), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n841), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1011), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n763), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n971), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1007), .A2(new_n1038), .ZN(G387));
  AND2_X1   g0839(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n756), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n270), .B1(new_n781), .B2(new_n790), .C1(new_n803), .C2(new_n490), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n799), .A2(new_n1029), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n793), .A2(new_n1027), .B1(new_n784), .B2(new_n778), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT115), .Z(new_n1045));
  AOI22_X1  g0845(.A1(G322), .A2(new_n812), .B1(new_n796), .B2(G311), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT48), .Z(new_n1048));
  AOI211_X1 g0848(.A(new_n1043), .B(new_n1048), .C1(G294), .C2(new_n805), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1042), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n289), .A2(new_n796), .B1(new_n791), .B2(G150), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n202), .B2(new_n793), .C1(new_n808), .C2(new_n780), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G77), .A2(new_n805), .B1(new_n785), .B2(G68), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(new_n264), .C1(new_n480), .C2(new_n803), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n799), .A2(new_n429), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n764), .B1(new_n1053), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n715), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1061), .A2(new_n767), .B1(new_n438), .B2(new_n712), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n236), .A2(new_n303), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT50), .B1(new_n291), .B2(G50), .ZN(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n715), .A3(new_n1065), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n291), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n771), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1062), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT114), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n766), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n758), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1060), .B(new_n1074), .C1(new_n702), .C2(new_n1037), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1004), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n713), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n752), .A2(new_n1040), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1041), .B(new_n1075), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  AND3_X1   g0879(.A1(new_n989), .A2(new_n995), .A3(new_n703), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n703), .B1(new_n989), .B2(new_n995), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1076), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n1005), .A3(new_n713), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT118), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n998), .A2(new_n756), .A3(new_n999), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n244), .A2(new_n1009), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n765), .B1(new_n480), .B2(new_n218), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n757), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G150), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n793), .A2(new_n808), .B1(new_n780), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G68), .A2(new_n805), .B1(new_n785), .B2(new_n289), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G50), .A2(new_n796), .B1(new_n791), .B2(G143), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n800), .A2(G77), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n270), .B1(new_n788), .B2(G87), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1092), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n264), .B(new_n804), .C1(new_n489), .C2(new_n800), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n785), .A2(G294), .B1(new_n791), .B2(G322), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n805), .A2(G283), .B1(new_n796), .B2(G303), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n793), .A2(new_n854), .B1(new_n780), .B2(new_n1027), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT52), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1099), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1089), .B1(new_n1107), .B2(new_n764), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT117), .Z(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n959), .B2(new_n1037), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1086), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1085), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G390));
  NAND4_X1  g0913(.A1(new_n944), .A2(G330), .A3(new_n929), .A4(new_n829), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n834), .A2(KEYINPUT104), .A3(new_n923), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT104), .B1(new_n834), .B2(new_n923), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n929), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n911), .B1(new_n1118), .B2(new_n913), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n929), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n920), .B1(new_n727), .B2(new_n829), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n908), .A2(new_n899), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n1123), .A3(new_n913), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1115), .B1(new_n1119), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n914), .B1(new_n925), .B2(new_n929), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1114), .B(new_n1124), .C1(new_n1127), .C2(new_n911), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1126), .A2(new_n1128), .A3(new_n756), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n757), .B1(new_n842), .B2(new_n289), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n803), .A2(new_n222), .B1(new_n1029), .B2(new_n780), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n264), .B(new_n1131), .C1(G87), .C2(new_n805), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G107), .A2(new_n796), .B1(new_n791), .B2(G294), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G116), .A2(new_n794), .B1(new_n785), .B2(G97), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1132), .A2(new_n1096), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n777), .A2(new_n1090), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT53), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n800), .A2(G159), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n791), .A2(G125), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n270), .B1(new_n788), .B2(G50), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT54), .B(G143), .Z(new_n1142));
  AOI22_X1  g0942(.A1(new_n785), .A2(new_n1142), .B1(new_n796), .B2(G137), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT120), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n793), .A2(new_n845), .B1(new_n780), .B2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT121), .Z(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1135), .B1(new_n1141), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1130), .B1(new_n1149), .B2(new_n764), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n911), .B2(new_n760), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT122), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G330), .B(new_n829), .C1(new_n747), .C2(new_n749), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1120), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1114), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1114), .A3(new_n1121), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n933), .A2(new_n640), .A3(new_n949), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT119), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n933), .A2(new_n949), .A3(KEYINPUT119), .A4(new_n640), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1158), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1126), .A2(new_n1163), .A3(new_n1128), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n713), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1129), .B(new_n1152), .C1(new_n1165), .C2(new_n1166), .ZN(G378));
  NAND2_X1  g0967(.A1(new_n639), .A2(new_n427), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n686), .A2(new_n414), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n948), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1172), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n947), .A2(G330), .A3(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1173), .A2(new_n930), .A3(new_n915), .A4(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n947), .A2(G330), .A3(new_n1174), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1174), .B1(new_n947), .B2(G330), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n931), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1172), .A2(new_n759), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n757), .B1(new_n842), .B2(G50), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT123), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n793), .A2(new_n1145), .B1(new_n795), .B2(new_n845), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n812), .A2(G125), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1142), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1185), .B1(new_n1013), .B2(new_n784), .C1(new_n777), .C2(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(G150), .C2(new_n800), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT59), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n788), .A2(G159), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n812), .A2(G116), .B1(new_n791), .B2(G283), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n480), .B2(new_n795), .C1(new_n438), .C2(new_n793), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n302), .B(new_n270), .C1(new_n777), .C2(new_n203), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n803), .A2(new_n221), .B1(new_n429), .B2(new_n784), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n1196), .A2(new_n1018), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G50), .B1(new_n266), .B2(new_n302), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n264), .B2(G41), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1194), .A2(new_n1200), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1183), .B1(new_n1204), .B2(new_n764), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1180), .A2(new_n756), .B1(new_n1181), .B2(new_n1205), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1162), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1164), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(KEYINPUT57), .A3(new_n1180), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n713), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1210), .B2(new_n1180), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1206), .B1(new_n1212), .B2(new_n1213), .ZN(G375));
  INV_X1    g1014(.A(new_n1163), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n984), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1120), .A2(new_n759), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n757), .B1(new_n842), .B2(G68), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n785), .A2(G150), .B1(new_n791), .B2(G128), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n808), .B2(new_n777), .C1(new_n795), .C2(new_n1186), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n794), .A2(G137), .B1(new_n812), .B2(G132), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n270), .B1(new_n788), .B2(G58), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n202), .C2(new_n799), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n489), .A2(new_n796), .B1(new_n791), .B2(G303), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n480), .B2(new_n777), .C1(new_n1029), .C2(new_n793), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n812), .A2(G294), .B1(new_n785), .B2(G107), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1058), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n270), .A3(new_n1012), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1222), .A2(new_n1225), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1220), .B1(new_n1231), .B2(new_n764), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1158), .A2(new_n756), .B1(new_n1219), .B2(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1218), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(G381));
  NAND2_X1  g1035(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT124), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n1206), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(G378), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1007), .A2(new_n1241), .A3(new_n1038), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1240), .A2(new_n1112), .A3(new_n1242), .A4(new_n1234), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT125), .B1(new_n1239), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT125), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1246), .B(new_n1243), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1245), .A2(new_n1247), .ZN(G407));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n704), .A2(G213), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(G378), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1249), .B1(new_n1239), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT126), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT126), .B(new_n1252), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(G409));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1206), .C1(new_n1212), .C2(new_n1213), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1210), .A2(new_n984), .A3(new_n1180), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1206), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1240), .A2(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1259), .A2(new_n1262), .B1(G213), .B2(new_n704), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1217), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1216), .B(KEYINPUT60), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n1215), .A3(new_n713), .A4(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G384), .B1(new_n1267), .B2(new_n1233), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(G384), .A3(new_n1233), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n704), .A2(G213), .A3(G2897), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1269), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1258), .B1(new_n1263), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1112), .A2(G387), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT127), .B1(new_n1112), .B2(G387), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1112), .A2(G387), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G393), .B(new_n821), .ZN(new_n1282));
  AND4_X1   g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .A4(new_n1282), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1279), .A2(new_n1281), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1250), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1286), .B1(new_n1288), .B2(new_n1271), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1271), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1278), .A2(new_n1285), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1263), .A2(new_n1293), .A3(new_n1290), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1293), .B1(new_n1263), .B2(new_n1290), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1294), .A2(new_n1277), .A3(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1296), .B2(new_n1285), .ZN(G405));
  NAND2_X1  g1097(.A1(G375), .A2(new_n1240), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1298), .A2(new_n1271), .A3(new_n1259), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1271), .B1(new_n1298), .B2(new_n1259), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1285), .ZN(G402));
endmodule


