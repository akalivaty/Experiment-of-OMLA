//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G2105), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(KEYINPUT64), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n469), .B2(new_n470), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND3_X1   g057(.A1(KEYINPUT64), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT3), .B1(KEYINPUT64), .B2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n475), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n468), .A2(new_n464), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(KEYINPUT4), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n475), .A2(G138), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n485), .A2(KEYINPUT4), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n475), .A2(G114), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT65), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n495), .A2(new_n494), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n476), .B2(G126), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n471), .B2(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n459), .A2(new_n460), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n498), .B(new_n500), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n497), .A2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n507), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT66), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n513), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  AND2_X1   g095(.A1(new_n507), .A2(new_n508), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT67), .B(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n511), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n528));
  AND4_X1   g103(.A1(new_n523), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(G168));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n509), .A2(new_n530), .B1(new_n511), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n507), .A2(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n514), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n536));
  OR3_X1    g111(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n532), .B2(new_n535), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(G171));
  XOR2_X1   g114(.A(KEYINPUT69), .B(G81), .Z(new_n540));
  NAND2_X1  g115(.A1(new_n521), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT5), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n541), .B(new_n550), .C1(new_n551), .C2(new_n511), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT70), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G188));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n514), .B1(new_n509), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n565), .A2(new_n567), .A3(G53), .A4(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n508), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n561), .B1(new_n564), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n544), .A2(new_n546), .A3(G65), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n521), .A2(G91), .B1(new_n576), .B2(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n569), .A2(new_n571), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(KEYINPUT71), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n573), .A2(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  NAND4_X1  g156(.A1(new_n525), .A2(new_n523), .A3(new_n527), .A4(new_n528), .ZN(G286));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n514), .B1(new_n547), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n524), .B2(G49), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT72), .B1(new_n509), .B2(new_n586), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(new_n521), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT74), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n521), .A2(new_n592), .A3(G86), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT73), .B1(new_n547), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n507), .A2(new_n598), .A3(G61), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(G47), .A2(new_n524), .B1(new_n521), .B2(G85), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n514), .B2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n547), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(G54), .A2(new_n524), .B1(new_n609), .B2(G651), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT10), .B1(new_n509), .B2(new_n611), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n509), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT75), .Z(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  NOR2_X1   g197(.A1(new_n615), .A2(G559), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(G860), .B2(new_n616), .ZN(G148));
  OAI21_X1  g199(.A(G868), .B1(new_n615), .B2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g202(.A1(new_n475), .A2(G111), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT77), .Z(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n476), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n471), .A2(G135), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT76), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n634), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT15), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2435), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(G14), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  NOR3_X1   g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT78), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n657), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n658), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n655), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n656), .C2(new_n658), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n672), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n682), .C1(new_n680), .C2(new_n679), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT80), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT32), .B(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1971), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n694), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT34), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G24), .ZN(new_n706));
  XOR2_X1   g281(.A(G290), .B(KEYINPUT82), .Z(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(G1986), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n476), .A2(G119), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n471), .A2(G131), .ZN(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT81), .B(G29), .ZN(new_n715));
  MUX2_X1   g290(.A(G25), .B(new_n714), .S(new_n715), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT35), .B(G1991), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  NAND3_X1  g293(.A1(new_n705), .A2(new_n709), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT36), .Z(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G33), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n471), .A2(G139), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT85), .ZN(new_n727));
  INV_X1    g302(.A(G127), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  OAI21_X1  g305(.A(G2105), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n721), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G2072), .Z(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT87), .B(KEYINPUT24), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G34), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n473), .A2(new_n737), .B1(new_n715), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n476), .A2(G129), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT26), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n471), .A2(G141), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n465), .A2(G105), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n743), .A2(new_n745), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT88), .Z(new_n749));
  MUX2_X1   g324(.A(G32), .B(new_n749), .S(G29), .Z(new_n750));
  XOR2_X1   g325(.A(KEYINPUT27), .B(G1996), .Z(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n736), .A2(new_n742), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT89), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n736), .A2(new_n755), .A3(new_n742), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n715), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n758), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G2090), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT93), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n633), .A2(new_n715), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT90), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT31), .B(G11), .ZN(new_n767));
  AND2_X1   g342(.A1(KEYINPUT30), .A2(G28), .ZN(new_n768));
  NOR2_X1   g343(.A1(KEYINPUT30), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n737), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT91), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n695), .A2(KEYINPUT23), .A3(G20), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT23), .ZN(new_n774));
  INV_X1    g349(.A(G20), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G16), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n776), .C1(new_n620), .C2(new_n695), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(G168), .A2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G16), .B2(G21), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n553), .A2(new_n695), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n695), .B2(G19), .ZN(new_n786));
  INV_X1    g361(.A(G1341), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n787), .B2(new_n786), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n740), .A2(new_n741), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n762), .B2(G2090), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n695), .A2(G5), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G171), .B2(new_n695), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n791), .B1(G1961), .B2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(G1961), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n715), .A2(G27), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G164), .B2(new_n715), .ZN(new_n797));
  INV_X1    g372(.A(G2078), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n789), .A2(new_n794), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n758), .A2(G26), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT84), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT28), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n804));
  INV_X1    g379(.A(G116), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(G2105), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT83), .ZN(new_n807));
  AOI22_X1  g382(.A1(G128), .A2(new_n476), .B1(new_n471), .B2(G140), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n803), .B1(G29), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G2067), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n812), .B(new_n813), .C1(new_n783), .C2(new_n782), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n750), .A2(new_n751), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n780), .A2(new_n800), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G4), .A2(G16), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n616), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(G1348), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n757), .A2(new_n764), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(KEYINPUT94), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(KEYINPUT94), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n720), .B1(new_n823), .B2(new_n824), .ZN(G311));
  INV_X1    g400(.A(new_n720), .ZN(new_n826));
  INV_X1    g401(.A(new_n824), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n822), .ZN(G150));
  XNOR2_X1  g403(.A(KEYINPUT95), .B(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n509), .A2(new_n829), .B1(new_n511), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n514), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(G860), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n616), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n831), .A2(new_n833), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n552), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT39), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n838), .B(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n836), .B1(new_n842), .B2(G860), .ZN(G145));
  XNOR2_X1  g418(.A(new_n481), .B(KEYINPUT96), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G160), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n714), .B(new_n636), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n471), .A2(G142), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n476), .A2(G130), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n475), .A2(G118), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n748), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n500), .B1(new_n502), .B2(new_n504), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n809), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n488), .A2(new_n490), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n807), .A2(new_n500), .A3(new_n860), .A4(new_n808), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT97), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(KEYINPUT97), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n855), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n748), .A3(new_n863), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n868), .A3(new_n732), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n749), .A2(new_n862), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n749), .A2(new_n862), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n734), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n870), .B1(new_n869), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n854), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n633), .ZN(new_n878));
  INV_X1    g453(.A(new_n854), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n878), .B1(new_n877), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n846), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n877), .A2(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n633), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n845), .A3(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g465(.A(new_n614), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(G299), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT100), .B1(new_n573), .B2(new_n579), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n893), .A2(new_n894), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n620), .A2(KEYINPUT100), .A3(new_n891), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT41), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT101), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n899), .A2(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n896), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n623), .B(new_n840), .ZN(new_n908));
  MUX2_X1   g483(.A(new_n906), .B(new_n907), .S(new_n908), .Z(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(KEYINPUT42), .ZN(new_n910));
  XNOR2_X1  g485(.A(G305), .B(G288), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G290), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(KEYINPUT42), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(G868), .B2(new_n839), .ZN(G295));
  OAI21_X1  g493(.A(new_n917), .B1(G868), .B2(new_n839), .ZN(G331));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g496(.A1(G171), .A2(G286), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n537), .A2(G168), .A3(new_n538), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT102), .B1(new_n924), .B2(new_n840), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n834), .B(new_n552), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n922), .A3(new_n927), .A4(new_n923), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n924), .B2(new_n840), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n537), .A2(G168), .A3(new_n538), .ZN(new_n931));
  AOI21_X1  g506(.A(G168), .B1(new_n537), .B2(new_n538), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n840), .B(new_n929), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n925), .B(new_n928), .C1(new_n930), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n902), .A2(new_n935), .A3(new_n905), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n913), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n924), .B(new_n926), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n903), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n902), .A2(new_n935), .A3(KEYINPUT104), .A4(new_n905), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n938), .A2(new_n939), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(new_n885), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n913), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n921), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n935), .A2(new_n907), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n940), .B1(new_n898), .B2(new_n901), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n913), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n885), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n920), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n946), .A2(new_n921), .A3(new_n885), .A4(new_n943), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT44), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(G397));
  NAND3_X1  g534(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n860), .B2(new_n500), .ZN(new_n961));
  INV_X1    g536(.A(G125), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n486), .B2(new_n487), .ZN(new_n963));
  INV_X1    g538(.A(new_n462), .ZN(new_n964));
  OAI21_X1  g539(.A(G2105), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n465), .A2(G101), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n965), .A2(new_n472), .A3(G40), .A4(new_n966), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(G1996), .A3(new_n748), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT106), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n749), .A2(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n809), .A2(G2067), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n960), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n968), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n714), .A2(new_n717), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(KEYINPUT126), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n960), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n968), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n968), .B1(new_n973), .B2(new_n748), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n968), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  INV_X1    g563(.A(new_n968), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n714), .B(new_n717), .ZN(new_n990));
  XOR2_X1   g565(.A(new_n990), .B(KEYINPUT107), .Z(new_n991));
  OAI21_X1  g566(.A(new_n975), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n989), .A2(G1986), .A3(G290), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT48), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n981), .B(new_n988), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  XNOR2_X1  g571(.A(G290), .B(G1986), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n992), .B1(new_n968), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT59), .ZN(new_n999));
  INV_X1    g574(.A(new_n967), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n961), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT58), .B(G1341), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(KEYINPUT119), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT45), .B(new_n1009), .C1(new_n491), .C2(new_n496), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n1000), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n497), .A2(new_n505), .A3(new_n1009), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n983), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1014), .B2(new_n983), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1008), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT120), .B1(new_n1018), .B2(new_n553), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1020), .B(new_n1000), .C1(new_n961), .C2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n466), .A2(new_n1021), .A3(G40), .A4(new_n472), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1009), .B1(new_n491), .B2(new_n496), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(KEYINPUT111), .C1(new_n1024), .C2(new_n967), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n497), .A2(new_n505), .A3(new_n1021), .A4(new_n1009), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n778), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(G2072), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1014), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n578), .A2(KEYINPUT114), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n569), .A2(new_n571), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n577), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT113), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n564), .A2(new_n572), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1038), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1044), .B(new_n1038), .C1(new_n1041), .C2(new_n1037), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1032), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1027), .A2(new_n778), .B1(new_n1014), .B2(new_n1030), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n569), .A2(new_n571), .A3(new_n1034), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1034), .B1(new_n569), .B2(new_n571), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT113), .B1(new_n1050), .B2(new_n577), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT57), .B1(new_n1051), .B2(new_n1039), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1044), .B1(new_n1052), .B2(new_n1038), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1045), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1047), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1046), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n999), .A2(new_n1019), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n1032), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1062), .A2(KEYINPUT117), .A3(new_n1047), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT61), .B(new_n1055), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1013), .A2(new_n1012), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1011), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT118), .B1(new_n1068), .B2(G1996), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1014), .A2(new_n1015), .A3(new_n983), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1007), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1065), .B1(new_n1071), .B2(new_n552), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1018), .A2(KEYINPUT120), .A3(new_n553), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(KEYINPUT59), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n961), .A2(new_n1021), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1000), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1001), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1077), .A2(new_n819), .B1(new_n811), .B2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1079), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n614), .B1(new_n1079), .B2(KEYINPUT60), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1080), .A2(new_n1081), .B1(KEYINPUT60), .B2(new_n1079), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1058), .A2(new_n1064), .A3(new_n1074), .A4(new_n1082), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1061), .A2(new_n1063), .B1(new_n614), .B2(new_n1079), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1055), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT108), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1068), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n798), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  INV_X1    g666(.A(G1961), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1091), .B1(new_n1092), .B2(new_n1077), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT45), .B1(new_n856), .B2(new_n1009), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(new_n967), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n967), .B1(new_n1024), .B2(new_n1012), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT112), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n497), .A2(new_n505), .A3(KEYINPUT45), .A4(new_n1009), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OR3_X1    g675(.A1(new_n1100), .A2(new_n1091), .A3(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1093), .A2(G301), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1097), .A2(KEYINPUT53), .A3(new_n798), .A4(new_n1010), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1102), .B(KEYINPUT54), .C1(new_n1106), .C2(G301), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT49), .ZN(new_n1108));
  INV_X1    g683(.A(G1981), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n594), .A2(new_n601), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n601), .B2(new_n590), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G8), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1078), .A2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n601), .A2(new_n590), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1110), .B(KEYINPUT49), .C1(new_n1116), .C2(new_n1109), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1113), .A2(KEYINPUT110), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1976), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1115), .B1(new_n1123), .B2(G288), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT52), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n700), .A2(G1976), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n1124), .A2(KEYINPUT52), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1122), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1971), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1066), .A2(KEYINPUT108), .A3(new_n1067), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT108), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1027), .A2(G2090), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1114), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(G303), .A2(G8), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT55), .Z(new_n1136));
  NOR2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1128), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT109), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1077), .A2(G2090), .ZN(new_n1141));
  OAI211_X1 g716(.A(KEYINPUT109), .B(new_n1129), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(G8), .A3(new_n1136), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1107), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(G286), .A2(G8), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT121), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT51), .B1(new_n1147), .B2(KEYINPUT122), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1075), .A2(new_n1000), .A3(new_n1076), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n741), .A2(new_n1150), .B1(new_n1100), .B2(new_n783), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1147), .B(new_n1149), .C1(new_n1151), .C2(new_n1114), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1099), .B1(new_n1097), .B2(KEYINPUT112), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1095), .A2(new_n1094), .A3(new_n967), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n783), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1075), .A2(new_n741), .A3(new_n1000), .A4(new_n1076), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1114), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1147), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1148), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1158), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1152), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1093), .A2(new_n1163), .A3(G301), .A4(new_n1105), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1093), .A2(G301), .A3(new_n1105), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1103), .A2(new_n1104), .A3(new_n1101), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1167), .B(KEYINPUT123), .C1(new_n1168), .C2(G301), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1162), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1086), .A2(new_n1145), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1143), .A2(G8), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1136), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1128), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1114), .B(G286), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT63), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1179), .B(new_n1176), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1144), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1122), .A2(new_n1123), .A3(new_n700), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1110), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1181), .A2(new_n1175), .B1(new_n1183), .B2(new_n1115), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT124), .B1(new_n1162), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1152), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(new_n1188), .A3(KEYINPUT62), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1168), .A2(G301), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1152), .A2(new_n1159), .A3(new_n1185), .A4(new_n1161), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1138), .A2(new_n1191), .A3(new_n1144), .A4(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1178), .B(new_n1184), .C1(new_n1190), .C2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g769(.A(KEYINPUT125), .B(new_n998), .C1(new_n1171), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1086), .A2(new_n1145), .A3(new_n1170), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1181), .A2(new_n1175), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1183), .A2(new_n1115), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1128), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1179), .B1(new_n1201), .B2(new_n1176), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1204), .A2(new_n1205), .A3(new_n1186), .A4(new_n1189), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1197), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(KEYINPUT125), .B1(new_n1207), .B2(new_n998), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n996), .B1(new_n1196), .B2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g784(.A(G319), .ZN(new_n1211));
  AOI211_X1 g785(.A(new_n1211), .B(G227), .C1(new_n653), .C2(G14), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1212), .A2(new_n889), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n947), .A2(new_n952), .ZN(new_n1214));
  NOR3_X1   g788(.A1(new_n1213), .A2(new_n1214), .A3(G229), .ZN(G308));
  NOR2_X1   g789(.A1(new_n1214), .A2(G229), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n1216), .A2(new_n889), .A3(new_n1212), .ZN(G225));
endmodule


