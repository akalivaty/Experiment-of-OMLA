

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595;

  AND2_X1 U326 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U327 ( .A(n360), .B(n329), .Z(n295) );
  XOR2_X1 U328 ( .A(KEYINPUT94), .B(n423), .Z(n296) );
  XNOR2_X1 U329 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n500) );
  XNOR2_X1 U330 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U331 ( .A(KEYINPUT0), .B(G127GAT), .Z(n409) );
  XNOR2_X1 U332 ( .A(n514), .B(KEYINPUT64), .ZN(n515) );
  XNOR2_X1 U333 ( .A(n365), .B(n294), .ZN(n366) );
  XNOR2_X1 U334 ( .A(n357), .B(n295), .ZN(n311) );
  XNOR2_X1 U335 ( .A(n516), .B(n515), .ZN(n546) );
  XNOR2_X1 U336 ( .A(n367), .B(n366), .ZN(n371) );
  XNOR2_X1 U337 ( .A(n312), .B(n311), .ZN(n477) );
  XNOR2_X1 U338 ( .A(n557), .B(n556), .ZN(n570) );
  XOR2_X1 U339 ( .A(n377), .B(n376), .Z(n494) );
  XOR2_X1 U340 ( .A(KEYINPUT98), .B(n448), .Z(n473) );
  XNOR2_X1 U341 ( .A(n454), .B(G50GAT), .ZN(n455) );
  XNOR2_X1 U342 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U343 ( .A(n456), .B(n455), .ZN(G1331GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT38), .B(KEYINPUT97), .Z(n447) );
  XNOR2_X1 U345 ( .A(G106GAT), .B(G78GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n297), .B(G148GAT), .ZN(n385) );
  INV_X1 U347 ( .A(n385), .ZN(n299) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G85GAT), .Z(n428) );
  INV_X1 U349 ( .A(n428), .ZN(n298) );
  NAND2_X1 U350 ( .A1(n299), .A2(n298), .ZN(n301) );
  NAND2_X1 U351 ( .A1(n428), .A2(n385), .ZN(n300) );
  NAND2_X1 U352 ( .A1(n301), .A2(n300), .ZN(n303) );
  AND2_X1 U353 ( .A1(G230GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U355 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n305) );
  XNOR2_X1 U356 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n304) );
  XOR2_X1 U357 ( .A(n305), .B(n304), .Z(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n312) );
  XOR2_X1 U359 ( .A(KEYINPUT72), .B(G64GAT), .Z(n309) );
  XNOR2_X1 U360 ( .A(G176GAT), .B(G92GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U362 ( .A(G204GAT), .B(n310), .Z(n357) );
  XOR2_X1 U363 ( .A(G120GAT), .B(G71GAT), .Z(n360) );
  XOR2_X1 U364 ( .A(G57GAT), .B(KEYINPUT13), .Z(n329) );
  XOR2_X1 U365 ( .A(G43GAT), .B(G29GAT), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U368 ( .A(n315), .B(KEYINPUT69), .Z(n317) );
  XNOR2_X1 U369 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n443) );
  XOR2_X1 U371 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n319) );
  XNOR2_X1 U372 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U374 ( .A(G141GAT), .B(G22GAT), .Z(n390) );
  XNOR2_X1 U375 ( .A(n320), .B(n390), .ZN(n324) );
  XOR2_X1 U376 ( .A(G113GAT), .B(G1GAT), .Z(n413) );
  XOR2_X1 U377 ( .A(n413), .B(KEYINPUT29), .Z(n322) );
  NAND2_X1 U378 ( .A1(G229GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U381 ( .A(G169GAT), .B(G8GAT), .Z(n347) );
  XOR2_X1 U382 ( .A(n325), .B(n347), .Z(n327) );
  XNOR2_X1 U383 ( .A(G15GAT), .B(G197GAT), .ZN(n326) );
  XOR2_X1 U384 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U385 ( .A(n443), .B(n328), .ZN(n531) );
  XOR2_X1 U386 ( .A(KEYINPUT71), .B(n531), .Z(n558) );
  INV_X1 U387 ( .A(n558), .ZN(n519) );
  NOR2_X1 U388 ( .A1(n477), .A2(n519), .ZN(n460) );
  XOR2_X1 U389 ( .A(KEYINPUT76), .B(n329), .Z(n331) );
  NAND2_X1 U390 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U392 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n333) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G1GAT), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U395 ( .A(n335), .B(n334), .Z(n337) );
  XNOR2_X1 U396 ( .A(G15GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n345) );
  XOR2_X1 U398 ( .A(G155GAT), .B(G78GAT), .Z(n339) );
  XNOR2_X1 U399 ( .A(G71GAT), .B(G127GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U401 ( .A(G64GAT), .B(KEYINPUT12), .Z(n341) );
  XNOR2_X1 U402 ( .A(G22GAT), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U404 ( .A(n343), .B(n342), .Z(n344) );
  XOR2_X1 U405 ( .A(n345), .B(n344), .Z(n589) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n346), .B(G211GAT), .ZN(n388) );
  XOR2_X1 U408 ( .A(n388), .B(n347), .Z(n349) );
  NAND2_X1 U409 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U411 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n351) );
  XNOR2_X1 U412 ( .A(G36GAT), .B(G218GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U414 ( .A(n353), .B(n352), .Z(n359) );
  XOR2_X1 U415 ( .A(KEYINPUT18), .B(G190GAT), .Z(n355) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U418 ( .A(KEYINPUT19), .B(n356), .Z(n375) );
  XNOR2_X1 U419 ( .A(n375), .B(n357), .ZN(n358) );
  XOR2_X1 U420 ( .A(n359), .B(n358), .Z(n474) );
  XOR2_X1 U421 ( .A(G99GAT), .B(n409), .Z(n362) );
  XNOR2_X1 U422 ( .A(G43GAT), .B(n360), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U424 ( .A(KEYINPUT77), .B(KEYINPUT82), .Z(n364) );
  XNOR2_X1 U425 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U427 ( .A(KEYINPUT80), .B(G176GAT), .Z(n369) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G134GAT), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U431 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n373) );
  XNOR2_X1 U432 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n372) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  INV_X1 U435 ( .A(n494), .ZN(n554) );
  NAND2_X1 U436 ( .A1(n474), .A2(n554), .ZN(n395) );
  XOR2_X1 U437 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n379) );
  XNOR2_X1 U438 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n394) );
  XOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n381) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U443 ( .A(n382), .B(G204GAT), .Z(n387) );
  XOR2_X1 U444 ( .A(G155GAT), .B(KEYINPUT2), .Z(n384) );
  XNOR2_X1 U445 ( .A(KEYINPUT3), .B(KEYINPUT83), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n417) );
  XNOR2_X1 U447 ( .A(n385), .B(n417), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U449 ( .A(n389), .B(n388), .Z(n392) );
  XOR2_X1 U450 ( .A(G218GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U451 ( .A(n390), .B(n439), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n549) );
  NAND2_X1 U454 ( .A1(n395), .A2(n549), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n396), .B(KEYINPUT25), .ZN(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT93), .B(n397), .ZN(n400) );
  NOR2_X1 U457 ( .A1(n554), .A2(n549), .ZN(n399) );
  XNOR2_X1 U458 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n579) );
  XNOR2_X1 U460 ( .A(n474), .B(KEYINPUT27), .ZN(n424) );
  NAND2_X1 U461 ( .A1(n579), .A2(n424), .ZN(n532) );
  NAND2_X1 U462 ( .A1(n400), .A2(n532), .ZN(n422) );
  XOR2_X1 U463 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n402) );
  XNOR2_X1 U464 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n421) );
  XOR2_X1 U466 ( .A(G85GAT), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(G120GAT), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U469 ( .A(KEYINPUT5), .B(G57GAT), .Z(n406) );
  XNOR2_X1 U470 ( .A(G141GAT), .B(G148GAT), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U472 ( .A(n408), .B(n407), .Z(n415) );
  XOR2_X1 U473 ( .A(G134GAT), .B(KEYINPUT74), .Z(n429) );
  XOR2_X1 U474 ( .A(n429), .B(n409), .Z(n411) );
  NAND2_X1 U475 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U479 ( .A(n416), .B(KEYINPUT86), .Z(n419) );
  XNOR2_X1 U480 ( .A(n417), .B(KEYINPUT6), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U482 ( .A(n421), .B(n420), .Z(n551) );
  NAND2_X1 U483 ( .A1(n422), .A2(n551), .ZN(n423) );
  XNOR2_X1 U484 ( .A(KEYINPUT28), .B(n549), .ZN(n497) );
  AND2_X1 U485 ( .A1(n424), .A2(n497), .ZN(n425) );
  INV_X1 U486 ( .A(n551), .ZN(n578) );
  NAND2_X1 U487 ( .A1(n425), .A2(n578), .ZN(n517) );
  NOR2_X1 U488 ( .A1(n554), .A2(n517), .ZN(n426) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(n426), .Z(n427) );
  NOR2_X1 U490 ( .A1(n296), .A2(n427), .ZN(n459) );
  XOR2_X1 U491 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U492 ( .A1(G232GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U494 ( .A(G92GAT), .B(KEYINPUT11), .Z(n433) );
  XNOR2_X1 U495 ( .A(G190GAT), .B(G106GAT), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U497 ( .A(n435), .B(n434), .Z(n441) );
  XOR2_X1 U498 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n437) );
  XNOR2_X1 U499 ( .A(KEYINPUT65), .B(KEYINPUT75), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n569) );
  XOR2_X1 U504 ( .A(n569), .B(KEYINPUT36), .Z(n593) );
  NOR2_X1 U505 ( .A1(n459), .A2(n593), .ZN(n444) );
  NAND2_X1 U506 ( .A1(n589), .A2(n444), .ZN(n445) );
  XNOR2_X1 U507 ( .A(KEYINPUT37), .B(n445), .ZN(n490) );
  NAND2_X1 U508 ( .A1(n460), .A2(n490), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  NAND2_X1 U510 ( .A1(n473), .A2(n554), .ZN(n452) );
  XOR2_X1 U511 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n450) );
  XNOR2_X1 U512 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(G1330GAT) );
  INV_X1 U514 ( .A(n497), .ZN(n453) );
  NAND2_X1 U515 ( .A1(n473), .A2(n453), .ZN(n456) );
  XOR2_X1 U516 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n454) );
  NOR2_X1 U517 ( .A1(n589), .A2(n569), .ZN(n457) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(n457), .Z(n458) );
  NOR2_X1 U519 ( .A1(n459), .A2(n458), .ZN(n478) );
  NAND2_X1 U520 ( .A1(n460), .A2(n478), .ZN(n467) );
  NOR2_X1 U521 ( .A1(n551), .A2(n467), .ZN(n461) );
  XOR2_X1 U522 ( .A(G1GAT), .B(n461), .Z(n462) );
  XNOR2_X1 U523 ( .A(KEYINPUT34), .B(n462), .ZN(G1324GAT) );
  INV_X1 U524 ( .A(n474), .ZN(n545) );
  NOR2_X1 U525 ( .A1(n545), .A2(n467), .ZN(n463) );
  XOR2_X1 U526 ( .A(G8GAT), .B(n463), .Z(G1325GAT) );
  NOR2_X1 U527 ( .A1(n494), .A2(n467), .ZN(n465) );
  XNOR2_X1 U528 ( .A(KEYINPUT95), .B(KEYINPUT35), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U530 ( .A(G15GAT), .B(n466), .Z(G1326GAT) );
  NOR2_X1 U531 ( .A1(n497), .A2(n467), .ZN(n468) );
  XOR2_X1 U532 ( .A(KEYINPUT96), .B(n468), .Z(n469) );
  XNOR2_X1 U533 ( .A(G22GAT), .B(n469), .ZN(G1327GAT) );
  XNOR2_X1 U534 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n578), .A2(n473), .ZN(n470) );
  XNOR2_X1 U536 ( .A(n470), .B(KEYINPUT39), .ZN(n471) );
  XNOR2_X1 U537 ( .A(n472), .B(n471), .ZN(G1328GAT) );
  NAND2_X1 U538 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n475), .B(KEYINPUT100), .ZN(n476) );
  XNOR2_X1 U540 ( .A(G36GAT), .B(n476), .ZN(G1329GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT41), .B(n477), .Z(n560) );
  INV_X1 U542 ( .A(n560), .ZN(n537) );
  NOR2_X1 U543 ( .A1(n531), .A2(n537), .ZN(n489) );
  NAND2_X1 U544 ( .A1(n478), .A2(n489), .ZN(n479) );
  XOR2_X1 U545 ( .A(KEYINPUT105), .B(n479), .Z(n486) );
  NOR2_X1 U546 ( .A1(n551), .A2(n486), .ZN(n481) );
  XNOR2_X1 U547 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n480) );
  XNOR2_X1 U548 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U549 ( .A(G57GAT), .B(n482), .Z(G1332GAT) );
  NOR2_X1 U550 ( .A1(n545), .A2(n486), .ZN(n483) );
  XOR2_X1 U551 ( .A(G64GAT), .B(n483), .Z(G1333GAT) );
  NOR2_X1 U552 ( .A1(n494), .A2(n486), .ZN(n485) );
  XNOR2_X1 U553 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n484) );
  XNOR2_X1 U554 ( .A(n485), .B(n484), .ZN(G1334GAT) );
  NOR2_X1 U555 ( .A1(n497), .A2(n486), .ZN(n488) );
  XNOR2_X1 U556 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n487) );
  XNOR2_X1 U557 ( .A(n488), .B(n487), .ZN(G1335GAT) );
  NAND2_X1 U558 ( .A1(n490), .A2(n489), .ZN(n496) );
  NOR2_X1 U559 ( .A1(n551), .A2(n496), .ZN(n491) );
  XOR2_X1 U560 ( .A(G85GAT), .B(n491), .Z(G1336GAT) );
  NOR2_X1 U561 ( .A1(n545), .A2(n496), .ZN(n492) );
  XOR2_X1 U562 ( .A(KEYINPUT108), .B(n492), .Z(n493) );
  XNOR2_X1 U563 ( .A(G92GAT), .B(n493), .ZN(G1337GAT) );
  NOR2_X1 U564 ( .A1(n494), .A2(n496), .ZN(n495) );
  XOR2_X1 U565 ( .A(G99GAT), .B(n495), .Z(G1338GAT) );
  NOR2_X1 U566 ( .A1(n497), .A2(n496), .ZN(n498) );
  XOR2_X1 U567 ( .A(KEYINPUT44), .B(n498), .Z(n499) );
  XNOR2_X1 U568 ( .A(G106GAT), .B(n499), .ZN(G1339GAT) );
  INV_X1 U569 ( .A(n589), .ZN(n566) );
  NAND2_X1 U570 ( .A1(n531), .A2(n560), .ZN(n501) );
  NOR2_X1 U571 ( .A1(n566), .A2(n502), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n503), .B(KEYINPUT110), .ZN(n504) );
  INV_X1 U573 ( .A(n569), .ZN(n543) );
  NAND2_X1 U574 ( .A1(n504), .A2(n543), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n505), .B(KEYINPUT111), .ZN(n506) );
  XNOR2_X1 U576 ( .A(KEYINPUT47), .B(n506), .ZN(n513) );
  XNOR2_X1 U577 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n508) );
  NOR2_X1 U578 ( .A1(n593), .A2(n589), .ZN(n507) );
  XOR2_X1 U579 ( .A(n508), .B(n507), .Z(n509) );
  NOR2_X1 U580 ( .A1(n477), .A2(n509), .ZN(n510) );
  XNOR2_X1 U581 ( .A(n510), .B(KEYINPUT112), .ZN(n511) );
  NAND2_X1 U582 ( .A1(n511), .A2(n519), .ZN(n512) );
  NAND2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n516) );
  INV_X1 U584 ( .A(KEYINPUT48), .ZN(n514) );
  NOR2_X1 U585 ( .A1(n546), .A2(n517), .ZN(n518) );
  NAND2_X1 U586 ( .A1(n554), .A2(n518), .ZN(n527) );
  NOR2_X1 U587 ( .A1(n519), .A2(n527), .ZN(n520) );
  XOR2_X1 U588 ( .A(G113GAT), .B(n520), .Z(G1340GAT) );
  NOR2_X1 U589 ( .A1(n537), .A2(n527), .ZN(n522) );
  XNOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U592 ( .A(G120GAT), .B(n523), .Z(G1341GAT) );
  NOR2_X1 U593 ( .A1(n589), .A2(n527), .ZN(n525) );
  XNOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U596 ( .A(G127GAT), .B(n526), .Z(G1342GAT) );
  NOR2_X1 U597 ( .A1(n543), .A2(n527), .ZN(n529) );
  XNOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n528) );
  XNOR2_X1 U599 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U600 ( .A(G134GAT), .B(n530), .Z(G1343GAT) );
  INV_X1 U601 ( .A(n531), .ZN(n581) );
  NOR2_X1 U602 ( .A1(n546), .A2(n532), .ZN(n533) );
  NAND2_X1 U603 ( .A1(n533), .A2(n578), .ZN(n542) );
  NOR2_X1 U604 ( .A1(n581), .A2(n542), .ZN(n534) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n534), .Z(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n536) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n535) );
  XNOR2_X1 U608 ( .A(n536), .B(n535), .ZN(n539) );
  NOR2_X1 U609 ( .A1(n537), .A2(n542), .ZN(n538) );
  XOR2_X1 U610 ( .A(n539), .B(n538), .Z(G1345GAT) );
  NOR2_X1 U611 ( .A1(n589), .A2(n542), .ZN(n541) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n540) );
  XNOR2_X1 U613 ( .A(n541), .B(n540), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U615 ( .A(G162GAT), .B(n544), .Z(G1347GAT) );
  NOR2_X1 U616 ( .A1(n546), .A2(n545), .ZN(n548) );
  INV_X1 U617 ( .A(KEYINPUT54), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n548), .B(n547), .ZN(n577) );
  INV_X1 U619 ( .A(n549), .ZN(n550) );
  NOR2_X1 U620 ( .A1(n577), .A2(n550), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n553), .B(KEYINPUT55), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U624 ( .A(KEYINPUT118), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n570), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n570), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n562) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n563), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT121), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n574) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT122), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT123), .B(n572), .Z(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1351GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n592) );
  NOR2_X1 U646 ( .A1(n581), .A2(n592), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1352GAT) );
  INV_X1 U648 ( .A(n477), .ZN(n584) );
  NOR2_X1 U649 ( .A1(n592), .A2(n584), .ZN(n588) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U654 ( .A1(n589), .A2(n592), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1354GAT) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT62), .B(n594), .Z(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

