//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n209));
  AND4_X1   g0009(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G250), .B1(G257), .B2(G264), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g0021(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n218), .A2(KEYINPUT0), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n218), .A2(KEYINPUT0), .ZN(new_n230));
  AND3_X1   g0030(.A1(new_n214), .A2(new_n229), .A3(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(G1), .B(G13), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  AND2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G226), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G77), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G1698), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n265), .B(new_n267), .C1(new_n260), .C2(new_n261), .ZN(new_n268));
  INV_X1    g0068(.A(G222), .ZN(new_n269));
  OR2_X1    g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n263), .B1(new_n268), .B2(new_n269), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n221), .A2(new_n222), .B1(G33), .B2(G41), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n259), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT73), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(G169), .B2(new_n277), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT70), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G58), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n224), .A2(G33), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n283), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n211), .B2(new_n249), .ZN(new_n294));
  NAND4_X1  g0094(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n294), .A2(new_n221), .A3(new_n222), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n215), .A2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G50), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n252), .A2(G20), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT71), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n303), .A2(new_n296), .A3(new_n300), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n301), .B1(new_n304), .B2(G50), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI211_X1 g0107(.A(KEYINPUT72), .B(new_n301), .C1(new_n304), .C2(G50), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n297), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n281), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n262), .A2(G107), .ZN(new_n312));
  INV_X1    g0112(.A(G232), .ZN(new_n313));
  INV_X1    g0113(.A(G238), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n312), .B1(new_n268), .B2(new_n313), .C1(new_n273), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n276), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n257), .B1(new_n254), .B2(G244), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G190), .B2(new_n318), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n223), .A2(new_n294), .A3(new_n295), .A4(new_n299), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n303), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G77), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G20), .A2(G77), .ZN(new_n325));
  INV_X1    g0125(.A(new_n282), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT15), .B(G87), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(new_n284), .B2(new_n326), .C1(new_n291), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n296), .ZN(new_n329));
  INV_X1    g0129(.A(G77), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n300), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n324), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n321), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n318), .A2(G169), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n278), .B2(new_n318), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n332), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n311), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n268), .A2(new_n274), .ZN(new_n339));
  OAI211_X1 g0139(.A(G226), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G87), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n276), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n251), .A2(G232), .A3(new_n253), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n258), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n341), .B(new_n340), .C1(new_n268), .C2(new_n274), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n345), .B1(new_n350), .B2(new_n276), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n278), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n290), .A2(new_n299), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n323), .B2(new_n290), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n270), .A2(new_n224), .A3(new_n271), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT77), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n224), .A4(new_n271), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n262), .A2(KEYINPUT77), .A3(KEYINPUT7), .A4(new_n224), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(G68), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G68), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n287), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n201), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n282), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT16), .B1(new_n364), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT7), .B1(new_n262), .B2(new_n224), .ZN(new_n372));
  INV_X1    g0172(.A(new_n361), .ZN(new_n373));
  OAI21_X1  g0173(.A(G68), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n296), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n356), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n354), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT18), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT78), .B(G190), .ZN(new_n381));
  AND4_X1   g0181(.A1(KEYINPUT79), .A2(new_n343), .A3(new_n346), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n351), .A2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT79), .B1(new_n351), .B2(G200), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n380), .B1(new_n385), .B2(new_n377), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n383), .ZN(new_n387));
  INV_X1    g0187(.A(new_n382), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n289), .A2(new_n300), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n304), .B2(new_n289), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n364), .A2(new_n370), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n296), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n359), .A2(new_n361), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n369), .B1(new_n396), .B2(G68), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n391), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n389), .A2(new_n399), .A3(KEYINPUT17), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n354), .A2(new_n377), .A3(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n379), .A2(new_n386), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n365), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n330), .B2(new_n291), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n406), .A2(new_n296), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n407), .A2(KEYINPUT11), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n323), .A2(G68), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(KEYINPUT11), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n298), .A2(G20), .A3(new_n365), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT12), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  INV_X1    g0215(.A(G226), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n415), .B1(new_n268), .B2(new_n416), .C1(new_n273), .C2(new_n313), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n276), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n257), .B1(new_n254), .B2(G238), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n419), .B1(new_n418), .B2(new_n420), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n422), .A2(new_n423), .A3(G190), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n418), .A2(new_n420), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n426));
  AOI21_X1  g0226(.A(G200), .B1(new_n426), .B2(new_n421), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n414), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n414), .C1(new_n424), .C2(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(G169), .B1(new_n422), .B2(new_n423), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(new_n421), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(G169), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n434), .B(new_n437), .C1(new_n278), .C2(new_n435), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n413), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n338), .A2(new_n404), .A3(new_n432), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT9), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n309), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT74), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n277), .A2(new_n443), .A3(G190), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n277), .B2(G190), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n277), .A2(new_n319), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(KEYINPUT9), .B(new_n297), .C1(new_n307), .C2(new_n308), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n449), .A2(KEYINPUT10), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT10), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n451), .B1(new_n449), .B2(KEYINPUT10), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n440), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT80), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT6), .ZN(new_n459));
  AND2_X1   g0259(.A1(G97), .A2(G107), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G97), .A2(G107), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G107), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(KEYINPUT6), .A3(G97), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n224), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n326), .A2(new_n330), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n466), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n463), .A2(KEYINPUT6), .A3(G97), .ZN(new_n469));
  XNOR2_X1  g0269(.A(G97), .B(G107), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(new_n459), .ZN(new_n471));
  OAI211_X1 g0271(.A(KEYINPUT80), .B(new_n468), .C1(new_n471), .C2(new_n224), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n362), .A2(G107), .A3(new_n363), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n395), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n299), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n249), .A2(G1), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n296), .A2(new_n300), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n479), .B2(new_n476), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  OAI21_X1  g0282(.A(G244), .B1(new_n260), .B2(new_n261), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n265), .A2(new_n267), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT68), .B(G1698), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n272), .A2(new_n486), .A3(KEYINPUT4), .A4(G244), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G250), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G283), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n485), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n276), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT81), .B1(new_n493), .B2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT81), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n250), .A3(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(G45), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G1), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n494), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n256), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n251), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G257), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n492), .A2(G179), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n348), .B1(new_n492), .B2(new_n503), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n475), .A2(new_n481), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n474), .A2(new_n467), .A3(new_n472), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n296), .ZN(new_n508));
  INV_X1    g0308(.A(G190), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n492), .A2(new_n509), .A3(new_n503), .ZN(new_n510));
  AOI21_X1  g0310(.A(G200), .B1(new_n492), .B2(new_n503), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n508), .B(new_n480), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n300), .A2(new_n327), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n479), .A2(G87), .ZN(new_n515));
  INV_X1    g0315(.A(new_n415), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n224), .ZN(new_n517));
  XNOR2_X1  g0317(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n272), .A2(new_n224), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n365), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT19), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT82), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT19), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(G20), .B1(new_n526), .B2(new_n516), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G87), .A2(G97), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n527), .A2(new_n528), .B1(new_n463), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n224), .B1(new_n518), .B2(new_n415), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n521), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n514), .B(new_n515), .C1(new_n533), .C2(new_n395), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n268), .C2(new_n314), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n252), .A2(G45), .A3(G274), .ZN(new_n538));
  INV_X1    g0338(.A(G250), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n499), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(new_n276), .B1(new_n251), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT84), .B1(new_n541), .B2(G190), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(KEYINPUT84), .A3(G190), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n534), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n319), .B2(new_n541), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n262), .A2(G20), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G68), .B1(new_n518), .B2(new_n517), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n529), .A2(new_n463), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n531), .B2(KEYINPUT83), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n527), .A2(new_n528), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n296), .B1(new_n300), .B2(new_n327), .ZN(new_n553));
  INV_X1    g0353(.A(new_n327), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n479), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n553), .A2(new_n555), .B1(new_n278), .B2(new_n541), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G169), .B2(new_n541), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n513), .A2(new_n546), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n479), .A2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n298), .A2(G20), .A3(new_n463), .ZN(new_n560));
  XOR2_X1   g0360(.A(new_n560), .B(KEYINPUT25), .Z(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n535), .A2(G20), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n224), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n463), .A2(KEYINPUT23), .A3(G20), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT22), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n547), .A2(new_n569), .A3(G87), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n272), .A2(new_n224), .A3(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT22), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n395), .B1(new_n573), .B2(KEYINPUT24), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n562), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n268), .A2(new_n539), .ZN(new_n578));
  OAI211_X1 g0378(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n579));
  AND2_X1   g0379(.A1(KEYINPUT88), .A2(G294), .ZN(new_n580));
  NOR2_X1   g0380(.A1(KEYINPUT88), .A2(G294), .ZN(new_n581));
  OAI21_X1  g0381(.A(G33), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT89), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n272), .A2(new_n486), .A3(G250), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT89), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n579), .A4(new_n582), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n276), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n502), .A2(G264), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n500), .A2(new_n256), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(G179), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT90), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(new_n276), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n579), .A2(new_n582), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n595), .B2(new_n585), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n589), .B(new_n590), .C1(new_n594), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G169), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n592), .A3(G169), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n577), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n562), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n570), .A2(new_n572), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(KEYINPUT24), .A3(new_n567), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n296), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n602), .B1(new_n605), .B2(new_n574), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n597), .A2(G190), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n597), .A2(new_n319), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n276), .ZN(new_n611));
  OAI21_X1  g0411(.A(G257), .B1(new_n260), .B2(new_n261), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT85), .B1(new_n612), .B2(new_n484), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n272), .A2(new_n486), .A3(new_n614), .A4(G257), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g0416(.A(KEYINPUT86), .B(G303), .Z(new_n617));
  AOI22_X1  g0417(.A1(G264), .A2(new_n488), .B1(new_n617), .B2(new_n262), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n611), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n500), .A2(new_n251), .ZN(new_n620));
  INV_X1    g0420(.A(G270), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n590), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(KEYINPUT21), .B(G169), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n616), .A2(new_n618), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n276), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n501), .B1(new_n502), .B2(G270), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G179), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT20), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n490), .B(new_n224), .C1(G33), .C2(new_n476), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT87), .ZN(new_n631));
  INV_X1    g0431(.A(G116), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n296), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n629), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT87), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n630), .B(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(KEYINPUT20), .A3(new_n296), .A4(new_n633), .ZN(new_n638));
  OAI21_X1  g0438(.A(G116), .B1(new_n322), .B2(new_n478), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n299), .A2(new_n632), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n635), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(G169), .B1(new_n619), .B2(new_n622), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n628), .A2(new_n641), .B1(new_n643), .B2(KEYINPUT21), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n625), .A2(new_n626), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n319), .ZN(new_n646));
  INV_X1    g0446(.A(new_n381), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n645), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n641), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n558), .A2(new_n610), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n457), .A2(new_n650), .ZN(G372));
  INV_X1    g0451(.A(new_n311), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT95), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n454), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(KEYINPUT95), .B(new_n450), .C1(new_n452), .C2(new_n453), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n439), .ZN(new_n657));
  INV_X1    g0457(.A(new_n337), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n432), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n400), .A2(new_n386), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n379), .B(new_n402), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n652), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n506), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n546), .A2(new_n663), .A3(new_n557), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n541), .A2(new_n278), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n540), .A2(new_n251), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT91), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n540), .A2(KEYINPUT91), .A3(new_n251), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n537), .A2(new_n276), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n348), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n514), .B1(new_n533), .B2(new_n395), .ZN(new_n675));
  INV_X1    g0475(.A(new_n555), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n666), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT92), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n673), .B2(G200), .ZN(new_n679));
  AOI211_X1 g0479(.A(KEYINPUT92), .B(new_n319), .C1(new_n671), .C2(new_n672), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n545), .A2(new_n681), .B1(new_n556), .B2(new_n674), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n663), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n665), .A2(new_n677), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n544), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n553), .B(new_n515), .C1(new_n686), .C2(new_n542), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n679), .A2(new_n680), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n677), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n506), .A2(new_n512), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n689), .A2(new_n690), .A3(new_n609), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT93), .B1(new_n601), .B2(new_n644), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n591), .A2(new_n592), .B1(new_n597), .B2(G169), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n597), .A2(new_n592), .A3(G169), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n606), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n348), .B1(new_n625), .B2(new_n626), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n635), .A2(new_n638), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n639), .A2(new_n640), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT21), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n641), .B1(new_n623), .B2(new_n627), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n695), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n691), .A2(new_n692), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT94), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT94), .A4(new_n704), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n685), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n662), .B1(new_n457), .B2(new_n709), .ZN(G369));
  INV_X1    g0510(.A(new_n298), .ZN(new_n711));
  OR3_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .A3(G20), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT27), .B1(new_n711), .B2(G20), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n641), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n649), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n702), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G330), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n610), .B1(new_n577), .B2(new_n717), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n601), .A2(new_n716), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n601), .A2(new_n717), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n644), .A2(new_n717), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(G399));
  NOR2_X1   g0531(.A1(new_n216), .A2(G41), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n529), .A2(new_n463), .A3(new_n632), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT96), .ZN(new_n734));
  OR3_X1    g0534(.A1(new_n732), .A2(new_n252), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n732), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n227), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  INV_X1    g0538(.A(new_n627), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT97), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT97), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n588), .A2(new_n589), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n492), .A2(new_n503), .ZN(new_n743));
  INV_X1    g0543(.A(new_n541), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n740), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(G179), .B1(new_n671), .B2(new_n672), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n645), .A2(new_n597), .A3(new_n743), .A4(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n746), .B2(new_n747), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n716), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT31), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n752), .B(KEYINPUT31), .C1(new_n650), .C2(new_n716), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G330), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n707), .A2(new_n708), .ZN(new_n758));
  INV_X1    g0558(.A(new_n685), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n716), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT29), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT98), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n690), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n695), .A2(new_n702), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n689), .A2(new_n609), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n546), .A2(new_n683), .A3(new_n663), .A4(new_n557), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT26), .B1(new_n689), .B2(new_n506), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n767), .A2(new_n677), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n716), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT29), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n757), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT99), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n738), .B1(new_n773), .B2(G1), .ZN(G364));
  NOR2_X1   g0574(.A1(new_n215), .A2(G20), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G45), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT101), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(KEYINPUT101), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(G1), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n732), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n216), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n272), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT102), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G355), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n216), .A2(new_n272), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n247), .A2(new_n498), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n228), .A2(G45), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n785), .B(new_n789), .C1(G116), .C2(new_n782), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n223), .B1(G20), .B2(new_n348), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT103), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n781), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n224), .A2(G190), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n278), .A3(new_n319), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G159), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT32), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n509), .A2(G179), .A3(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n224), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G97), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n319), .A2(G179), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n798), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n262), .B1(new_n809), .B2(G107), .ZN(new_n810));
  INV_X1    g0610(.A(G87), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n807), .A2(G20), .A3(G190), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n806), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(G20), .A2(G179), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT104), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(new_n647), .A3(G200), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n509), .A3(G200), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n202), .A2(new_n816), .B1(new_n817), .B2(new_n365), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n802), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n815), .B(KEYINPUT105), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(new_n319), .A3(new_n647), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n820), .A2(new_n509), .A3(new_n319), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n819), .B1(new_n287), .B2(new_n821), .C1(new_n330), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n821), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G322), .ZN(new_n827));
  INV_X1    g0627(.A(G303), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n262), .B1(new_n812), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT106), .ZN(new_n830));
  INV_X1    g0630(.A(new_n816), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(G326), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G329), .A2(new_n800), .B1(new_n809), .B2(G283), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n580), .A2(new_n581), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n833), .B1(new_n835), .B2(new_n804), .ZN(new_n836));
  INV_X1    g0636(.A(new_n817), .ZN(new_n837));
  XNOR2_X1  g0637(.A(KEYINPUT33), .B(G317), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n827), .A2(new_n832), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n823), .B1(new_n825), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT107), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n791), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(new_n721), .ZN(new_n845));
  INV_X1    g0645(.A(new_n794), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n797), .B1(new_n843), .B2(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(G330), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT100), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n780), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n723), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n848), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n847), .B1(new_n851), .B2(new_n853), .ZN(G396));
  AOI22_X1  g0654(.A1(G132), .A2(new_n800), .B1(new_n809), .B2(G68), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n855), .B(new_n272), .C1(new_n202), .C2(new_n812), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G137), .A2(new_n831), .B1(new_n837), .B2(G150), .ZN(new_n857));
  INV_X1    g0657(.A(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n822), .B2(new_n858), .C1(new_n859), .C2(new_n821), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT34), .Z(new_n861));
  AOI211_X1 g0661(.A(new_n856), .B(new_n861), .C1(G58), .C2(new_n805), .ZN(new_n862));
  INV_X1    g0662(.A(G294), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n821), .A2(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n812), .A2(new_n463), .B1(new_n799), .B2(new_n824), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n808), .A2(new_n811), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n865), .A2(new_n272), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n806), .ZN(new_n868));
  INV_X1    g0668(.A(G283), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n868), .B1(new_n869), .B2(new_n817), .C1(new_n828), .C2(new_n816), .ZN(new_n870));
  INV_X1    g0670(.A(new_n822), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n864), .B(new_n870), .C1(G116), .C2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n791), .B1(new_n862), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n791), .A2(new_n792), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n781), .B1(new_n330), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n334), .B1(new_n333), .B2(new_n717), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n337), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n658), .A2(new_n717), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n873), .B(new_n875), .C1(new_n793), .C2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n760), .A2(new_n880), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n709), .A2(new_n716), .A3(new_n879), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n781), .B1(new_n885), .B2(new_n756), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n884), .A2(new_n757), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(G384));
  OR2_X1    g0688(.A1(new_n397), .A2(KEYINPUT16), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n391), .B1(new_n889), .B2(new_n398), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n353), .B2(new_n714), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n385), .A2(new_n377), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n389), .A2(new_n399), .ZN(new_n894));
  INV_X1    g0694(.A(new_n714), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n377), .A2(KEYINPUT108), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT108), .B1(new_n377), .B2(new_n895), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n378), .B(new_n894), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n893), .B1(new_n898), .B2(KEYINPUT37), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n890), .A2(new_n714), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n403), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(KEYINPUT109), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT109), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT108), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n399), .B2(new_n714), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n377), .A2(KEYINPUT108), .A3(new_n895), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n394), .A2(new_n398), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n353), .B1(new_n910), .B2(new_n356), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n892), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT37), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(new_n893), .B1(new_n403), .B2(new_n900), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n905), .B1(new_n915), .B2(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(KEYINPUT38), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n904), .A2(new_n916), .A3(KEYINPUT39), .A4(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n439), .A2(new_n716), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n914), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n403), .A2(new_n907), .A3(new_n908), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n918), .A2(new_n919), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n379), .A2(new_n402), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n714), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT110), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n414), .A2(new_n717), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n432), .A2(new_n439), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n432), .B2(new_n439), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n902), .A2(new_n903), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n925), .B1(new_n938), .B2(new_n905), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n904), .ZN(new_n940));
  INV_X1    g0740(.A(new_n878), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n937), .B(new_n940), .C1(new_n883), .C2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n930), .A2(new_n931), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n931), .B1(new_n930), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n761), .A2(new_n456), .A3(new_n771), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n662), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n945), .B(new_n947), .Z(new_n948));
  NOR2_X1   g0748(.A1(new_n936), .A2(new_n879), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n755), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(KEYINPUT40), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n940), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n924), .A2(new_n925), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT40), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n456), .A2(new_n755), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n722), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n948), .A2(new_n958), .B1(new_n252), .B2(new_n775), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n948), .B2(new_n958), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n227), .A2(new_n330), .A3(new_n366), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n202), .A2(G68), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n252), .B(G13), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n471), .ZN(new_n964));
  OAI211_X1 g0764(.A(G116), .B(new_n225), .C1(new_n964), .C2(KEYINPUT35), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(KEYINPUT35), .B2(new_n964), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT36), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n960), .A2(new_n963), .A3(new_n967), .ZN(G367));
  AOI22_X1  g0768(.A1(new_n786), .A2(new_n239), .B1(new_n216), .B2(new_n554), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n781), .B1(new_n796), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n534), .A2(new_n716), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n556), .B2(new_n674), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n689), .B2(new_n971), .ZN(new_n973));
  INV_X1    g0773(.A(new_n812), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G58), .A2(new_n974), .B1(new_n800), .B2(G137), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT112), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n859), .A2(new_n816), .B1(new_n817), .B2(new_n858), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n809), .A2(G77), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n272), .C1(new_n365), .C2(new_n804), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(G150), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n982), .B1(new_n202), .B2(new_n822), .C1(new_n983), .C2(new_n821), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n812), .A2(new_n632), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT46), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n824), .A2(new_n816), .B1(new_n817), .B2(new_n835), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n262), .B1(new_n808), .B2(new_n476), .C1(new_n988), .C2(new_n799), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n804), .A2(new_n463), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n986), .A2(new_n987), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n617), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n869), .B2(new_n822), .C1(new_n992), .C2(new_n821), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n984), .A2(KEYINPUT47), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n791), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT47), .B1(new_n984), .B2(new_n993), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n970), .B1(new_n973), .B2(new_n846), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n730), .A2(new_n728), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n716), .B1(new_n475), .B2(new_n481), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n763), .A2(new_n999), .B1(new_n663), .B2(new_n716), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT44), .Z(new_n1002));
  NOR2_X1   g0802(.A1(new_n998), .A2(new_n1000), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n727), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n729), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n730), .B1(new_n726), .B2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(new_n723), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n773), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n732), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n779), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n730), .B1(new_n998), .B2(new_n1000), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT42), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n763), .A2(new_n601), .A3(new_n999), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1019), .A2(new_n506), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1017), .B(new_n1018), .C1(new_n716), .C2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n973), .B(KEYINPUT111), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT43), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1025), .A3(new_n1023), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n727), .A2(new_n1000), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n997), .B1(new_n1014), .B2(new_n1031), .ZN(G387));
  INV_X1    g0832(.A(new_n1010), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n736), .B1(new_n773), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n773), .B2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n262), .B1(new_n808), .B2(new_n632), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n805), .A2(G283), .B1(new_n974), .B2(new_n834), .ZN(new_n1037));
  XOR2_X1   g0837(.A(KEYINPUT115), .B(G322), .Z(new_n1038));
  AOI22_X1  g0838(.A1(new_n831), .A2(new_n1038), .B1(new_n837), .B2(G311), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n822), .B2(new_n992), .C1(new_n988), .C2(new_n821), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1044));
  XNOR2_X1  g0844(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1036), .B(new_n1045), .C1(G326), .C2(new_n800), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n821), .A2(new_n202), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n272), .B1(new_n808), .B2(new_n476), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n812), .A2(new_n330), .B1(new_n799), .B2(new_n983), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n554), .C2(new_n805), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n858), .B2(new_n816), .C1(new_n290), .C2(new_n817), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1047), .B(new_n1051), .C1(G68), .C2(new_n871), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n791), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n784), .A2(new_n734), .B1(new_n463), .B2(new_n216), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G45), .B(new_n734), .C1(G68), .C2(G77), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n284), .A2(G50), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT114), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT50), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n236), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n786), .B1(new_n1061), .B2(new_n498), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1054), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n781), .B1(new_n1063), .B2(new_n796), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1053), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n724), .A2(new_n725), .A3(new_n794), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1065), .A2(new_n1066), .B1(new_n1033), .B2(new_n779), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1035), .A2(new_n1067), .ZN(G393));
  OAI22_X1  g0868(.A1(new_n821), .A2(new_n858), .B1(new_n983), .B2(new_n816), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n822), .A2(new_n284), .B1(new_n202), .B2(new_n817), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT117), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n812), .A2(new_n365), .B1(new_n799), .B2(new_n859), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n804), .A2(new_n330), .ZN(new_n1076));
  NOR4_X1   g0876(.A1(new_n1075), .A2(new_n1076), .A3(new_n262), .A4(new_n866), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1070), .A2(new_n1073), .A3(new_n1074), .A4(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT118), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT118), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n821), .A2(new_n824), .B1(new_n988), .B2(new_n816), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G283), .A2(new_n974), .B1(new_n800), .B2(new_n1038), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n272), .B1(new_n809), .B2(G107), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n632), .C2(new_n804), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n617), .B2(new_n837), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1082), .B(new_n1086), .C1(new_n863), .C2(new_n822), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1079), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n791), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n244), .A2(new_n216), .A3(new_n272), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n796), .B1(new_n476), .B2(new_n782), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n780), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n794), .B2(new_n1000), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1005), .B(new_n727), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n779), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n773), .A3(new_n1033), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n732), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1094), .B1(new_n773), .B2(new_n1033), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(G390));
  AOI21_X1  g0899(.A(new_n262), .B1(new_n800), .B2(G125), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n202), .B2(new_n808), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n974), .A2(G150), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G159), .C2(new_n805), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n826), .A2(G132), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT54), .B(G143), .Z(new_n1106));
  NAND2_X1  g0906(.A1(new_n871), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G128), .A2(new_n831), .B1(new_n837), .B2(G137), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n822), .A2(new_n476), .B1(new_n463), .B2(new_n817), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT122), .Z(new_n1111));
  OAI22_X1  g0911(.A1(new_n799), .A2(new_n863), .B1(new_n808), .B2(new_n365), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n262), .B1(new_n812), .B2(new_n811), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n1112), .A2(new_n1076), .A3(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1114), .B1(new_n869), .B2(new_n816), .C1(new_n821), .C2(new_n632), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1109), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1116), .A2(new_n791), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n874), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n780), .B1(new_n1118), .B2(new_n289), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n918), .A2(new_n926), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1117), .B(new_n1119), .C1(new_n1120), .C2(new_n792), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n919), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n941), .B1(new_n760), .B2(new_n880), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n936), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n766), .A2(new_n769), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n717), .A3(new_n877), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n936), .B1(new_n1128), .B2(new_n878), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1123), .B1(new_n924), .B2(new_n925), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1130), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n941), .B1(new_n770), .B2(new_n877), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(KEYINPUT119), .C1(new_n936), .C2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1125), .A2(new_n1120), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n755), .A2(G330), .A3(new_n949), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n607), .A2(new_n608), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n577), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n682), .A2(new_n513), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n703), .B1(new_n695), .B2(new_n702), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT94), .B1(new_n1142), .B2(new_n704), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n708), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n759), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n717), .A3(new_n880), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n936), .B1(new_n1146), .B2(new_n878), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1120), .B1(new_n1147), .B2(new_n919), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1136), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT120), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT120), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1153), .B(new_n1136), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1137), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n779), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1122), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n956), .A2(G330), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n946), .A3(new_n662), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n753), .A2(new_n754), .A3(G330), .A4(new_n880), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n936), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1136), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n941), .B2(new_n883), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(KEYINPUT121), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT121), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1165), .A3(new_n936), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n1133), .A3(new_n1136), .A4(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1159), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n1137), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n736), .B1(new_n1155), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1157), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G378));
  NAND2_X1  g0973(.A1(new_n955), .A2(G330), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  XOR2_X1   g0975(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n654), .A2(new_n311), .A3(new_n655), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n310), .A2(new_n714), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1179), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n654), .A2(new_n311), .A3(new_n655), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1177), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1177), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n943), .A2(new_n944), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1185), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n1183), .ZN(new_n1189));
  AOI221_X4 g0989(.A(new_n936), .B1(new_n939), .B2(new_n904), .C1(new_n1146), .C2(new_n878), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n927), .A2(new_n929), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT110), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n930), .A2(new_n931), .A3(new_n942), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1189), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1175), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1186), .B1(new_n943), .B2(new_n944), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1192), .A2(new_n1193), .A3(new_n1189), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1174), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n779), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n780), .B1(new_n1118), .B2(G50), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n262), .A2(new_n250), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n974), .B2(G77), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n287), .B2(new_n808), .C1(new_n869), .C2(new_n799), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT123), .Z(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n476), .B2(new_n817), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n816), .A2(new_n632), .B1(new_n365), .B2(new_n804), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n463), .A2(new_n821), .B1(new_n822), .B2(new_n327), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G50), .B1(new_n249), .B2(new_n250), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1208), .A2(KEYINPUT58), .B1(new_n1201), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n871), .A2(G137), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n826), .A2(G128), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n805), .A2(G150), .B1(new_n974), .B2(new_n1106), .ZN(new_n1213));
  INV_X1    g1013(.A(G132), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n817), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G125), .B2(new_n831), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1211), .A2(new_n1212), .A3(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(G33), .B(G41), .C1(new_n809), .C2(G159), .ZN(new_n1220));
  INV_X1    g1020(.A(G124), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n799), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1210), .B1(KEYINPUT58), .B2(new_n1208), .C1(new_n1219), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1200), .B1(new_n1223), .B2(new_n791), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1186), .B2(new_n793), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1199), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT125), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT57), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1153), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1150), .A2(KEYINPUT120), .A3(new_n1151), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1159), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1227), .B(new_n1228), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1159), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1169), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1238), .A2(KEYINPUT57), .A3(new_n1195), .A4(new_n1198), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n732), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1227), .B1(new_n1241), .B2(new_n1228), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1226), .B1(new_n1240), .B2(new_n1242), .ZN(G375));
  NAND2_X1  g1043(.A1(new_n936), .A2(new_n792), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n780), .B1(new_n1118), .B2(G68), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G294), .A2(new_n831), .B1(new_n837), .B2(G116), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n822), .B2(new_n463), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT126), .Z(new_n1248));
  NAND2_X1  g1048(.A1(new_n980), .A2(new_n262), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n812), .A2(new_n476), .B1(new_n799), .B2(new_n828), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT127), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1249), .B(new_n1251), .C1(new_n554), .C2(new_n805), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n869), .B2(new_n821), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n822), .A2(new_n983), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G128), .A2(new_n800), .B1(new_n974), .B2(G159), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n262), .B1(new_n809), .B2(G58), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n202), .C2(new_n804), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G132), .B2(new_n831), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n826), .A2(G137), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n837), .A2(new_n1106), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1248), .A2(new_n1253), .B1(new_n1254), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1245), .B1(new_n1262), .B2(new_n791), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1233), .A2(new_n779), .B1(new_n1244), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1170), .A2(new_n1013), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1237), .A2(new_n1233), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(G381));
  OR2_X1    g1067(.A1(G375), .A2(G378), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G387), .A2(G390), .ZN(new_n1270));
  INV_X1    g1070(.A(G396), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1035), .A2(new_n1271), .A3(new_n1067), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1272), .A2(G384), .A3(G381), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1270), .A3(new_n1273), .ZN(G407));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(G343), .C2(new_n1268), .ZN(G409));
  AND2_X1   g1075(.A1(new_n715), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1266), .A2(new_n1277), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1237), .A2(new_n1233), .A3(KEYINPUT60), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n732), .B(new_n1170), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1264), .ZN(new_n1281));
  INV_X1    g1081(.A(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(G384), .A3(new_n1264), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1226), .C1(new_n1240), .C2(new_n1242), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1226), .B1(new_n1012), .B2(new_n1241), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1172), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1276), .B(new_n1285), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1276), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1276), .A2(G2897), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1285), .B(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT63), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G393), .A2(G396), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1272), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G387), .A2(G390), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1298), .B1(new_n1300), .B2(new_n1270), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1270), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1297), .A3(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1301), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n1289), .B2(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1295), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1285), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1291), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1304), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1291), .B2(new_n1309), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1307), .B1(new_n1313), .B2(new_n1315), .ZN(G405));
  XNOR2_X1  g1116(.A(new_n1314), .B(new_n1285), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G375), .A2(G378), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1317), .B1(new_n1269), .B2(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1314), .B(new_n1309), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1268), .A3(new_n1318), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(G402));
endmodule


