

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  NOR2_X1 U322 ( .A1(n488), .A2(n578), .ZN(n413) );
  INV_X1 U323 ( .A(KEYINPUT83), .ZN(n369) );
  XOR2_X1 U324 ( .A(KEYINPUT28), .B(n471), .Z(n514) );
  INV_X1 U325 ( .A(KEYINPUT33), .ZN(n424) );
  INV_X1 U326 ( .A(KEYINPUT100), .ZN(n412) );
  XOR2_X1 U327 ( .A(G190GAT), .B(KEYINPUT73), .Z(n352) );
  XNOR2_X1 U328 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U329 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U330 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U331 ( .A(G218GAT), .B(G162GAT), .Z(n364) );
  XNOR2_X1 U332 ( .A(n372), .B(n371), .ZN(n375) );
  NOR2_X1 U333 ( .A1(n391), .A2(n390), .ZN(n488) );
  XOR2_X1 U334 ( .A(n431), .B(n430), .Z(n574) );
  NOR2_X1 U335 ( .A1(n530), .A2(n473), .ZN(n562) );
  XOR2_X1 U336 ( .A(KEYINPUT108), .B(n480), .Z(n525) );
  XNOR2_X1 U337 ( .A(n446), .B(n445), .ZN(n503) );
  XNOR2_X1 U338 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U339 ( .A(n481), .B(G106GAT), .ZN(n482) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n447) );
  XNOR2_X1 U341 ( .A(n477), .B(n476), .ZN(G1349GAT) );
  XNOR2_X1 U342 ( .A(n448), .B(n447), .ZN(G1330GAT) );
  XNOR2_X1 U343 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n446) );
  XNOR2_X1 U344 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n290) );
  XNOR2_X1 U345 ( .A(n290), .B(G29GAT), .ZN(n291) );
  XOR2_X1 U346 ( .A(n291), .B(KEYINPUT8), .Z(n293) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G50GAT), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n444) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .ZN(n430) );
  XNOR2_X1 U350 ( .A(n430), .B(n352), .ZN(n295) );
  NAND2_X1 U351 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U353 ( .A(KEYINPUT11), .B(G92GAT), .Z(n297) );
  XNOR2_X1 U354 ( .A(G134GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U356 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U357 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n301) );
  XNOR2_X1 U358 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n364), .B(n302), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n444), .B(n305), .ZN(n563) );
  INV_X1 U363 ( .A(n563), .ZN(n484) );
  XNOR2_X1 U364 ( .A(KEYINPUT36), .B(n484), .ZN(n583) );
  XOR2_X1 U365 ( .A(KEYINPUT81), .B(KEYINPUT17), .Z(n307) );
  XNOR2_X1 U366 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U368 ( .A(KEYINPUT19), .B(n308), .Z(n356) );
  XOR2_X1 U369 ( .A(G127GAT), .B(KEYINPUT0), .Z(n310) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n323) );
  XOR2_X1 U372 ( .A(G120GAT), .B(G71GAT), .Z(n429) );
  XOR2_X1 U373 ( .A(n323), .B(n429), .Z(n312) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G99GAT), .ZN(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U376 ( .A(KEYINPUT20), .B(KEYINPUT65), .Z(n314) );
  NAND2_X1 U377 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U379 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U380 ( .A(G176GAT), .B(KEYINPUT80), .Z(n318) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(G190GAT), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U383 ( .A(G15GAT), .B(n319), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n356), .B(n322), .ZN(n530) );
  INV_X1 U386 ( .A(n530), .ZN(n524) );
  XOR2_X1 U387 ( .A(n323), .B(KEYINPUT88), .Z(n325) );
  NAND2_X1 U388 ( .A1(G225GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U390 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n327) );
  XNOR2_X1 U391 ( .A(KEYINPUT87), .B(KEYINPUT6), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U394 ( .A(G57GAT), .B(G148GAT), .Z(n331) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(G1GAT), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U398 ( .A(G85GAT), .B(G162GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n334), .B(KEYINPUT2), .ZN(n373) );
  XNOR2_X1 U401 ( .A(G29GAT), .B(n373), .ZN(n335) );
  XNOR2_X1 U402 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U403 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U404 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n340) );
  XNOR2_X1 U405 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(n341), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n519) );
  XOR2_X1 U409 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n345) );
  NAND2_X1 U410 ( .A1(G226GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U411 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U412 ( .A(n346), .B(KEYINPUT93), .Z(n351) );
  XOR2_X1 U413 ( .A(G211GAT), .B(KEYINPUT84), .Z(n348) );
  XNOR2_X1 U414 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n348), .B(n347), .ZN(n378) );
  XNOR2_X1 U416 ( .A(G176GAT), .B(G92GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n349), .B(G64GAT), .ZN(n419) );
  XNOR2_X1 U418 ( .A(n378), .B(n419), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n360) );
  XOR2_X1 U420 ( .A(KEYINPUT92), .B(n352), .Z(n354) );
  XOR2_X1 U421 ( .A(G169GAT), .B(G8GAT), .Z(n439) );
  XNOR2_X1 U422 ( .A(n439), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U424 ( .A(n355), .B(G218GAT), .Z(n358) );
  XNOR2_X1 U425 ( .A(G36GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X2 U427 ( .A(n360), .B(n359), .Z(n522) );
  XNOR2_X1 U428 ( .A(n522), .B(KEYINPUT96), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n361), .B(KEYINPUT27), .ZN(n386) );
  NAND2_X1 U430 ( .A1(n519), .A2(n386), .ZN(n543) );
  XOR2_X1 U431 ( .A(KEYINPUT85), .B(KEYINPUT24), .Z(n363) );
  XNOR2_X1 U432 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U434 ( .A(KEYINPUT86), .B(n364), .Z(n366) );
  XOR2_X1 U435 ( .A(G141GAT), .B(G22GAT), .Z(n440) );
  XNOR2_X1 U436 ( .A(G50GAT), .B(n440), .ZN(n365) );
  XNOR2_X1 U437 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U438 ( .A(n368), .B(n367), .Z(n372) );
  NAND2_X1 U439 ( .A1(G228GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n373), .B(KEYINPUT82), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U442 ( .A(G78GAT), .B(G148GAT), .Z(n377) );
  XNOR2_X1 U443 ( .A(G106GAT), .B(G204GAT), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n420) );
  XOR2_X1 U445 ( .A(n378), .B(n420), .Z(n379) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n471) );
  NOR2_X1 U447 ( .A1(n543), .A2(n514), .ZN(n528) );
  XNOR2_X1 U448 ( .A(KEYINPUT97), .B(n528), .ZN(n381) );
  NOR2_X1 U449 ( .A1(n524), .A2(n381), .ZN(n391) );
  NAND2_X1 U450 ( .A1(n522), .A2(n524), .ZN(n382) );
  NAND2_X1 U451 ( .A1(n382), .A2(n471), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n383), .B(KEYINPUT25), .ZN(n384) );
  XNOR2_X1 U453 ( .A(KEYINPUT98), .B(n384), .ZN(n388) );
  NOR2_X1 U454 ( .A1(n524), .A2(n471), .ZN(n385) );
  XNOR2_X1 U455 ( .A(KEYINPUT26), .B(n385), .ZN(n567) );
  AND2_X1 U456 ( .A1(n386), .A2(n567), .ZN(n387) );
  NOR2_X1 U457 ( .A1(n388), .A2(n387), .ZN(n389) );
  NOR2_X1 U458 ( .A1(n519), .A2(n389), .ZN(n390) );
  XOR2_X1 U459 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n393) );
  XNOR2_X1 U460 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U462 ( .A(KEYINPUT13), .B(G57GAT), .Z(n423) );
  XOR2_X1 U463 ( .A(n423), .B(G71GAT), .Z(n396) );
  XNOR2_X1 U464 ( .A(G15GAT), .B(G1GAT), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n394), .B(KEYINPUT67), .ZN(n432) );
  XNOR2_X1 U466 ( .A(n432), .B(G183GAT), .ZN(n395) );
  XNOR2_X1 U467 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(n397), .ZN(n411) );
  XOR2_X1 U469 ( .A(G155GAT), .B(G211GAT), .Z(n400) );
  XNOR2_X1 U470 ( .A(G22GAT), .B(G127GAT), .ZN(n399) );
  XNOR2_X1 U471 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U472 ( .A(KEYINPUT77), .B(G64GAT), .Z(n402) );
  XNOR2_X1 U473 ( .A(G8GAT), .B(G78GAT), .ZN(n401) );
  XNOR2_X1 U474 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U475 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U476 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n406) );
  NAND2_X1 U477 ( .A1(G231GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U478 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U479 ( .A(KEYINPUT12), .B(n407), .ZN(n408) );
  XNOR2_X1 U480 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n411), .B(n410), .ZN(n460) );
  INV_X1 U482 ( .A(n460), .ZN(n578) );
  XNOR2_X1 U483 ( .A(n413), .B(n412), .ZN(n414) );
  NOR2_X1 U484 ( .A1(n583), .A2(n414), .ZN(n415) );
  XOR2_X1 U485 ( .A(KEYINPUT37), .B(n415), .Z(n479) );
  XOR2_X1 U486 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n417) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U488 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U489 ( .A(n418), .B(KEYINPUT69), .Z(n422) );
  XNOR2_X1 U490 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n423), .B(KEYINPUT70), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U494 ( .A(n432), .B(KEYINPUT66), .Z(n434) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U497 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n436) );
  XNOR2_X1 U498 ( .A(G113GAT), .B(G197GAT), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U500 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n568) );
  XNOR2_X1 U504 ( .A(KEYINPUT68), .B(n568), .ZN(n558) );
  INV_X1 U505 ( .A(n558), .ZN(n463) );
  NOR2_X1 U506 ( .A1(n574), .A2(n463), .ZN(n489) );
  NAND2_X1 U507 ( .A1(n479), .A2(n489), .ZN(n445) );
  NAND2_X1 U508 ( .A1(n503), .A2(n524), .ZN(n448) );
  XOR2_X1 U509 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n469) );
  XNOR2_X1 U510 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n449), .B(n574), .ZN(n478) );
  INV_X1 U512 ( .A(n478), .ZN(n550) );
  NAND2_X1 U513 ( .A1(n550), .A2(n568), .ZN(n454) );
  INV_X1 U514 ( .A(n454), .ZN(n452) );
  XOR2_X1 U515 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n450) );
  XNOR2_X1 U516 ( .A(KEYINPUT112), .B(n450), .ZN(n453) );
  INV_X1 U517 ( .A(n453), .ZN(n451) );
  NAND2_X1 U518 ( .A1(n452), .A2(n451), .ZN(n456) );
  NAND2_X1 U519 ( .A1(n454), .A2(n453), .ZN(n455) );
  NAND2_X1 U520 ( .A1(n456), .A2(n455), .ZN(n458) );
  NOR2_X1 U521 ( .A1(n563), .A2(n578), .ZN(n457) );
  AND2_X1 U522 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U523 ( .A(n459), .B(KEYINPUT47), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n460), .A2(n583), .ZN(n461) );
  XOR2_X1 U525 ( .A(KEYINPUT45), .B(n461), .Z(n462) );
  NOR2_X1 U526 ( .A1(n574), .A2(n462), .ZN(n464) );
  NAND2_X1 U527 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U529 ( .A(KEYINPUT48), .B(n467), .ZN(n545) );
  NAND2_X1 U530 ( .A1(n545), .A2(n522), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n470), .A2(n519), .ZN(n566) );
  AND2_X1 U533 ( .A1(n566), .A2(n471), .ZN(n472) );
  XNOR2_X1 U534 ( .A(KEYINPUT55), .B(n472), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n562), .A2(n550), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n475) );
  XOR2_X1 U537 ( .A(G176GAT), .B(KEYINPUT123), .Z(n474) );
  NOR2_X1 U538 ( .A1(n478), .A2(n568), .ZN(n506) );
  NAND2_X1 U539 ( .A1(n506), .A2(n479), .ZN(n480) );
  NAND2_X1 U540 ( .A1(n525), .A2(n514), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n481) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1339GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n491) );
  XOR2_X1 U544 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n486) );
  NAND2_X1 U545 ( .A1(n484), .A2(n578), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  NOR2_X1 U547 ( .A1(n488), .A2(n487), .ZN(n505) );
  AND2_X1 U548 ( .A1(n489), .A2(n505), .ZN(n496) );
  NAND2_X1 U549 ( .A1(n496), .A2(n519), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U552 ( .A1(n496), .A2(n522), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U555 ( .A1(n496), .A2(n524), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U557 ( .A1(n514), .A2(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n499) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n501) );
  NAND2_X1 U562 ( .A1(n503), .A2(n519), .ZN(n500) );
  XOR2_X1 U563 ( .A(n501), .B(n500), .Z(G1328GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n522), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n503), .A2(n514), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U568 ( .A1(n506), .A2(n505), .ZN(n515) );
  NAND2_X1 U569 ( .A1(n515), .A2(n519), .ZN(n510) );
  XOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n508) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n515), .A2(n522), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n515), .A2(n524), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  XOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT109), .Z(n521) );
  NAND2_X1 U584 ( .A1(n519), .A2(n525), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n525), .A2(n522), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(KEYINPUT110), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n545), .A2(n528), .ZN(n529) );
  NOR2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n539), .A2(n558), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n531), .B(KEYINPUT114), .ZN(n532) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U597 ( .A1(n539), .A2(n550), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U599 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n537) );
  NAND2_X1 U601 ( .A1(n539), .A2(n578), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n538), .Z(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U605 ( .A1(n539), .A2(n563), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U607 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  XOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT119), .Z(n549) );
  INV_X1 U609 ( .A(n567), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(n547), .Z(n556) );
  NAND2_X1 U613 ( .A1(n556), .A2(n568), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U617 ( .A1(n556), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n556), .A2(n578), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n563), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n562), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT122), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n578), .A2(n562), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n570) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n582) );
  INV_X1 U634 ( .A(n582), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n579), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(n571), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U641 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

