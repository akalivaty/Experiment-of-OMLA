//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n438, new_n439, new_n444, new_n445, new_n446, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n551, new_n552, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n588,
    new_n591, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(G69), .ZN(new_n438));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(G69), .ZN(new_n439));
  NOR2_X1   g014(.A1(new_n438), .A2(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT68), .ZN(new_n456));
  XOR2_X1   g031(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n457));
  XNOR2_X1  g032(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  NAND2_X1  g037(.A1(new_n458), .A2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G567), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g041(.A(new_n466), .B(KEYINPUT70), .Z(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(G319));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n470), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(new_n470), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n472), .A2(G136), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n469), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n470), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n480), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n492), .B(new_n497), .C1(new_n494), .C2(new_n493), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n490), .B1(new_n496), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n500), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n512), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  AND2_X1   g093(.A1(new_n508), .A2(new_n512), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n513), .A2(G51), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n520), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  AOI22_X1  g101(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n510), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n515), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G171));
  AOI22_X1  g107(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n510), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n519), .A2(G81), .B1(G43), .B2(new_n513), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT72), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(G860), .A3(new_n539), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(G188));
  AOI22_X1  g119(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n510), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n513), .A2(G53), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT9), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n519), .A2(G91), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(G299));
  OR3_X1    g125(.A1(new_n528), .A2(new_n531), .A3(KEYINPUT73), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT73), .B1(new_n528), .B2(new_n531), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(G301));
  OR2_X1    g128(.A1(new_n511), .A2(new_n517), .ZN(G303));
  INV_X1    g129(.A(G74), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n510), .B1(new_n507), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(G49), .B2(new_n513), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n505), .A2(G87), .A3(new_n506), .A4(new_n512), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G288));
  NAND2_X1  g135(.A1(new_n513), .A2(G48), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n505), .A2(G86), .A3(new_n506), .A4(new_n512), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n505), .A2(G61), .A3(new_n506), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n510), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G305));
  NAND2_X1  g144(.A1(new_n513), .A2(G47), .ZN(new_n570));
  INV_X1    g145(.A(G85), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n515), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n572), .A2(KEYINPUT75), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n572), .A2(KEYINPUT75), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n573), .A2(new_n574), .B1(new_n510), .B2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(new_n519), .A2(G92), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT10), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n507), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  MUX2_X1   g159(.A(new_n584), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g160(.A(new_n584), .B(G301), .S(G868), .Z(G321));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(G299), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n587), .B2(G168), .ZN(G297));
  OAI21_X1  g164(.A(new_n588), .B1(new_n587), .B2(G168), .ZN(G280));
  INV_X1    g165(.A(new_n584), .ZN(new_n591));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n537), .A2(new_n539), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  MUX2_X1   g170(.A(new_n594), .B(new_n595), .S(G868), .Z(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g172(.A1(new_n469), .A2(new_n473), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT12), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT13), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(G2100), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT76), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n481), .A2(G123), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT77), .Z(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OR2_X1    g181(.A1(new_n606), .A2(KEYINPUT78), .ZN(new_n607));
  INV_X1    g182(.A(G111), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n606), .A2(KEYINPUT78), .B1(new_n608), .B2(G2105), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n472), .A2(G135), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G2096), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(new_n612), .B1(new_n601), .B2(G2100), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n603), .B(new_n613), .C1(new_n612), .C2(new_n611), .ZN(G156));
  XNOR2_X1  g189(.A(G2427), .B(G2438), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2430), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(KEYINPUT14), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G1341), .B(G1348), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n620), .B(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G2443), .B(G2446), .Z(new_n626));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(G14), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n625), .ZN(G401));
  NOR2_X1   g206(.A1(G2072), .A2(G2078), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n446), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT17), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT80), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2084), .B(G2090), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n635), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT82), .Z(new_n641));
  OAI21_X1  g216(.A(KEYINPUT81), .B1(new_n446), .B2(new_n632), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n446), .A2(KEYINPUT81), .A3(new_n632), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n637), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(new_n639), .C1(new_n634), .C2(new_n637), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n637), .A2(new_n633), .A3(new_n639), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2096), .B(G2100), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1971), .B(G1976), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT19), .ZN(new_n652));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT83), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n653), .A2(new_n654), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(new_n656), .ZN(new_n662));
  MUX2_X1   g237(.A(new_n662), .B(new_n661), .S(new_n652), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1991), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G229));
  INV_X1    g246(.A(G29), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(G32), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n472), .A2(G141), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n481), .A2(G129), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n473), .A2(G105), .ZN(new_n676));
  NAND3_X1  g251(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT26), .Z(new_n678));
  NAND4_X1  g253(.A1(new_n674), .A2(new_n675), .A3(new_n676), .A4(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n673), .B1(new_n679), .B2(G29), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT27), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT97), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT31), .B(G11), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(KEYINPUT98), .ZN(new_n686));
  INV_X1    g261(.A(G28), .ZN(new_n687));
  AOI21_X1  g262(.A(G29), .B1(new_n687), .B2(KEYINPUT30), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(KEYINPUT30), .B2(new_n687), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT98), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n684), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT85), .B(G29), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n686), .B(new_n691), .C1(new_n611), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n680), .A2(new_n682), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G1961), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NOR2_X1   g273(.A1(G171), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G5), .B2(new_n698), .ZN(new_n700));
  AOI211_X1 g275(.A(new_n683), .B(new_n696), .C1(new_n697), .C2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n672), .A2(G33), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT25), .ZN(new_n703));
  NAND2_X1  g278(.A1(G103), .A2(G2104), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n470), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n472), .A2(G139), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n470), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT95), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n702), .B1(new_n710), .B2(G29), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(new_n444), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT96), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n698), .A2(G21), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G168), .B2(new_n698), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1966), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT24), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G34), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n692), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n477), .B2(new_n672), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(G2084), .Z(new_n722));
  NOR2_X1   g297(.A1(new_n693), .A2(G27), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n693), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2078), .ZN(new_n725));
  NOR3_X1   g300(.A1(new_n716), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n700), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n727), .A2(G1961), .B1(new_n444), .B2(new_n711), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n701), .A2(new_n713), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n729), .A2(KEYINPUT99), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(KEYINPUT99), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n692), .A2(G26), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(G128), .A2(new_n481), .B1(new_n472), .B2(G140), .ZN(new_n735));
  NOR2_X1   g310(.A1(G104), .A2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(new_n470), .B2(G116), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(new_n672), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT94), .B(G2067), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n693), .A2(G35), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n693), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT29), .B(G2090), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n591), .A2(G16), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G4), .B2(G16), .ZN(new_n750));
  INV_X1    g325(.A(G1348), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n744), .B(new_n748), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n698), .A2(G20), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT23), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n752), .B(new_n756), .C1(new_n751), .C2(new_n750), .ZN(new_n757));
  MUX2_X1   g332(.A(G19), .B(new_n594), .S(G16), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1341), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n730), .A2(new_n731), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G22), .ZN(new_n761));
  OR3_X1    g336(.A1(new_n761), .A2(KEYINPUT89), .A3(G16), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT89), .B1(new_n761), .B2(G16), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n762), .B(new_n763), .C1(G166), .C2(new_n698), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT90), .B(G1971), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT33), .B(G1976), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT88), .ZN(new_n768));
  INV_X1    g343(.A(G288), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n766), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n768), .B2(new_n771), .ZN(new_n773));
  MUX2_X1   g348(.A(G6), .B(G305), .S(G16), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT32), .ZN(new_n775));
  INV_X1    g350(.A(G1981), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT34), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT34), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n773), .A2(new_n780), .A3(new_n777), .ZN(new_n781));
  MUX2_X1   g356(.A(G24), .B(G290), .S(G16), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G1986), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(G1986), .ZN(new_n784));
  OR2_X1    g359(.A1(G95), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n786));
  INV_X1    g361(.A(G131), .ZN(new_n787));
  INV_X1    g362(.A(G119), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n786), .B1(new_n471), .B2(new_n787), .C1(new_n788), .C2(new_n480), .ZN(new_n789));
  MUX2_X1   g364(.A(G25), .B(new_n789), .S(new_n693), .Z(new_n790));
  XOR2_X1   g365(.A(KEYINPUT35), .B(G1991), .Z(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n790), .B(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(KEYINPUT91), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n784), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n795), .A2(KEYINPUT91), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n760), .A2(new_n800), .A3(new_n801), .ZN(G311));
  NAND3_X1  g377(.A1(new_n760), .A2(new_n800), .A3(new_n801), .ZN(G150));
  NOR2_X1   g378(.A1(new_n584), .A2(new_n592), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n510), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT101), .B(G55), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n513), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n515), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n536), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n594), .B2(new_n813), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n806), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n817));
  AOI21_X1  g392(.A(G860), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n813), .A2(G860), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT102), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n819), .A2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(new_n477), .B(new_n485), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n611), .B(new_n824), .Z(new_n825));
  INV_X1    g400(.A(KEYINPUT103), .ZN(new_n826));
  INV_X1    g401(.A(new_n498), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n497), .B1(new_n469), .B2(new_n492), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n496), .A2(KEYINPUT103), .A3(new_n498), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n490), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n741), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n679), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n710), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n709), .B2(new_n833), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n789), .B(new_n599), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n472), .A2(G142), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT104), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n481), .A2(G130), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n470), .A2(G118), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n836), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n835), .A2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n825), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  INV_X1    g423(.A(new_n825), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n844), .B(new_n849), .C1(new_n846), .C2(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n835), .A2(KEYINPUT105), .A3(new_n843), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n847), .B(new_n848), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g429(.A1(new_n584), .A2(G299), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n548), .A2(new_n549), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n579), .A2(new_n546), .A3(new_n856), .A4(new_n583), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(KEYINPUT41), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT41), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n595), .B(new_n815), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n857), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n864), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT42), .ZN(new_n866));
  XNOR2_X1  g441(.A(G290), .B(G166), .ZN(new_n867));
  XOR2_X1   g442(.A(G288), .B(G305), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n862), .B(new_n871), .C1(new_n864), .C2(new_n861), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n866), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n870), .B1(new_n866), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(G868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n813), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(G868), .B2(new_n876), .ZN(G295));
  OAI21_X1  g452(.A(new_n875), .B1(G868), .B2(new_n876), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n879));
  NAND3_X1  g454(.A1(G301), .A2(new_n879), .A3(G168), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(G171), .B2(G286), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n551), .A2(new_n552), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(G286), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n815), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n883), .ZN(new_n887));
  INV_X1    g462(.A(new_n815), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n880), .A2(new_n815), .A3(KEYINPUT107), .A4(new_n883), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n886), .A2(new_n889), .A3(new_n864), .A4(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n858), .A2(new_n859), .ZN(new_n892));
  INV_X1    g467(.A(new_n884), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n815), .B1(new_n883), .B2(new_n880), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n895), .A3(new_n869), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n848), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n870), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT43), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n886), .A2(new_n889), .A3(new_n890), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n892), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n889), .A2(new_n864), .A3(new_n884), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n869), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n905), .A2(new_n897), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT44), .B1(new_n901), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n906), .B1(new_n898), .B2(new_n900), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n905), .A2(new_n897), .A3(KEYINPUT43), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(G397));
  INV_X1    g488(.A(new_n490), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n496), .A2(KEYINPUT103), .A3(new_n498), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT103), .B1(new_n496), .B2(new_n498), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT45), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n474), .A2(new_n476), .A3(G40), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(G290), .A2(G1986), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(G290), .A2(G1986), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G2067), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n741), .B(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT109), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n929), .B2(new_n679), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(G1996), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n921), .A2(G1996), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT108), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n930), .A2(new_n931), .B1(new_n679), .B2(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n936));
  INV_X1    g511(.A(new_n791), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n789), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n789), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n922), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND4_X1   g515(.A1(new_n926), .A2(new_n935), .A3(new_n936), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n942));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n943));
  NOR3_X1   g518(.A1(G164), .A2(new_n943), .A3(G1384), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT111), .B1(new_n831), .B2(G1384), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n917), .A2(new_n946), .A3(new_n918), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n944), .B1(new_n948), .B2(new_n943), .ZN(new_n949));
  INV_X1    g524(.A(new_n920), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n697), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT45), .B1(new_n945), .B2(new_n947), .ZN(new_n952));
  NOR2_X1   g527(.A1(G164), .A2(G1384), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n920), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(G2078), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n917), .A2(KEYINPUT45), .A3(new_n918), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(G164), .B2(G1384), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n960), .A2(new_n962), .A3(new_n445), .A4(new_n920), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT124), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n957), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n957), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT124), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n951), .A2(new_n959), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n882), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT50), .B1(new_n945), .B2(new_n947), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n920), .B1(new_n970), .B2(new_n944), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n971), .A2(new_n697), .B1(KEYINPUT124), .B2(new_n966), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n919), .A2(new_n957), .A3(G2078), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(new_n920), .A3(new_n960), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n972), .A2(G301), .A3(new_n974), .A4(new_n965), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n942), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1966), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n952), .B2(new_n955), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n950), .A2(G2084), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n970), .B2(new_n944), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT112), .B(G8), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(G168), .A2(new_n982), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(KEYINPUT51), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n978), .B2(new_n980), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT51), .B1(new_n989), .B2(new_n985), .ZN(new_n990));
  AOI211_X1 g565(.A(G168), .B(new_n982), .C1(new_n978), .C2(new_n980), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n976), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n945), .A2(new_n947), .A3(new_n920), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n769), .A2(G1976), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n995), .A3(new_n983), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT52), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n994), .A2(new_n995), .A3(new_n999), .A4(new_n983), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n564), .A2(new_n776), .A3(new_n568), .ZN(new_n1001));
  OAI21_X1  g576(.A(G1981), .B1(new_n563), .B2(new_n567), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1001), .A2(KEYINPUT49), .A3(new_n1002), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n994), .A3(new_n983), .A4(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n997), .A2(new_n1000), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT114), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n997), .A2(new_n1010), .A3(new_n1000), .A4(new_n1007), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT55), .Z(new_n1014));
  AND3_X1   g589(.A1(new_n960), .A2(new_n920), .A3(new_n962), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n971), .A2(G2090), .B1(G1971), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1016), .A3(G8), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n943), .B1(new_n945), .B2(new_n947), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n953), .A2(new_n943), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n920), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1018), .A2(new_n1020), .A3(G2090), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1015), .A2(G1971), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n983), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1013), .B(KEYINPUT55), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT125), .B1(new_n1012), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT125), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n1017), .A4(new_n1025), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n972), .A2(new_n965), .A3(new_n974), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G171), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(KEYINPUT54), .C1(new_n882), .C2(new_n968), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n993), .A2(new_n1027), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n831), .A2(KEYINPUT111), .A3(G1384), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n946), .B1(new_n917), .B2(new_n918), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n943), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n944), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1348), .B1(new_n1039), .B2(new_n920), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n945), .A2(new_n947), .A3(new_n927), .A4(new_n920), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT116), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT117), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1041), .B(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n971), .A2(new_n751), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n591), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n548), .B2(KEYINPUT115), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G299), .B(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1956), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1015), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1049), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT118), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1059), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n1061), .B(new_n1062), .C1(new_n1049), .C2(new_n1057), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1062), .A2(new_n1056), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT119), .B(G1996), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1015), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n994), .A2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n1071), .C2(new_n594), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n594), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n1075), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT121), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1066), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1048), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1047), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT60), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1043), .A2(new_n1085), .A3(new_n1048), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n591), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1065), .B1(new_n1062), .B2(new_n1056), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT122), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n1065), .C1(new_n1062), .C2(new_n1056), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT60), .B(new_n584), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1081), .A2(new_n1087), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1034), .B1(new_n1064), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n984), .A2(G286), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1028), .A2(new_n1017), .A3(new_n1025), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT63), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1016), .A2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1024), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1008), .A2(new_n1098), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1101), .A2(new_n1096), .A3(new_n1017), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1007), .A2(new_n998), .A3(new_n769), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1001), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n994), .A3(new_n983), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1017), .B2(new_n1008), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n992), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n987), .B(KEYINPUT62), .C1(new_n990), .C2(new_n991), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n882), .A3(new_n968), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1104), .B(new_n1110), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n941), .B1(new_n1095), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n924), .A2(new_n922), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT48), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n935), .A2(new_n936), .A3(new_n940), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT46), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n933), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(new_n930), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n933), .A2(new_n1121), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(KEYINPUT126), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(KEYINPUT126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1123), .B(new_n1124), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1125), .B(KEYINPUT126), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1124), .B1(new_n1130), .B2(new_n1123), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1120), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n741), .A2(new_n927), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n921), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1117), .A2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g712(.A1(G229), .A2(new_n467), .A3(G401), .A4(G227), .ZN(new_n1139));
  OAI211_X1 g713(.A(new_n853), .B(new_n1139), .C1(new_n910), .C2(new_n911), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


