//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT65), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n469), .B1(new_n467), .B2(new_n462), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n467), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT64), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(G113), .A2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n474), .B1(new_n485), .B2(new_n473), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  XOR2_X1   g062(.A(KEYINPUT65), .B(G2104), .Z(new_n488));
  AOI22_X1  g063(.A1(new_n488), .A2(KEYINPUT3), .B1(new_n465), .B2(new_n468), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n489), .B2(new_n473), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n470), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(G124), .A2(new_n492), .B1(new_n497), .B2(G136), .ZN(new_n498));
  OR2_X1    g073(.A1(G100), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  AOI21_X1  g077(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT4), .B1(new_n503), .B2(G138), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n469), .B(G126), .C1(new_n467), .C2(new_n462), .ZN(new_n505));
  NAND2_X1  g080(.A1(G114), .A2(G2104), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n473), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT4), .A2(G138), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n469), .B(new_n508), .C1(new_n467), .C2(new_n462), .ZN(new_n509));
  NAND2_X1  g084(.A1(G102), .A2(G2104), .ZN(new_n510));
  AOI21_X1  g085(.A(G2105), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n504), .A2(new_n507), .A3(new_n511), .ZN(G164));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n513), .A2(new_n514), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT69), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n518), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G166));
  NAND2_X1  g109(.A1(new_n517), .A2(G51), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n524), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(new_n522), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT7), .Z(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT70), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n523), .A2(new_n524), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n524), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n543), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n532), .ZN(new_n555));
  AOI211_X1 g130(.A(new_n553), .B(new_n555), .C1(G43), .C2(new_n517), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT72), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n517), .A2(G53), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT9), .Z(new_n566));
  AOI22_X1  g141(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n567), .A2(new_n532), .B1(new_n544), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n566), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n530), .A2(new_n533), .ZN(G303));
  OAI21_X1  g147(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n517), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n523), .A2(new_n524), .A3(G87), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n523), .A2(KEYINPUT73), .A3(G61), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n522), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n544), .A2(new_n584), .B1(new_n546), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  XOR2_X1   g163(.A(KEYINPUT74), .B(G85), .Z(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n544), .A2(new_n589), .B1(new_n546), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n532), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G290));
  NAND3_X1  g172(.A1(new_n523), .A2(new_n524), .A3(G92), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n517), .A2(G54), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n532), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n566), .A2(new_n569), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  INV_X1    g186(.A(new_n603), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n492), .A2(G123), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n497), .A2(G135), .ZN(new_n620));
  OR2_X1    g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT76), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n503), .A2(new_n462), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2451), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT78), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2430), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n638), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n650), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n654), .B(new_n657), .Z(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT22), .B(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G32), .ZN(new_n679));
  NAND3_X1  g254(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT26), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n492), .B2(G129), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n497), .A2(G141), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n462), .A2(G105), .A3(new_n473), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(KEYINPUT87), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n682), .A2(new_n687), .A3(new_n683), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n686), .A2(KEYINPUT88), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n679), .B1(new_n693), .B2(new_n678), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT27), .B(G1996), .Z(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G6), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n586), .B1(G651), .B2(new_n582), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT80), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n697), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n697), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT34), .B1(new_n706), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n710), .A2(new_n715), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n718), .A2(new_n719), .A3(new_n704), .A4(new_n705), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n721));
  AOI22_X1  g296(.A1(G119), .A2(new_n492), .B1(new_n497), .B2(G131), .ZN(new_n722));
  OR2_X1    g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G25), .B(new_n725), .S(G29), .Z(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT35), .B(G1991), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n717), .A2(new_n720), .A3(new_n721), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n697), .A2(G24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n596), .B2(new_n697), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT79), .B(G1986), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  OR3_X1    g309(.A1(new_n730), .A2(KEYINPUT36), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT36), .B1(new_n730), .B2(new_n734), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n696), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  NAND2_X1  g313(.A1(G171), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G5), .B2(G16), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n694), .A2(new_n695), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G34), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G160), .B2(G29), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G2084), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT89), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n741), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT90), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n752));
  INV_X1    g327(.A(G20), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G16), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n754), .C1(new_n609), .C2(new_n697), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT92), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1956), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n678), .A2(G35), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n501), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT29), .ZN(new_n760));
  INV_X1    g335(.A(G2090), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n697), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n697), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n737), .A2(new_n750), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n740), .A2(new_n738), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n678), .A2(G26), .ZN(new_n773));
  AOI22_X1  g348(.A1(G128), .A2(new_n492), .B1(new_n497), .B2(G140), .ZN(new_n774));
  OR2_X1    g349(.A1(G104), .A2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n775), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n772), .B(new_n773), .C1(new_n777), .C2(G29), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n772), .B2(new_n773), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT84), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT83), .B(G2067), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n697), .A2(G4), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n612), .B2(new_n697), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1348), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n760), .A2(new_n761), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT91), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n678), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n678), .ZN(new_n789));
  INV_X1    g364(.A(G2078), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n745), .A2(G2084), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT31), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT30), .B(G28), .Z(new_n794));
  OAI221_X1 g369(.A(new_n792), .B1(new_n793), .B2(G11), .C1(G29), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n762), .B2(new_n763), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n787), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n793), .A2(G11), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n678), .A2(G33), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT25), .Z(new_n801));
  INV_X1    g376(.A(G139), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n496), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT85), .Z(new_n804));
  INV_X1    g379(.A(G127), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n480), .B2(new_n481), .ZN(new_n806));
  AND2_X1   g381(.A1(G115), .A2(G2104), .ZN(new_n807));
  OAI21_X1  g382(.A(G2105), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n799), .B1(new_n810), .B2(new_n678), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(G2072), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n697), .A2(G19), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n556), .B2(new_n697), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT82), .B(G1341), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n623), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(G29), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n797), .A2(new_n798), .A3(new_n812), .A4(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n771), .A2(new_n782), .A3(new_n785), .A4(new_n820), .ZN(G150));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n822));
  NAND2_X1  g397(.A1(G150), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n769), .A2(new_n819), .A3(new_n770), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n824), .A2(KEYINPUT94), .A3(new_n782), .A4(new_n785), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(G311));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n522), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT95), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n532), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n544), .A2(new_n832), .B1(new_n546), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n612), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT39), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n556), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n831), .A2(new_n834), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(KEYINPUT96), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n844), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n840), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n837), .B1(new_n848), .B2(G860), .ZN(G145));
  NAND3_X1  g424(.A1(new_n691), .A2(new_n810), .A3(new_n692), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n809), .A2(new_n686), .A3(new_n688), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n627), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n722), .A2(new_n854), .A3(new_n724), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n854), .B1(new_n722), .B2(new_n724), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n857), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n855), .A3(new_n627), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n862));
  INV_X1    g437(.A(G106), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n473), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n492), .B2(G130), .ZN(new_n865));
  INV_X1    g440(.A(G142), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n496), .A2(KEYINPUT97), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT97), .B1(new_n496), .B2(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(G164), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(G164), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n871), .A2(new_n774), .A3(new_n776), .A4(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n777), .B1(new_n874), .B2(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n861), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n861), .B1(new_n875), .B2(new_n873), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n852), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n873), .A2(new_n875), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n858), .A2(new_n860), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n883), .A2(new_n851), .A3(new_n876), .A4(new_n850), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n817), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n879), .A2(new_n884), .A3(new_n880), .A4(new_n623), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n501), .B(new_n486), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(new_n889), .A3(new_n887), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n891), .A2(KEYINPUT100), .A3(new_n892), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT40), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(G395));
  NAND2_X1  g477(.A1(new_n835), .A2(new_n604), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n847), .B(new_n615), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n612), .B(new_n609), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT101), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  MUX2_X1   g483(.A(KEYINPUT101), .B(new_n906), .S(new_n908), .Z(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT42), .ZN(new_n910));
  XNOR2_X1  g485(.A(G303), .B(new_n712), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(G305), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(new_n596), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n910), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n903), .B1(new_n914), .B2(new_n604), .ZN(G295));
  OAI21_X1  g490(.A(new_n903), .B1(new_n914), .B2(new_n604), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  INV_X1    g492(.A(new_n913), .ZN(new_n918));
  XNOR2_X1  g493(.A(G301), .B(G168), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n847), .B(new_n919), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n905), .A2(KEYINPUT103), .A3(KEYINPUT41), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n907), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT104), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n920), .A2(new_n926), .A3(new_n921), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n845), .A2(new_n846), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(new_n919), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n847), .A2(KEYINPUT102), .A3(new_n919), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n905), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n918), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n920), .A2(new_n905), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n907), .A3(new_n933), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(new_n913), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n892), .A4(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n892), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n913), .B1(new_n936), .B2(new_n937), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT44), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n935), .A2(new_n940), .A3(new_n892), .A4(new_n938), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n941), .B2(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n917), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n939), .B2(new_n943), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n946), .B2(new_n947), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT105), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n951), .A2(new_n954), .ZN(G397));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G164), .B2(G1384), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n505), .A2(new_n506), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G2105), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n509), .A2(new_n510), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n473), .ZN(new_n962));
  INV_X1    g537(.A(new_n481), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT64), .B1(new_n476), .B2(new_n477), .ZN(new_n964));
  OAI211_X1 g539(.A(G138), .B(new_n473), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT4), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(KEYINPUT106), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n957), .A2(new_n958), .A3(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n474), .B(G40), .C1(new_n485), .C2(new_n473), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n507), .A2(new_n511), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n973), .B2(new_n967), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n972), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n790), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n971), .A2(KEYINPUT121), .A3(new_n790), .A4(new_n975), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(KEYINPUT53), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n968), .A2(new_n969), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n958), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n975), .A2(new_n790), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT50), .B1(new_n957), .B2(new_n970), .ZN(new_n986));
  INV_X1    g561(.A(new_n972), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n974), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n738), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n980), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G171), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT122), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n968), .A2(KEYINPUT106), .A3(new_n969), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT106), .B1(new_n968), .B2(new_n969), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n988), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n972), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(KEYINPUT122), .A3(new_n738), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n482), .A2(KEYINPUT123), .A3(new_n484), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT123), .B1(new_n482), .B2(new_n484), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(G2105), .A3(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1005), .A2(G40), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(new_n982), .A3(new_n474), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT124), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT124), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1006), .A2(new_n982), .A3(new_n1009), .A4(new_n474), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n984), .B(G2078), .C1(new_n974), .C2(KEYINPUT45), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1002), .A2(G301), .A3(new_n985), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n993), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n986), .A2(new_n989), .ZN(new_n1016));
  INV_X1    g591(.A(G2084), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n971), .A2(new_n975), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n767), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(G168), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G168), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  OAI211_X1 g598(.A(G8), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT51), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1014), .A2(new_n1015), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT122), .B1(new_n1000), .B2(new_n738), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n994), .B(G1961), .C1(new_n998), .C2(new_n999), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n985), .B(new_n1012), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G171), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT125), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n980), .A2(new_n991), .A3(G301), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1034), .A2(KEYINPUT54), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1030), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(G166), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(G303), .A2(KEYINPUT107), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n975), .A2(new_n982), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(G1971), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n987), .B1(new_n996), .B2(new_n997), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n987), .A2(new_n988), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT113), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n957), .A2(new_n970), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(new_n987), .C1(new_n1053), .C2(new_n988), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n974), .A2(new_n988), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1051), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1057), .A2(new_n761), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1051), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT114), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1048), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1046), .B1(new_n1061), .B2(new_n1042), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1000), .A2(G2090), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1063), .B2(new_n1048), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1045), .B(KEYINPUT108), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1042), .B1(new_n1053), .B2(new_n987), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(G288), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT52), .ZN(new_n1070));
  INV_X1    g645(.A(G1981), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n699), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(G305), .B2(G1981), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n699), .A2(KEYINPUT109), .A3(new_n1071), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n1077));
  OR3_X1    g652(.A1(new_n1076), .A2(new_n1077), .A3(KEYINPUT49), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1076), .B2(KEYINPUT49), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(KEYINPUT49), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1067), .A4(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1067), .B(new_n1082), .C1(new_n1068), .C2(G288), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1070), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1066), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1027), .A2(new_n1037), .A3(new_n1062), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g663(.A(KEYINPUT118), .B1(G2067), .B2(new_n1049), .C1(new_n1016), .C2(G1348), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1348), .B1(new_n998), .B2(new_n999), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1049), .A2(G2067), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n603), .B1(new_n1094), .B2(KEYINPUT60), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1096), .B(new_n612), .C1(new_n1089), .C2(new_n1093), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1095), .A2(new_n1097), .B1(KEYINPUT60), .B2(new_n1094), .ZN(new_n1098));
  INV_X1    g673(.A(G1996), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1047), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1049), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT119), .B(G1341), .Z(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT58), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n556), .ZN(new_n1105));
  OR2_X1    g680(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1059), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n1114));
  OAI21_X1  g689(.A(G299), .B1(KEYINPUT117), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1047), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1117), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1111), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1122), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(KEYINPUT61), .A3(new_n1120), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1098), .A2(new_n1110), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1121), .A2(new_n603), .A3(new_n1094), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(new_n1122), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1066), .A2(new_n1084), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1060), .A2(new_n761), .A3(new_n1057), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1048), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1042), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1134), .B2(new_n1046), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(KEYINPUT126), .A3(new_n1027), .A4(new_n1037), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1088), .A2(new_n1129), .A3(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(new_n1042), .B(G286), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1085), .B(new_n1138), .C1(new_n1133), .C2(new_n1045), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT115), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1062), .A2(KEYINPUT115), .A3(new_n1085), .A4(new_n1138), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1084), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1064), .A2(new_n1046), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1070), .A2(new_n1081), .A3(KEYINPUT111), .A4(new_n1083), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1150), .A2(KEYINPUT63), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1066), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT116), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1138), .A4(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1144), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1146), .A2(new_n1066), .A3(new_n1149), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n712), .A2(new_n1068), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT112), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1081), .A2(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1067), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1026), .A2(new_n1024), .A3(new_n1164), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1085), .C1(new_n1133), .C2(new_n1045), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1026), .B2(new_n1024), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n993), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1137), .A2(new_n1156), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n982), .A2(new_n972), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n777), .B(G2067), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1099), .B1(new_n686), .B2(new_n688), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1173), .B(new_n1174), .C1(new_n693), .C2(new_n1099), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n725), .B(new_n728), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G1986), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n596), .B(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1172), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1171), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1172), .B1(new_n1173), .B2(new_n689), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1172), .A2(new_n1099), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT46), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT47), .Z(new_n1186));
  NAND3_X1  g761(.A1(new_n1172), .A2(new_n1178), .A3(new_n596), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT48), .Z(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n1177), .B2(new_n1172), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1175), .A2(new_n728), .A3(new_n722), .A4(new_n724), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(G2067), .B2(new_n777), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1186), .B(new_n1189), .C1(new_n1172), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1181), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1181), .A2(KEYINPUT127), .A3(new_n1192), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1195), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g772(.A(new_n460), .B(G229), .C1(new_n946), .C2(new_n947), .ZN(new_n1199));
  INV_X1    g773(.A(G227), .ZN(new_n1200));
  NAND4_X1  g774(.A1(new_n898), .A2(new_n1199), .A3(new_n645), .A4(new_n1200), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


