//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n566,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT70), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  OR2_X1    g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n466), .A2(KEYINPUT71), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  INV_X1    g059(.A(G137), .ZN(new_n485));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT71), .B(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n486), .B(new_n471), .C1(new_n487), .C2(new_n468), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n484), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n478), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G160));
  INV_X1    g067(.A(new_n488), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT72), .Z(new_n495));
  OAI21_X1  g070(.A(KEYINPUT73), .B1(G100), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g072(.A1(KEYINPUT73), .A2(G100), .A3(G2105), .ZN(new_n498));
  OAI221_X1 g073(.A(G2104), .B1(G112), .B2(new_n486), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G2105), .B(new_n471), .C1(new_n487), .C2(new_n468), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G124), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n495), .A2(new_n499), .A3(new_n502), .ZN(G162));
  NAND2_X1  g078(.A1(new_n470), .A2(new_n474), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G138), .A4(new_n486), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT4), .B1(new_n488), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G126), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT74), .B1(new_n500), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n467), .B1(new_n482), .B2(KEYINPUT3), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G126), .A4(G2105), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(G102), .A2(G2105), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n516), .B(G2104), .C1(G114), .C2(new_n486), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n509), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G50), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n527), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(G89), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n528), .A2(G543), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(G51), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT75), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  AOI22_X1  g123(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n526), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n529), .A2(new_n551), .B1(new_n531), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  AOI22_X1  g132(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n526), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  INV_X1    g135(.A(G43), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n529), .A2(new_n560), .B1(new_n531), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT78), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  NAND2_X1  g145(.A1(new_n543), .A2(G53), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT9), .Z(new_n572));
  AOI22_X1  g147(.A1(new_n524), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n573), .A2(new_n526), .B1(new_n529), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n572), .A2(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n543), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n529), .ZN(G288));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n521), .A2(new_n523), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n529), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n543), .A2(G48), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n584), .A2(KEYINPUT79), .A3(G651), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n587), .A2(new_n589), .A3(new_n590), .A4(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n543), .A2(G47), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT80), .B(G85), .Z(new_n594));
  AOI22_X1  g169(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n529), .B2(new_n594), .C1(new_n595), .C2(new_n526), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT82), .Z(new_n599));
  AND3_X1   g174(.A1(new_n521), .A2(new_n523), .A3(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n531), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT83), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n588), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n597), .B1(new_n608), .B2(G868), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n572), .A2(new_n575), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(G868), .B2(new_n612), .ZN(G297));
  OAI21_X1  g188(.A(new_n611), .B1(G868), .B2(new_n612), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n608), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n501), .A2(G123), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n493), .A2(G135), .ZN(new_n622));
  NOR2_X1   g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n486), .A2(KEYINPUT85), .A3(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT85), .B1(new_n486), .B2(G111), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(G2104), .A3(new_n625), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n504), .A2(new_n483), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT84), .B(G2100), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2435), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2438), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n640), .B(new_n645), .Z(new_n646));
  AND2_X1   g221(.A1(new_n646), .A2(G14), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT87), .Z(new_n654));
  XOR2_X1   g229(.A(new_n652), .B(KEYINPUT17), .Z(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n650), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n652), .A3(new_n648), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n650), .A3(new_n648), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2096), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2100), .Z(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n665), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  AOI22_X1  g246(.A1(new_n669), .A2(KEYINPUT20), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n665), .A3(new_n668), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n674), .C1(KEYINPUT20), .C2(new_n669), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G229));
  MUX2_X1   g257(.A(G24), .B(G290), .S(G16), .Z(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(G1986), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(G1986), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n686));
  INV_X1    g261(.A(G119), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n500), .B2(new_n687), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n512), .A2(KEYINPUT89), .A3(G119), .A4(G2105), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(G95), .A2(G2105), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n691), .B(G2104), .C1(G107), .C2(new_n486), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n493), .A2(G131), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n690), .A2(new_n696), .A3(new_n692), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G25), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT91), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n684), .B(new_n685), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G22), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT92), .B1(G16), .B2(G23), .ZN(new_n712));
  OR3_X1    g287(.A1(KEYINPUT92), .A2(G16), .A3(G23), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n712), .B(new_n713), .C1(G288), .C2(new_n707), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n707), .A2(G6), .ZN(new_n717));
  INV_X1    g292(.A(G305), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n707), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT32), .B(G1981), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n711), .A2(new_n716), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT34), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n706), .B(new_n724), .C1(new_n705), .C2(new_n702), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT36), .Z(new_n726));
  AND2_X1   g301(.A1(new_n700), .A2(G26), .ZN(new_n727));
  OR2_X1    g302(.A1(G104), .A2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT94), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n466), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n730), .B1(new_n729), .B2(new_n728), .C1(G116), .C2(new_n486), .ZN(new_n731));
  INV_X1    g306(.A(G128), .ZN(new_n732));
  INV_X1    g307(.A(G140), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n731), .B1(new_n732), .B2(new_n500), .C1(new_n733), .C2(new_n488), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(G29), .ZN(new_n735));
  MUX2_X1   g310(.A(new_n727), .B(new_n735), .S(KEYINPUT28), .Z(new_n736));
  XOR2_X1   g311(.A(KEYINPUT95), .B(G2067), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n700), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n700), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2090), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n743), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n707), .A2(G20), .ZN(new_n746));
  NAND2_X1  g321(.A1(G299), .A2(G16), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(KEYINPUT23), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(KEYINPUT23), .B2(new_n746), .ZN(new_n749));
  INV_X1    g324(.A(G1956), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n744), .B(new_n745), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n608), .A2(new_n707), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G4), .B2(new_n707), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT93), .B(G1348), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G5), .B2(G16), .ZN(new_n758));
  OR3_X1    g333(.A1(new_n757), .A2(G5), .A3(G16), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n758), .B(new_n759), .C1(G301), .C2(new_n707), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n749), .B2(new_n750), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n707), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n707), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1966), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n700), .B1(new_n767), .B2(G28), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(G28), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n563), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G16), .B2(G19), .ZN(new_n771));
  INV_X1    g346(.A(G1341), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  NOR2_X1   g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n774), .A2(new_n775), .A3(G29), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n491), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n773), .B1(new_n772), .B2(new_n771), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n755), .A2(new_n756), .A3(new_n763), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n627), .A2(new_n700), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT97), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n778), .B2(new_n777), .ZN(new_n784));
  NAND2_X1  g359(.A1(G164), .A2(G29), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G27), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(G2078), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G29), .A2(G32), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n493), .A2(G141), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n501), .A2(G129), .ZN(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT26), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n483), .A2(G105), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n790), .A2(new_n791), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n789), .B1(new_n796), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT27), .B(G1996), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n786), .A2(new_n787), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n784), .A2(new_n788), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n504), .A2(G127), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n803));
  NAND2_X1  g378(.A1(G115), .A2(G2104), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G127), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n470), .B2(new_n474), .ZN(new_n807));
  INV_X1    g382(.A(new_n804), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT96), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n805), .A2(new_n809), .A3(G2105), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n493), .A2(G139), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n486), .A2(G103), .A3(G2104), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT25), .Z(new_n813));
  NAND3_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G33), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(G2072), .Z(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n753), .B2(new_n754), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n781), .A2(new_n801), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n726), .A2(new_n738), .A3(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n529), .A2(new_n821), .B1(new_n531), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(KEYINPUT100), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OAI22_X1  g401(.A1(new_n824), .A2(new_n825), .B1(new_n526), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G860), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n607), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n615), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n827), .A2(KEYINPUT101), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n559), .B2(new_n562), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n827), .A2(KEYINPUT101), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n833), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n829), .B1(new_n840), .B2(G860), .ZN(G145));
  NAND2_X1  g416(.A1(new_n501), .A2(G130), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n493), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(G106), .A2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(new_n486), .B2(G118), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n630), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n734), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n814), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n810), .A2(new_n734), .A3(new_n811), .A4(new_n813), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n698), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n698), .B1(new_n850), .B2(new_n851), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n518), .B(new_n795), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n850), .A2(new_n851), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n699), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n855), .B1(new_n859), .B2(new_n852), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n848), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n856), .B1(new_n853), .B2(new_n854), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n859), .A2(new_n855), .A3(new_n852), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n847), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n491), .B(new_n627), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n861), .A2(new_n865), .A3(new_n862), .A4(new_n867), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n872));
  XOR2_X1   g447(.A(G162), .B(new_n872), .Z(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT104), .B(G37), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n873), .A3(new_n870), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT106), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n875), .A2(new_n880), .A3(new_n876), .A4(new_n877), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n879), .A2(KEYINPUT40), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT40), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(G395));
  XNOR2_X1  g459(.A(new_n839), .B(new_n617), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n608), .A2(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n830), .A2(new_n612), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(KEYINPUT41), .A3(new_n887), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n890), .A2(KEYINPUT107), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n889), .B1(new_n885), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(G303), .B(G288), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G290), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n899), .A2(G305), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(G305), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(KEYINPUT42), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n897), .B(new_n903), .ZN(new_n904));
  MUX2_X1   g479(.A(new_n827), .B(new_n904), .S(G868), .Z(G295));
  MUX2_X1   g480(.A(new_n827), .B(new_n904), .S(G868), .Z(G331));
  XNOR2_X1  g481(.A(G286), .B(G301), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n839), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n837), .A2(new_n838), .A3(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n888), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(new_n902), .C1(new_n896), .C2(new_n911), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n909), .A2(new_n910), .B1(new_n887), .B2(new_n886), .ZN(new_n915));
  INV_X1    g490(.A(new_n896), .ZN(new_n916));
  INV_X1    g491(.A(new_n911), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n902), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n900), .A2(KEYINPUT108), .A3(new_n901), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n913), .B(new_n914), .C1(new_n918), .C2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n894), .A2(new_n909), .A3(new_n910), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n922), .B1(new_n926), .B2(new_n915), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n876), .A3(new_n913), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n925), .A2(new_n931), .A3(KEYINPUT44), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n927), .A2(new_n913), .A3(new_n935), .A4(new_n876), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(KEYINPUT44), .B2(new_n937), .ZN(G397));
  INV_X1    g513(.A(KEYINPUT60), .ZN(new_n939));
  INV_X1    g514(.A(G40), .ZN(new_n940));
  AOI211_X1 g515(.A(new_n940), .B(new_n489), .C1(new_n477), .C2(G2105), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n508), .A2(new_n506), .B1(new_n511), .B2(new_n514), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n942), .B2(new_n517), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n518), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT119), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n478), .A2(new_n490), .A3(G40), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n518), .A2(new_n946), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(KEYINPUT50), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT119), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n947), .ZN(new_n954));
  AOI21_X1  g529(.A(G1348), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n943), .A2(new_n941), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(G2067), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n608), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1348), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n944), .B1(new_n518), .B2(new_n946), .ZN(new_n960));
  NOR4_X1   g535(.A1(new_n948), .A2(new_n960), .A3(KEYINPUT119), .A4(new_n950), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n953), .B1(new_n952), .B2(new_n947), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n957), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n830), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n939), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n951), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n518), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT120), .B(G1996), .Z(new_n970));
  NAND4_X1  g545(.A1(new_n968), .A2(new_n941), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT58), .B(G1341), .Z(new_n972));
  NAND2_X1  g547(.A1(new_n956), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n563), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT59), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT59), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n977), .A3(new_n563), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n963), .A2(new_n939), .A3(new_n608), .A4(new_n964), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n966), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT61), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT115), .B1(new_n943), .B2(new_n944), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n947), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n952), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT116), .B(G1956), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(G299), .A2(KEYINPUT117), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n572), .A2(KEYINPUT117), .A3(new_n575), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(KEYINPUT57), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n612), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n996), .B2(new_n991), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT56), .B(G2072), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n968), .A2(new_n941), .A3(new_n999), .A4(new_n969), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n518), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT45), .B1(new_n518), .B2(new_n946), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1005), .A2(KEYINPUT118), .A3(new_n941), .A4(new_n999), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n989), .A2(new_n998), .A3(new_n1002), .A4(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT122), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n983), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n993), .A2(new_n997), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1002), .ZN(new_n1011));
  INV_X1    g586(.A(new_n988), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n947), .B(new_n985), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(new_n952), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1010), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(KEYINPUT122), .A3(new_n998), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1009), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1007), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n983), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT121), .B(KEYINPUT61), .C1(new_n1015), .C2(new_n1007), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n982), .B(new_n1018), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1015), .A2(new_n958), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1007), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1961), .B1(new_n949), .B2(new_n954), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1003), .A2(new_n1004), .A3(new_n950), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n1028), .B2(new_n787), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n968), .A2(new_n941), .A3(new_n969), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(G2078), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1027), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G301), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n486), .B1(new_n477), .B2(KEYINPUT123), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n475), .A2(KEYINPUT123), .A3(new_n476), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n940), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(new_n490), .C1(KEYINPUT45), .C2(new_n943), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT124), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1031), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n968), .A2(KEYINPUT124), .A3(new_n490), .A4(new_n1037), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n787), .A3(new_n969), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1029), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n761), .B1(new_n961), .B2(new_n962), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1034), .B(KEYINPUT54), .C1(G301), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n587), .A2(new_n1047), .A3(new_n591), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G1981), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n718), .ZN(new_n1050));
  NAND3_X1  g625(.A1(G305), .A2(G1981), .A3(new_n1048), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT49), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n951), .A2(new_n950), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1050), .A2(KEYINPUT49), .A3(new_n1051), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(KEYINPUT114), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1054), .A2(new_n1053), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT112), .B1(G288), .B2(new_n1061), .ZN(new_n1062));
  OR3_X1    g637(.A1(G288), .A2(KEYINPUT112), .A3(new_n1061), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .A4(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1059), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n951), .A2(KEYINPUT50), .ZN(new_n1069));
  INV_X1    g644(.A(G2090), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n941), .A4(new_n947), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1030), .A2(new_n710), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n952), .A2(KEYINPUT110), .A3(new_n1070), .A4(new_n947), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G303), .A2(G8), .ZN(new_n1077));
  XOR2_X1   g652(.A(new_n1077), .B(KEYINPUT55), .Z(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(G8), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT111), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1076), .A2(new_n1081), .A3(G8), .A4(new_n1078), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1068), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1074), .B1(new_n987), .B2(G2090), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n1084), .B2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1046), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1042), .A2(G301), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1033), .B2(G301), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G286), .A2(G8), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n948), .A2(new_n960), .A3(new_n950), .ZN(new_n1094));
  INV_X1    g669(.A(G1966), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1094), .A2(new_n778), .B1(new_n1030), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1092), .B(new_n1093), .C1(new_n1096), .C2(new_n1053), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n952), .A2(new_n778), .A3(new_n947), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1028), .B2(G1966), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT51), .B(G8), .C1(new_n1099), .C2(G286), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(G8), .A3(G286), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1091), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1087), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1026), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G288), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G305), .A2(G1981), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1060), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1068), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1080), .A2(new_n1111), .A3(new_n1082), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1101), .A2(new_n1114), .A3(new_n1102), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1033), .A2(G301), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1083), .A2(new_n1115), .A3(new_n1116), .A4(new_n1086), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1085), .B(new_n1068), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(KEYINPUT125), .A3(new_n1116), .A4(new_n1115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1096), .A2(new_n1053), .A3(G286), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1078), .B1(new_n1076), .B2(G8), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n1124), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1083), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1106), .A2(new_n1113), .A3(new_n1123), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n968), .A2(new_n950), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n734), .B(G2067), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n795), .A2(G1996), .ZN(new_n1136));
  INV_X1    g711(.A(G1996), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n796), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n699), .A2(new_n705), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n698), .A2(new_n704), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G290), .B(G1986), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1134), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1133), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1134), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1135), .B2(new_n796), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1134), .A2(KEYINPUT46), .A3(new_n1137), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT46), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT47), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1139), .A2(new_n1141), .B1(G2067), .B2(new_n734), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1134), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT126), .Z(new_n1155));
  NOR3_X1   g730(.A1(new_n1147), .A2(G1986), .A3(G290), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT127), .ZN(new_n1157));
  XOR2_X1   g732(.A(new_n1157), .B(KEYINPUT48), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1143), .A2(new_n1134), .ZN(new_n1159));
  AOI211_X1 g734(.A(new_n1152), .B(new_n1155), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1146), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g736(.A(G319), .ZN(new_n1163));
  NOR2_X1   g737(.A1(G229), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g738(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g739(.A(new_n1165), .B1(new_n934), .B2(new_n936), .ZN(new_n1166));
  NOR2_X1   g740(.A1(G227), .A2(G401), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n1166), .A2(new_n878), .A3(new_n1167), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


