

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X2 U320 ( .A(n403), .B(KEYINPUT113), .ZN(n404) );
  XOR2_X2 U321 ( .A(G99GAT), .B(G85GAT), .Z(n361) );
  XNOR2_X1 U322 ( .A(n380), .B(n379), .ZN(n381) );
  INV_X1 U323 ( .A(KEYINPUT45), .ZN(n379) );
  NOR2_X1 U324 ( .A1(n577), .A2(n400), .ZN(n401) );
  XNOR2_X1 U325 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n407) );
  INV_X1 U327 ( .A(KEYINPUT124), .ZN(n449) );
  OR2_X2 U328 ( .A1(n448), .A2(n529), .ZN(n450) );
  AND2_X1 U329 ( .A1(G230GAT), .A2(G233GAT), .ZN(n288) );
  AND2_X1 U330 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U331 ( .A(n418), .B(n391), .Z(n290) );
  XNOR2_X1 U332 ( .A(n361), .B(n289), .ZN(n363) );
  XNOR2_X1 U333 ( .A(n363), .B(n362), .ZN(n366) );
  INV_X1 U334 ( .A(KEYINPUT75), .ZN(n351) );
  XNOR2_X1 U335 ( .A(n295), .B(n288), .ZN(n296) );
  XNOR2_X1 U336 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n301) );
  XNOR2_X1 U338 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U339 ( .A(n374), .B(n373), .Z(n377) );
  XNOR2_X1 U340 ( .A(n305), .B(n304), .ZN(n574) );
  XOR2_X1 U341 ( .A(n358), .B(n357), .Z(n555) );
  XNOR2_X1 U342 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U343 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n292) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U345 ( .A(n439), .B(n361), .ZN(n291) );
  XNOR2_X1 U346 ( .A(n292), .B(n291), .ZN(n297) );
  XOR2_X1 U347 ( .A(KEYINPUT32), .B(KEYINPUT70), .Z(n294) );
  XNOR2_X1 U348 ( .A(KEYINPUT71), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U350 ( .A(KEYINPUT72), .B(G64GAT), .Z(n299) );
  XNOR2_X1 U351 ( .A(G204GAT), .B(G92GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U353 ( .A(G176GAT), .B(n300), .Z(n329) );
  XNOR2_X1 U354 ( .A(n301), .B(n329), .ZN(n305) );
  XNOR2_X1 U355 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n302), .B(G148GAT), .ZN(n426) );
  XNOR2_X1 U357 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n303), .B(KEYINPUT13), .ZN(n350) );
  XOR2_X1 U359 ( .A(n426), .B(n350), .Z(n304) );
  XNOR2_X1 U360 ( .A(KEYINPUT41), .B(n574), .ZN(n550) );
  INV_X1 U361 ( .A(n550), .ZN(n534) );
  XOR2_X1 U362 ( .A(G134GAT), .B(KEYINPUT74), .Z(n375) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n306), .B(G127GAT), .ZN(n438) );
  XOR2_X1 U365 ( .A(n375), .B(n438), .Z(n308) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U368 ( .A(n309), .B(KEYINPUT1), .Z(n312) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n310), .B(KEYINPUT2), .ZN(n425) );
  XNOR2_X1 U371 ( .A(n425), .B(KEYINPUT88), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U373 ( .A(G85GAT), .B(G162GAT), .Z(n314) );
  XNOR2_X1 U374 ( .A(G29GAT), .B(G148GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U376 ( .A(n316), .B(n315), .Z(n324) );
  XOR2_X1 U377 ( .A(KEYINPUT4), .B(KEYINPUT87), .Z(n318) );
  XNOR2_X1 U378 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U380 ( .A(G57GAT), .B(G155GAT), .Z(n320) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(G120GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n515) );
  XNOR2_X1 U385 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n325), .B(KEYINPUT18), .ZN(n326) );
  XOR2_X1 U387 ( .A(n326), .B(KEYINPUT83), .Z(n328) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(G183GAT), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n443) );
  XNOR2_X1 U390 ( .A(n443), .B(n329), .ZN(n339) );
  XNOR2_X1 U391 ( .A(G36GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n330), .B(G218GAT), .ZN(n362) );
  XOR2_X1 U393 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n332) );
  NAND2_X1 U394 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U396 ( .A(n362), .B(n333), .Z(n337) );
  XOR2_X1 U397 ( .A(G211GAT), .B(KEYINPUT21), .Z(n335) );
  XNOR2_X1 U398 ( .A(G197GAT), .B(KEYINPUT86), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n414) );
  XNOR2_X1 U400 ( .A(G8GAT), .B(n414), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n517) );
  XOR2_X1 U403 ( .A(G64GAT), .B(KEYINPUT79), .Z(n341) );
  XNOR2_X1 U404 ( .A(KEYINPUT76), .B(KEYINPUT78), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n358) );
  XOR2_X1 U406 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n343) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(KEYINPUT14), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U409 ( .A(G211GAT), .B(G78GAT), .Z(n345) );
  XNOR2_X1 U410 ( .A(G127GAT), .B(G71GAT), .ZN(n344) );
  XNOR2_X1 U411 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n356) );
  XOR2_X1 U413 ( .A(G22GAT), .B(G155GAT), .Z(n418) );
  XNOR2_X1 U414 ( .A(G15GAT), .B(G1GAT), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n348), .B(G8GAT), .ZN(n391) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n290), .B(n349), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n350), .B(KEYINPUT15), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U420 ( .A(G92GAT), .B(KEYINPUT9), .Z(n360) );
  XNOR2_X1 U421 ( .A(G106GAT), .B(KEYINPUT10), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n374) );
  INV_X1 U423 ( .A(n366), .ZN(n364) );
  NAND2_X1 U424 ( .A1(n364), .A2(KEYINPUT11), .ZN(n368) );
  INV_X1 U425 ( .A(KEYINPUT11), .ZN(n365) );
  NAND2_X1 U426 ( .A1(n366), .A2(n365), .ZN(n367) );
  NAND2_X1 U427 ( .A1(n368), .A2(n367), .ZN(n372) );
  XOR2_X1 U428 ( .A(G29GAT), .B(G43GAT), .Z(n370) );
  XNOR2_X1 U429 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n392) );
  XNOR2_X1 U431 ( .A(n392), .B(KEYINPUT73), .ZN(n371) );
  XOR2_X1 U432 ( .A(G50GAT), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U433 ( .A(n413), .B(n375), .ZN(n376) );
  XOR2_X2 U434 ( .A(n377), .B(n376), .Z(n564) );
  INV_X1 U435 ( .A(KEYINPUT36), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n564), .B(n378), .ZN(n581) );
  NOR2_X1 U437 ( .A1(n555), .A2(n581), .ZN(n380) );
  NOR2_X1 U438 ( .A1(n574), .A2(n381), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT114), .ZN(n397) );
  XOR2_X1 U440 ( .A(G36GAT), .B(G50GAT), .Z(n384) );
  NAND2_X1 U441 ( .A1(G229GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n396) );
  XOR2_X1 U443 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n386) );
  XNOR2_X1 U444 ( .A(G169GAT), .B(KEYINPUT67), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U446 ( .A(G113GAT), .B(G22GAT), .Z(n388) );
  XNOR2_X1 U447 ( .A(G141GAT), .B(G197GAT), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U449 ( .A(n390), .B(n389), .Z(n394) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U452 ( .A(n396), .B(n395), .Z(n571) );
  INV_X1 U453 ( .A(n571), .ZN(n548) );
  NAND2_X1 U454 ( .A1(n397), .A2(n548), .ZN(n406) );
  INV_X1 U455 ( .A(n555), .ZN(n577) );
  NOR2_X1 U456 ( .A1(n550), .A2(n548), .ZN(n399) );
  XOR2_X1 U457 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U459 ( .A(KEYINPUT112), .B(n401), .ZN(n402) );
  INV_X1 U460 ( .A(n564), .ZN(n558) );
  NAND2_X1 U461 ( .A1(n402), .A2(n558), .ZN(n403) );
  XNOR2_X1 U462 ( .A(KEYINPUT47), .B(n404), .ZN(n405) );
  NAND2_X1 U463 ( .A1(n406), .A2(n405), .ZN(n408) );
  XNOR2_X2 U464 ( .A(n408), .B(n407), .ZN(n546) );
  AND2_X2 U465 ( .A1(n517), .A2(n546), .ZN(n410) );
  XNOR2_X1 U466 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  NOR2_X1 U468 ( .A1(n515), .A2(n411), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n412), .B(KEYINPUT65), .ZN(n569) );
  XOR2_X1 U470 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U473 ( .A(n417), .B(KEYINPUT23), .Z(n420) );
  XNOR2_X1 U474 ( .A(G218GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U476 ( .A(KEYINPUT85), .B(KEYINPUT22), .Z(n422) );
  XNOR2_X1 U477 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U479 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n466) );
  NOR2_X1 U482 ( .A1(n569), .A2(n466), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n429), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U484 ( .A(KEYINPUT80), .B(KEYINPUT84), .Z(n431) );
  XNOR2_X1 U485 ( .A(G15GAT), .B(KEYINPUT66), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n447) );
  XOR2_X1 U487 ( .A(G134GAT), .B(G99GAT), .Z(n433) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G190GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U490 ( .A(KEYINPUT81), .B(G176GAT), .Z(n435) );
  XNOR2_X1 U491 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n445) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n520) );
  INV_X1 U500 ( .A(n520), .ZN(n529) );
  XNOR2_X2 U501 ( .A(n450), .B(n449), .ZN(n563) );
  NAND2_X1 U502 ( .A1(n534), .A2(n563), .ZN(n454) );
  XOR2_X1 U503 ( .A(G176GAT), .B(KEYINPUT56), .Z(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n451) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(G1349GAT) );
  XOR2_X1 U506 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n474) );
  NOR2_X1 U507 ( .A1(n574), .A2(n548), .ZN(n486) );
  AND2_X1 U508 ( .A1(n520), .A2(n517), .ZN(n455) );
  NOR2_X1 U509 ( .A1(n466), .A2(n455), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(KEYINPUT25), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT93), .ZN(n462) );
  NAND2_X1 U512 ( .A1(n466), .A2(n529), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT26), .ZN(n570) );
  XNOR2_X1 U514 ( .A(n517), .B(KEYINPUT27), .ZN(n465) );
  INV_X1 U515 ( .A(n465), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n570), .A2(n459), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n460), .B(KEYINPUT92), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT94), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n515), .A2(n464), .ZN(n469) );
  NAND2_X1 U521 ( .A1(n515), .A2(n465), .ZN(n545) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT28), .ZN(n522) );
  NOR2_X1 U523 ( .A1(n545), .A2(n522), .ZN(n527) );
  XNOR2_X1 U524 ( .A(KEYINPUT91), .B(n527), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n520), .A2(n467), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n483) );
  NOR2_X1 U527 ( .A1(n555), .A2(n564), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  NOR2_X1 U529 ( .A1(n483), .A2(n471), .ZN(n502) );
  NAND2_X1 U530 ( .A1(n486), .A2(n502), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT95), .B(n472), .ZN(n481) );
  NAND2_X1 U532 ( .A1(n481), .A2(n515), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U534 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  NAND2_X1 U535 ( .A1(n481), .A2(n517), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n478) );
  NAND2_X1 U538 ( .A1(n481), .A2(n520), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n480) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT97), .Z(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U542 ( .A1(n522), .A2(n481), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U544 ( .A1(n483), .A2(n581), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n484), .A2(n555), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n485), .B(KEYINPUT37), .ZN(n514) );
  NAND2_X1 U547 ( .A1(n486), .A2(n514), .ZN(n487) );
  XOR2_X1 U548 ( .A(KEYINPUT38), .B(n487), .Z(n498) );
  NAND2_X1 U549 ( .A1(n498), .A2(n515), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n489) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT99), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n517), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(KEYINPUT102), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n496) );
  NAND2_X1 U559 ( .A1(n498), .A2(n520), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n498), .A2(n522), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  NAND2_X1 U565 ( .A1(n548), .A2(n534), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(KEYINPUT105), .ZN(n513) );
  AND2_X1 U567 ( .A1(n502), .A2(n513), .ZN(n509) );
  NAND2_X1 U568 ( .A1(n515), .A2(n509), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n517), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n507) );
  NAND2_X1 U574 ( .A1(n509), .A2(n520), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U578 ( .A1(n509), .A2(n522), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  AND2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n523), .A2(n515), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U584 ( .A(G92GAT), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U585 ( .A1(n523), .A2(n517), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n523), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n525) );
  NAND2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n532) );
  NAND2_X1 U594 ( .A1(n527), .A2(n546), .ZN(n528) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(n530), .Z(n541) );
  NAND2_X1 U597 ( .A1(n541), .A2(n571), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n536) );
  NAND2_X1 U601 ( .A1(n541), .A2(n534), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n539) );
  NAND2_X1 U605 ( .A1(n541), .A2(n577), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U609 ( .A1(n541), .A2(n564), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n570), .A2(n545), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n548), .A2(n557), .ZN(n549) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U616 ( .A1(n557), .A2(n550), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n552) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n557), .ZN(n556) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT122), .B(n559), .Z(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n571), .A2(n563), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n577), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT60), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(n568), .Z(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U640 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n579), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U644 ( .A(n579), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

