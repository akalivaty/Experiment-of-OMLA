

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761;

  NOR2_X1 U376 ( .A1(n680), .A2(n681), .ZN(n578) );
  XNOR2_X1 U377 ( .A(n617), .B(KEYINPUT38), .ZN(n678) );
  XNOR2_X1 U378 ( .A(G107), .B(G104), .ZN(n438) );
  INV_X1 U379 ( .A(G119), .ZN(n376) );
  XNOR2_X2 U380 ( .A(n388), .B(n571), .ZN(n617) );
  XNOR2_X1 U381 ( .A(n375), .B(n432), .ZN(n436) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n514) );
  INV_X1 U383 ( .A(G953), .ZN(n482) );
  XNOR2_X1 U384 ( .A(G137), .B(G119), .ZN(n487) );
  XNOR2_X1 U385 ( .A(G113), .B(G104), .ZN(n518) );
  OR2_X2 U386 ( .A1(n711), .A2(KEYINPUT2), .ZN(n353) );
  XNOR2_X2 U387 ( .A(n626), .B(n625), .ZN(n412) );
  NAND2_X2 U388 ( .A1(n379), .A2(n377), .ZN(n626) );
  XNOR2_X2 U389 ( .A(n555), .B(n469), .ZN(n552) );
  OR2_X1 U390 ( .A1(n394), .A2(n396), .ZN(n402) );
  XNOR2_X1 U391 ( .A(n391), .B(KEYINPUT107), .ZN(n390) );
  AND2_X1 U392 ( .A1(n421), .A2(n420), .ZN(n419) );
  NAND2_X1 U393 ( .A1(n760), .A2(n662), .ZN(n559) );
  XNOR2_X1 U394 ( .A(n530), .B(n431), .ZN(n541) );
  OR2_X1 U395 ( .A1(n545), .A2(n537), .ZN(n538) );
  XNOR2_X1 U396 ( .A(n406), .B(n405), .ZN(n669) );
  NOR2_X1 U397 ( .A1(n600), .A2(n452), .ZN(n453) );
  XNOR2_X1 U398 ( .A(n402), .B(n447), .ZN(n600) );
  OR2_X1 U399 ( .A1(n688), .A2(n687), .ZN(n501) );
  OR2_X1 U400 ( .A1(n640), .A2(G902), .ZN(n496) );
  XNOR2_X1 U401 ( .A(n414), .B(n413), .ZN(n640) );
  XNOR2_X1 U402 ( .A(n490), .B(n360), .ZN(n414) );
  XNOR2_X1 U403 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U404 ( .A(n436), .B(n435), .ZN(n475) );
  XNOR2_X1 U405 ( .A(n426), .B(n439), .ZN(n425) );
  XNOR2_X1 U406 ( .A(n510), .B(n458), .ZN(n473) );
  XNOR2_X1 U407 ( .A(n744), .B(n484), .ZN(n413) );
  XNOR2_X1 U408 ( .A(n455), .B(n454), .ZN(n510) );
  XNOR2_X1 U409 ( .A(n376), .B(G113), .ZN(n375) );
  INV_X2 U410 ( .A(G143), .ZN(n369) );
  XNOR2_X1 U411 ( .A(n697), .B(n410), .ZN(n589) );
  NOR2_X1 U412 ( .A1(n682), .A2(n557), .ZN(n558) );
  NOR2_X1 U413 ( .A1(n669), .A2(n355), .ZN(n557) );
  XNOR2_X1 U414 ( .A(n613), .B(n366), .ZN(n385) );
  INV_X1 U415 ( .A(G134), .ZN(n454) );
  INV_X1 U416 ( .A(KEYINPUT82), .ZN(n373) );
  NOR2_X1 U417 ( .A1(n675), .A2(KEYINPUT80), .ZN(n384) );
  NOR2_X1 U418 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U419 ( .A(n637), .ZN(n381) );
  NOR2_X1 U420 ( .A1(n619), .A2(n620), .ZN(n382) );
  NAND2_X1 U421 ( .A1(n368), .A2(n392), .ZN(n391) );
  XNOR2_X1 U422 ( .A(KEYINPUT24), .B(G128), .ZN(n486) );
  NAND2_X1 U423 ( .A1(n690), .A2(n589), .ZN(n409) );
  NAND2_X1 U424 ( .A1(n399), .A2(n397), .ZN(n396) );
  NOR2_X1 U425 ( .A1(n398), .A2(n403), .ZN(n397) );
  NAND2_X1 U426 ( .A1(n651), .A2(n400), .ZN(n399) );
  AND2_X1 U427 ( .A1(n571), .A2(n401), .ZN(n398) );
  XNOR2_X1 U428 ( .A(n453), .B(KEYINPUT0), .ZN(n533) );
  XNOR2_X1 U429 ( .A(n434), .B(n433), .ZN(n435) );
  INV_X1 U430 ( .A(KEYINPUT3), .ZN(n433) );
  XNOR2_X1 U431 ( .A(n483), .B(KEYINPUT8), .ZN(n508) );
  AND2_X1 U432 ( .A1(G234), .A2(n482), .ZN(n483) );
  XNOR2_X1 U433 ( .A(G116), .B(G107), .ZN(n504) );
  XOR2_X1 U434 ( .A(n459), .B(n473), .Z(n746) );
  XNOR2_X1 U435 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U436 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n440) );
  NAND2_X1 U437 ( .A1(n430), .A2(n362), .ZN(n429) );
  NOR2_X1 U438 ( .A1(n361), .A2(n371), .ZN(n370) );
  OR2_X1 U439 ( .A1(G902), .A2(G237), .ZN(n446) );
  NOR2_X1 U440 ( .A1(n571), .A2(n401), .ZN(n400) );
  INV_X1 U441 ( .A(n677), .ZN(n403) );
  XOR2_X1 U442 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n471) );
  AND2_X1 U443 ( .A1(n544), .A2(n364), .ZN(n420) );
  NAND2_X1 U444 ( .A1(G237), .A2(G234), .ZN(n448) );
  AND2_X1 U445 ( .A1(n621), .A2(n656), .ZN(n682) );
  NAND2_X1 U446 ( .A1(n378), .A2(KEYINPUT80), .ZN(n377) );
  AND2_X1 U447 ( .A1(n383), .A2(n380), .ZN(n379) );
  INV_X1 U448 ( .A(n571), .ZN(n395) );
  INV_X1 U449 ( .A(G902), .ZN(n525) );
  XNOR2_X1 U450 ( .A(KEYINPUT94), .B(KEYINPUT23), .ZN(n484) );
  XNOR2_X1 U451 ( .A(G110), .B(KEYINPUT93), .ZN(n485) );
  XOR2_X1 U452 ( .A(KEYINPUT98), .B(G131), .Z(n521) );
  XNOR2_X1 U453 ( .A(G143), .B(G122), .ZN(n520) );
  XOR2_X1 U454 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n516) );
  NOR2_X1 U455 ( .A1(n552), .A2(n409), .ZN(n408) );
  INV_X1 U456 ( .A(KEYINPUT6), .ZN(n410) );
  XNOR2_X1 U457 ( .A(n534), .B(KEYINPUT22), .ZN(n545) );
  XNOR2_X1 U458 ( .A(n550), .B(n404), .ZN(n554) );
  INV_X1 U459 ( .A(KEYINPUT89), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n374), .B(n509), .ZN(n726) );
  XNOR2_X1 U461 ( .A(n424), .B(n444), .ZN(n389) );
  XNOR2_X1 U462 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n405) );
  NAND2_X1 U463 ( .A1(n356), .A2(n553), .ZN(n406) );
  NOR2_X2 U464 ( .A1(n601), .A2(n600), .ZN(n665) );
  AND2_X1 U465 ( .A1(n549), .A2(n548), .ZN(n670) );
  XNOR2_X1 U466 ( .A(n546), .B(KEYINPUT106), .ZN(n757) );
  AND2_X1 U467 ( .A1(n428), .A2(n427), .ZN(n546) );
  XNOR2_X1 U468 ( .A(n429), .B(KEYINPUT81), .ZN(n428) );
  XNOR2_X1 U469 ( .A(n722), .B(n721), .ZN(n723) );
  XOR2_X1 U470 ( .A(n358), .B(n506), .Z(n354) );
  NOR2_X1 U471 ( .A1(n554), .A2(n359), .ZN(n355) );
  NOR2_X1 U472 ( .A1(n552), .A2(n551), .ZN(n356) );
  AND2_X1 U473 ( .A1(n713), .A2(n401), .ZN(n357) );
  XOR2_X1 U474 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n358) );
  OR2_X1 U475 ( .A1(n556), .A2(n697), .ZN(n359) );
  AND2_X2 U476 ( .A1(n357), .A2(n353), .ZN(n725) );
  AND2_X1 U477 ( .A1(n508), .A2(G221), .ZN(n360) );
  AND2_X1 U478 ( .A1(KEYINPUT78), .A2(n682), .ZN(n361) );
  NOR2_X1 U479 ( .A1(n691), .A2(n589), .ZN(n362) );
  AND2_X1 U480 ( .A1(G217), .A2(n508), .ZN(n363) );
  OR2_X1 U481 ( .A1(n559), .A2(KEYINPUT64), .ZN(n364) );
  XOR2_X1 U482 ( .A(n502), .B(KEYINPUT71), .Z(n365) );
  XNOR2_X1 U483 ( .A(n408), .B(n365), .ZN(n676) );
  XOR2_X1 U484 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n366) );
  INV_X1 U485 ( .A(KEYINPUT47), .ZN(n371) );
  XNOR2_X1 U486 ( .A(KEYINPUT15), .B(G902), .ZN(n624) );
  XNOR2_X1 U487 ( .A(n445), .B(n443), .ZN(n424) );
  NAND2_X1 U488 ( .A1(n651), .A2(n624), .ZN(n388) );
  XNOR2_X2 U489 ( .A(n732), .B(n389), .ZN(n651) );
  XNOR2_X1 U490 ( .A(n477), .B(n476), .ZN(n627) );
  XNOR2_X1 U491 ( .A(n386), .B(KEYINPUT39), .ZN(n573) );
  XNOR2_X1 U492 ( .A(n367), .B(KEYINPUT46), .ZN(n612) );
  NOR2_X2 U493 ( .A1(n639), .A2(n761), .ZN(n367) );
  NOR2_X1 U494 ( .A1(n570), .A2(n415), .ZN(n387) );
  XNOR2_X1 U495 ( .A(n510), .B(n363), .ZN(n374) );
  NOR2_X1 U496 ( .A1(n673), .A2(n610), .ZN(n611) );
  NAND2_X1 U497 ( .A1(n370), .A2(n665), .ZN(n603) );
  INV_X1 U498 ( .A(n757), .ZN(n368) );
  XNOR2_X2 U499 ( .A(n369), .B(G128), .ZN(n455) );
  NAND2_X1 U500 ( .A1(n588), .A2(n697), .ZN(n580) );
  XNOR2_X2 U501 ( .A(n478), .B(n479), .ZN(n697) );
  NAND2_X1 U502 ( .A1(n423), .A2(n422), .ZN(n421) );
  INV_X1 U503 ( .A(n680), .ZN(n577) );
  XNOR2_X1 U504 ( .A(n531), .B(KEYINPUT105), .ZN(n680) );
  NAND2_X1 U505 ( .A1(n372), .A2(n541), .ZN(n411) );
  XNOR2_X1 U506 ( .A(n559), .B(n373), .ZN(n372) );
  XNOR2_X1 U507 ( .A(n746), .B(n466), .ZN(n720) );
  INV_X1 U508 ( .A(n385), .ZN(n378) );
  NAND2_X1 U509 ( .A1(n385), .A2(n384), .ZN(n383) );
  INV_X1 U510 ( .A(n573), .ZN(n622) );
  NAND2_X1 U511 ( .A1(n417), .A2(n387), .ZN(n386) );
  XNOR2_X2 U512 ( .A(n475), .B(n425), .ZN(n732) );
  NAND2_X1 U513 ( .A1(n419), .A2(n390), .ZN(n561) );
  XNOR2_X1 U514 ( .A(n558), .B(n393), .ZN(n392) );
  INV_X1 U515 ( .A(KEYINPUT104), .ZN(n393) );
  NOR2_X1 U516 ( .A1(n651), .A2(n395), .ZN(n394) );
  INV_X1 U517 ( .A(n624), .ZN(n401) );
  OR2_X2 U518 ( .A1(n707), .A2(n601), .ZN(n585) );
  NOR2_X1 U519 ( .A1(n547), .A2(n549), .ZN(n531) );
  OR2_X2 U520 ( .A1(n738), .A2(n407), .ZN(n713) );
  NAND2_X1 U521 ( .A1(n623), .A2(KEYINPUT2), .ZN(n407) );
  XNOR2_X2 U522 ( .A(n561), .B(n560), .ZN(n738) );
  INV_X1 U523 ( .A(n541), .ZN(n759) );
  NAND2_X1 U524 ( .A1(n411), .A2(KEYINPUT64), .ZN(n423) );
  NOR2_X2 U525 ( .A1(n412), .A2(n738), .ZN(n711) );
  XNOR2_X1 U526 ( .A(n412), .B(n747), .ZN(n748) );
  INV_X1 U527 ( .A(n570), .ZN(n418) );
  NAND2_X1 U528 ( .A1(n678), .A2(n555), .ZN(n415) );
  INV_X1 U529 ( .A(n569), .ZN(n417) );
  NOR2_X1 U530 ( .A1(n416), .A2(n569), .ZN(n597) );
  NAND2_X1 U531 ( .A1(n418), .A2(n555), .ZN(n416) );
  INV_X1 U532 ( .A(KEYINPUT44), .ZN(n422) );
  INV_X1 U533 ( .A(n464), .ZN(n426) );
  INV_X1 U534 ( .A(n688), .ZN(n427) );
  INV_X1 U535 ( .A(n545), .ZN(n430) );
  INV_X1 U536 ( .A(n626), .ZN(n623) );
  XNOR2_X1 U537 ( .A(n464), .B(n465), .ZN(n466) );
  XNOR2_X1 U538 ( .A(KEYINPUT35), .B(KEYINPUT73), .ZN(n431) );
  INV_X1 U539 ( .A(KEYINPUT17), .ZN(n441) );
  INV_X1 U540 ( .A(KEYINPUT79), .ZN(n625) );
  XNOR2_X1 U541 ( .A(n437), .B(G122), .ZN(n439) );
  XNOR2_X1 U542 ( .A(n474), .B(n463), .ZN(n465) );
  INV_X1 U543 ( .A(KEYINPUT83), .ZN(n535) );
  INV_X1 U544 ( .A(KEYINPUT19), .ZN(n447) );
  INV_X1 U545 ( .A(n726), .ZN(n727) );
  XNOR2_X1 U546 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U547 ( .A(KEYINPUT86), .B(KEYINPUT70), .ZN(n432) );
  XNOR2_X1 U548 ( .A(G116), .B(KEYINPUT69), .ZN(n434) );
  XOR2_X1 U549 ( .A(KEYINPUT16), .B(KEYINPUT72), .Z(n437) );
  XNOR2_X1 U550 ( .A(n438), .B(G110), .ZN(n464) );
  XNOR2_X1 U551 ( .A(KEYINPUT65), .B(G101), .ZN(n460) );
  XOR2_X1 U552 ( .A(n440), .B(n460), .Z(n444) );
  NAND2_X1 U553 ( .A1(G224), .A2(n482), .ZN(n442) );
  XNOR2_X1 U554 ( .A(G146), .B(G125), .ZN(n481) );
  XNOR2_X1 U555 ( .A(n455), .B(n481), .ZN(n445) );
  NAND2_X1 U556 ( .A1(G210), .A2(n446), .ZN(n571) );
  NAND2_X1 U557 ( .A1(G214), .A2(n446), .ZN(n677) );
  XNOR2_X1 U558 ( .A(n448), .B(KEYINPUT14), .ZN(n449) );
  NAND2_X1 U559 ( .A1(G952), .A2(n449), .ZN(n706) );
  NOR2_X1 U560 ( .A1(G953), .A2(n706), .ZN(n566) );
  NAND2_X1 U561 ( .A1(G902), .A2(n449), .ZN(n563) );
  XNOR2_X1 U562 ( .A(G898), .B(KEYINPUT87), .ZN(n737) );
  NAND2_X1 U563 ( .A1(G953), .A2(n737), .ZN(n733) );
  NOR2_X1 U564 ( .A1(n563), .A2(n733), .ZN(n450) );
  NOR2_X1 U565 ( .A1(n566), .A2(n450), .ZN(n451) );
  XNOR2_X1 U566 ( .A(n451), .B(KEYINPUT88), .ZN(n452) );
  INV_X1 U567 ( .A(n533), .ZN(n550) );
  INV_X1 U568 ( .A(KEYINPUT90), .ZN(n459) );
  XOR2_X1 U569 ( .A(G137), .B(KEYINPUT67), .Z(n457) );
  XNOR2_X1 U570 ( .A(KEYINPUT4), .B(G131), .ZN(n456) );
  XNOR2_X1 U571 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U572 ( .A(G146), .B(n460), .ZN(n474) );
  XOR2_X1 U573 ( .A(G140), .B(KEYINPUT91), .Z(n462) );
  NAND2_X1 U574 ( .A1(G227), .A2(n482), .ZN(n461) );
  XNOR2_X1 U575 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U576 ( .A1(n720), .A2(G902), .ZN(n468) );
  INV_X1 U577 ( .A(G469), .ZN(n467) );
  XNOR2_X2 U578 ( .A(n468), .B(n467), .ZN(n555) );
  INV_X1 U579 ( .A(KEYINPUT1), .ZN(n469) );
  INV_X1 U580 ( .A(G472), .ZN(n479) );
  NAND2_X1 U581 ( .A1(n514), .A2(G210), .ZN(n470) );
  XNOR2_X1 U582 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U583 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U584 ( .A1(G902), .A2(n627), .ZN(n478) );
  XNOR2_X1 U585 ( .A(KEYINPUT10), .B(G140), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n744) );
  XNOR2_X1 U587 ( .A(n486), .B(n485), .ZN(n489) );
  XNOR2_X1 U588 ( .A(n487), .B(KEYINPUT92), .ZN(n488) );
  XNOR2_X1 U589 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U590 ( .A1(n624), .A2(G234), .ZN(n492) );
  INV_X1 U591 ( .A(KEYINPUT20), .ZN(n491) );
  XNOR2_X1 U592 ( .A(n492), .B(n491), .ZN(n498) );
  INV_X1 U593 ( .A(G217), .ZN(n493) );
  OR2_X1 U594 ( .A1(n498), .A2(n493), .ZN(n494) );
  XNOR2_X1 U595 ( .A(n494), .B(KEYINPUT25), .ZN(n495) );
  XNOR2_X2 U596 ( .A(n496), .B(n495), .ZN(n688) );
  INV_X1 U597 ( .A(G221), .ZN(n497) );
  OR2_X1 U598 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U599 ( .A(n499), .B(KEYINPUT21), .ZN(n687) );
  INV_X1 U600 ( .A(KEYINPUT66), .ZN(n500) );
  XNOR2_X2 U601 ( .A(n501), .B(n500), .ZN(n690) );
  XNOR2_X1 U602 ( .A(KEYINPUT108), .B(KEYINPUT33), .ZN(n502) );
  NOR2_X1 U603 ( .A1(n554), .A2(n676), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n503), .B(KEYINPUT34), .ZN(n529) );
  XOR2_X1 U605 ( .A(KEYINPUT101), .B(G122), .Z(n505) );
  XNOR2_X1 U606 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U607 ( .A(KEYINPUT99), .B(KEYINPUT7), .ZN(n506) );
  XNOR2_X1 U608 ( .A(n507), .B(n354), .ZN(n509) );
  NOR2_X1 U609 ( .A1(n726), .A2(G902), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n511), .B(KEYINPUT102), .ZN(n513) );
  INV_X1 U611 ( .A(G478), .ZN(n512) );
  XNOR2_X1 U612 ( .A(n513), .B(n512), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n514), .A2(G214), .ZN(n515) );
  XNOR2_X1 U614 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U615 ( .A(n517), .B(KEYINPUT11), .Z(n519) );
  XNOR2_X1 U616 ( .A(n519), .B(n518), .ZN(n524) );
  XNOR2_X1 U617 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U618 ( .A(n744), .B(n522), .ZN(n523) );
  XNOR2_X1 U619 ( .A(n524), .B(n523), .ZN(n645) );
  NAND2_X1 U620 ( .A1(n645), .A2(n525), .ZN(n527) );
  XOR2_X1 U621 ( .A(KEYINPUT13), .B(G475), .Z(n526) );
  XNOR2_X1 U622 ( .A(n527), .B(n526), .ZN(n547) );
  NAND2_X1 U623 ( .A1(n549), .A2(n547), .ZN(n595) );
  XOR2_X1 U624 ( .A(n595), .B(KEYINPUT74), .Z(n528) );
  NAND2_X1 U625 ( .A1(n529), .A2(n528), .ZN(n530) );
  INV_X1 U626 ( .A(n687), .ZN(n579) );
  AND2_X1 U627 ( .A1(n579), .A2(n577), .ZN(n532) );
  NAND2_X1 U628 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n552), .B(n535), .ZN(n594) );
  NOR2_X1 U630 ( .A1(n594), .A2(n589), .ZN(n536) );
  NAND2_X1 U631 ( .A1(n688), .A2(n536), .ZN(n537) );
  XNOR2_X2 U632 ( .A(n538), .B(KEYINPUT32), .ZN(n760) );
  INV_X1 U633 ( .A(n552), .ZN(n691) );
  NOR2_X1 U634 ( .A1(n697), .A2(n691), .ZN(n539) );
  NAND2_X1 U635 ( .A1(n688), .A2(n539), .ZN(n540) );
  OR2_X1 U636 ( .A1(n545), .A2(n540), .ZN(n662) );
  NAND2_X1 U637 ( .A1(KEYINPUT64), .A2(n559), .ZN(n542) );
  NAND2_X1 U638 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n543), .A2(KEYINPUT44), .ZN(n544) );
  INV_X1 U640 ( .A(n547), .ZN(n548) );
  XNOR2_X1 U641 ( .A(n670), .B(KEYINPUT103), .ZN(n621) );
  OR2_X1 U642 ( .A1(n549), .A2(n548), .ZN(n656) );
  INV_X1 U643 ( .A(n550), .ZN(n553) );
  NAND2_X1 U644 ( .A1(n697), .A2(n690), .ZN(n551) );
  NAND2_X1 U645 ( .A1(n555), .A2(n690), .ZN(n556) );
  INV_X1 U646 ( .A(KEYINPUT45), .ZN(n560) );
  NAND2_X1 U647 ( .A1(n697), .A2(n677), .ZN(n562) );
  XNOR2_X1 U648 ( .A(n562), .B(KEYINPUT30), .ZN(n570) );
  OR2_X1 U649 ( .A1(n482), .A2(n563), .ZN(n564) );
  NOR2_X1 U650 ( .A1(G900), .A2(n564), .ZN(n565) );
  OR2_X1 U651 ( .A1(n566), .A2(n565), .ZN(n568) );
  INV_X1 U652 ( .A(KEYINPUT75), .ZN(n567) );
  XNOR2_X1 U653 ( .A(n568), .B(n567), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n690), .A2(n586), .ZN(n569) );
  INV_X1 U655 ( .A(n656), .ZN(n572) );
  NAND2_X1 U656 ( .A1(n573), .A2(n572), .ZN(n576) );
  INV_X1 U657 ( .A(KEYINPUT110), .ZN(n574) );
  XNOR2_X1 U658 ( .A(n574), .B(KEYINPUT40), .ZN(n575) );
  XNOR2_X1 U659 ( .A(n576), .B(n575), .ZN(n639) );
  NAND2_X1 U660 ( .A1(n678), .A2(n677), .ZN(n681) );
  XNOR2_X1 U661 ( .A(n578), .B(KEYINPUT41), .ZN(n707) );
  INV_X1 U662 ( .A(n586), .ZN(n581) );
  AND2_X1 U663 ( .A1(n688), .A2(n579), .ZN(n588) );
  NOR2_X1 U664 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U665 ( .A(KEYINPUT28), .B(n582), .ZN(n583) );
  NAND2_X1 U666 ( .A1(n555), .A2(n583), .ZN(n601) );
  INV_X1 U667 ( .A(KEYINPUT42), .ZN(n584) );
  XNOR2_X2 U668 ( .A(n585), .B(n584), .ZN(n761) );
  NAND2_X1 U669 ( .A1(n586), .A2(n677), .ZN(n587) );
  NOR2_X1 U670 ( .A1(n656), .A2(n587), .ZN(n591) );
  AND2_X1 U671 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n614) );
  NOR2_X1 U673 ( .A1(n617), .A2(n614), .ZN(n592) );
  XOR2_X1 U674 ( .A(KEYINPUT36), .B(n592), .Z(n593) );
  NOR2_X1 U675 ( .A1(n594), .A2(n593), .ZN(n673) );
  NOR2_X1 U676 ( .A1(n617), .A2(n595), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n599) );
  INV_X1 U678 ( .A(KEYINPUT109), .ZN(n598) );
  XNOR2_X1 U679 ( .A(n599), .B(n598), .ZN(n758) );
  NAND2_X1 U680 ( .A1(n371), .A2(KEYINPUT78), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n371), .A2(n665), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n604), .A2(KEYINPUT78), .ZN(n606) );
  INV_X1 U684 ( .A(n682), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n607) );
  AND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n758), .A2(n609), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n691), .A2(n614), .ZN(n616) );
  INV_X1 U690 ( .A(KEYINPUT43), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n616), .B(n615), .ZN(n618) );
  AND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n675) );
  INV_X1 U693 ( .A(n675), .ZN(n619) );
  INV_X1 U694 ( .A(KEYINPUT80), .ZN(n620) );
  OR2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n637) );
  NAND2_X1 U696 ( .A1(n725), .A2(G472), .ZN(n630) );
  XNOR2_X1 U697 ( .A(n627), .B(KEYINPUT62), .ZN(n628) );
  XNOR2_X1 U698 ( .A(n628), .B(KEYINPUT111), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n634) );
  INV_X1 U700 ( .A(G952), .ZN(n631) );
  NAND2_X1 U701 ( .A1(n631), .A2(G953), .ZN(n633) );
  INV_X1 U702 ( .A(KEYINPUT85), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(n729) );
  NAND2_X1 U704 ( .A1(n634), .A2(n729), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U706 ( .A(G134), .B(KEYINPUT116), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(G36) );
  XNOR2_X1 U708 ( .A(G131), .B(KEYINPUT127), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(G33) );
  NAND2_X1 U710 ( .A1(n725), .A2(G217), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n642) );
  INV_X1 U712 ( .A(n729), .ZN(n724) );
  NOR2_X1 U713 ( .A1(n642), .A2(n724), .ZN(G66) );
  NAND2_X1 U714 ( .A1(n725), .A2(G475), .ZN(n647) );
  XNOR2_X1 U715 ( .A(KEYINPUT84), .B(KEYINPUT120), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(KEYINPUT59), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X2 U719 ( .A1(n648), .A2(n724), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U721 ( .A1(n725), .A2(G210), .ZN(n653) );
  XNOR2_X1 U722 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X2 U725 ( .A1(n654), .A2(n724), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U727 ( .A1(n355), .A2(n572), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(G104), .ZN(G6) );
  XOR2_X1 U729 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n659) );
  NAND2_X1 U730 ( .A1(n355), .A2(n670), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(n661) );
  XOR2_X1 U732 ( .A(G107), .B(KEYINPUT27), .Z(n660) );
  XNOR2_X1 U733 ( .A(n661), .B(n660), .ZN(G9) );
  XNOR2_X1 U734 ( .A(G110), .B(n662), .ZN(G12) );
  XOR2_X1 U735 ( .A(G128), .B(KEYINPUT29), .Z(n664) );
  NAND2_X1 U736 ( .A1(n665), .A2(n670), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(G30) );
  NAND2_X1 U738 ( .A1(n665), .A2(n572), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n666), .B(KEYINPUT114), .ZN(n667) );
  XNOR2_X1 U740 ( .A(G146), .B(n667), .ZN(G48) );
  NAND2_X1 U741 ( .A1(n669), .A2(n572), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n668), .B(G113), .ZN(G15) );
  XOR2_X1 U743 ( .A(G116), .B(KEYINPUT115), .Z(n672) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(G18) );
  XNOR2_X1 U746 ( .A(G125), .B(n673), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n674), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U748 ( .A(G140), .B(n675), .Z(G42) );
  NOR2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U753 ( .A(KEYINPUT119), .B(n685), .Z(n686) );
  NOR2_X1 U754 ( .A1(n676), .A2(n686), .ZN(n703) );
  NAND2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U756 ( .A(KEYINPUT49), .B(n689), .Z(n695) );
  XOR2_X1 U757 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n693) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U759 ( .A(n693), .B(n692), .Z(n694) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U762 ( .A1(n356), .A2(n698), .ZN(n699) );
  XOR2_X1 U763 ( .A(n699), .B(KEYINPUT51), .Z(n700) );
  XNOR2_X1 U764 ( .A(KEYINPUT118), .B(n700), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n707), .A2(n701), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U767 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n676), .A2(n707), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n716) );
  XOR2_X1 U771 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n710) );
  NOR2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U773 ( .A(KEYINPUT76), .B(n712), .Z(n714) );
  NAND2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U775 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U776 ( .A1(n717), .A2(G953), .ZN(n718) );
  XNOR2_X1 U777 ( .A(n718), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U778 ( .A1(n725), .A2(G469), .ZN(n722) );
  XOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n719) );
  NOR2_X1 U780 ( .A1(n724), .A2(n723), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n725), .A2(G478), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT121), .ZN(G63) );
  XNOR2_X1 U785 ( .A(n732), .B(G101), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n734), .A2(n733), .ZN(n743) );
  NAND2_X1 U787 ( .A1(G953), .A2(G224), .ZN(n735) );
  XOR2_X1 U788 ( .A(KEYINPUT61), .B(n735), .Z(n736) );
  NOR2_X1 U789 ( .A1(n737), .A2(n736), .ZN(n741) );
  NOR2_X1 U790 ( .A1(G953), .A2(n738), .ZN(n739) );
  XNOR2_X1 U791 ( .A(n739), .B(KEYINPUT122), .ZN(n740) );
  NOR2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n744), .B(KEYINPUT123), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n746), .B(n745), .ZN(n750) );
  XOR2_X1 U796 ( .A(n750), .B(KEYINPUT124), .Z(n747) );
  NOR2_X1 U797 ( .A1(n748), .A2(G953), .ZN(n749) );
  XNOR2_X1 U798 ( .A(n749), .B(KEYINPUT125), .ZN(n755) );
  XNOR2_X1 U799 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U800 ( .A1(n751), .A2(G900), .ZN(n752) );
  XNOR2_X1 U801 ( .A(KEYINPUT126), .B(n752), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(G953), .ZN(n754) );
  NAND2_X1 U803 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U804 ( .A(G101), .B(KEYINPUT112), .Z(n756) );
  XNOR2_X1 U805 ( .A(n757), .B(n756), .ZN(G3) );
  XNOR2_X1 U806 ( .A(G143), .B(n758), .ZN(G45) );
  XOR2_X1 U807 ( .A(G122), .B(n759), .Z(G24) );
  XNOR2_X1 U808 ( .A(G119), .B(n760), .ZN(G21) );
  XOR2_X1 U809 ( .A(n761), .B(G137), .Z(G39) );
endmodule

