//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n217), .B1(new_n201), .B2(new_n218), .C1(new_n206), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n210), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n210), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT64), .Z(new_n233));
  AOI21_X1  g0033(.A(new_n228), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  AND3_X1   g0034(.A1(new_n224), .A2(new_n225), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n229), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n230), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n261), .A2(new_n262), .B1(G20), .B2(new_n204), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n255), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G13), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n266), .A2(new_n230), .A3(G1), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n254), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G50), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n267), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(G50), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g0074(.A(new_n274), .B(KEYINPUT9), .Z(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G222), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G223), .A2(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n229), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n280), .B(new_n282), .C1(G77), .C2(new_n276), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT68), .B1(new_n281), .B2(new_n229), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT68), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(G1), .A4(G13), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n286), .A3(G274), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n285), .A3(new_n289), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n283), .B(new_n290), .C1(new_n218), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(G200), .B2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n275), .A2(new_n298), .A3(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n268), .ZN(new_n302));
  INV_X1    g0102(.A(new_n256), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n270), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n302), .A2(new_n304), .B1(new_n272), .B2(new_n303), .ZN(new_n305));
  XNOR2_X1  g0105(.A(G58), .B(G68), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n306), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT74), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n312));
  AOI21_X1  g0112(.A(G20), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n308), .B1(new_n313), .B2(KEYINPUT7), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT7), .ZN(new_n315));
  OAI211_X1 g0115(.A(KEYINPUT74), .B(new_n315), .C1(new_n276), .C2(G20), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(G20), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n310), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n309), .A2(KEYINPUT75), .A3(G33), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n312), .A3(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n314), .A2(new_n316), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n307), .B1(new_n322), .B2(new_n203), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n255), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n311), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT72), .B1(new_n311), .B2(KEYINPUT3), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n310), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT73), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n317), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n311), .A2(KEYINPUT3), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT72), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n309), .B2(G33), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n311), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n315), .B1(new_n335), .B2(G20), .ZN(new_n336));
  INV_X1    g0136(.A(new_n317), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT73), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n330), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G68), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(KEYINPUT16), .A3(new_n307), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n305), .B1(new_n325), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n333), .A2(new_n334), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G223), .A2(G1698), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n218), .B2(G1698), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n345), .A3(new_n310), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n282), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n284), .A2(G232), .A3(new_n285), .A4(new_n289), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n290), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  INV_X1    g0154(.A(new_n282), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n346), .B2(new_n347), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n290), .A2(new_n351), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT76), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n356), .A2(new_n357), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n342), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT18), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n314), .A2(new_n316), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n321), .A2(new_n317), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n203), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n307), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n324), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n341), .A2(new_n370), .A3(new_n254), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n353), .A2(new_n372), .A3(new_n358), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n293), .A2(KEYINPUT77), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n293), .A2(KEYINPUT77), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n360), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n305), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n371), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n365), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT71), .B1(new_n272), .B2(G68), .ZN(new_n384));
  XOR2_X1   g0184(.A(new_n384), .B(KEYINPUT12), .Z(new_n385));
  NAND3_X1  g0185(.A1(new_n268), .A2(G68), .A3(new_n270), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n260), .A2(new_n201), .B1(new_n230), .B2(G68), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n257), .A2(new_n212), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n254), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g0190(.A(new_n390), .B(KEYINPUT11), .Z(new_n391));
  NOR2_X1   g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n284), .A2(G238), .A3(new_n285), .A4(new_n289), .ZN(new_n394));
  NOR2_X1   g0194(.A1(G226), .A2(G1698), .ZN(new_n395));
  INV_X1    g0195(.A(G232), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(G1698), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n276), .B1(G33), .B2(G97), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n290), .B(new_n394), .C1(new_n398), .C2(new_n355), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT13), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G169), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n401), .A2(KEYINPUT14), .B1(new_n361), .B2(new_n400), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n393), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(G200), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n392), .B(new_n405), .C1(new_n293), .C2(new_n400), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT15), .B(G87), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n408), .A2(new_n257), .B1(new_n230), .B2(new_n212), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n256), .A2(new_n260), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n254), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n270), .A2(G77), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT70), .B1(new_n267), .B2(new_n212), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n267), .A2(KEYINPUT70), .A3(new_n212), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OAI221_X1 g0215(.A(new_n411), .B1(new_n302), .B2(new_n412), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G238), .A2(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n276), .B(new_n417), .C1(new_n396), .C2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n282), .C1(G107), .C2(new_n276), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n290), .C1(new_n213), .C2(new_n291), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n420), .B2(G200), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n293), .B2(new_n420), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n354), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n416), .C1(G179), .C2(new_n420), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n292), .A2(new_n354), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n426), .B1(G179), .B2(new_n292), .C1(new_n265), .C2(new_n273), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n301), .A2(new_n383), .A3(new_n407), .A4(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT21), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n269), .A2(G33), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n268), .A2(G116), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G116), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n267), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G283), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT80), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n436), .B(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(KEYINPUT78), .A2(G97), .ZN(new_n439));
  NAND2_X1  g0239(.A1(KEYINPUT78), .A2(G97), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(new_n230), .C1(new_n441), .C2(G33), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n255), .B1(G20), .B2(new_n433), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT20), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(KEYINPUT20), .A3(new_n443), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n435), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n284), .A2(G274), .A3(new_n289), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  INV_X1    g0250(.A(G41), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT5), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G41), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n455), .A2(new_n284), .A3(new_n289), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G270), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  MUX2_X1   g0259(.A(G257), .B(G264), .S(G1698), .Z(new_n460));
  INV_X1    g0260(.A(new_n276), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n335), .A2(new_n460), .B1(new_n461), .B2(G303), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n355), .ZN(new_n463));
  OAI21_X1  g0263(.A(G169), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n430), .B1(new_n447), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n459), .A2(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n376), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n467), .B(new_n447), .C1(new_n372), .C2(new_n466), .ZN(new_n468));
  INV_X1    g0268(.A(new_n446), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n434), .B(new_n432), .C1(new_n469), .C2(new_n444), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G179), .A3(new_n466), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n459), .A2(new_n463), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT21), .A4(G169), .ZN(new_n473));
  AND4_X1   g0273(.A1(new_n465), .A2(new_n468), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n335), .A2(new_n230), .A3(G68), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n441), .B2(new_n257), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G97), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n230), .B1(new_n478), .B2(new_n476), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n439), .A2(new_n214), .A3(new_n207), .A4(new_n440), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n475), .B(new_n477), .C1(new_n481), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n254), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT83), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n268), .A2(new_n431), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(new_n408), .ZN(new_n489));
  INV_X1    g0289(.A(new_n408), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n268), .A2(KEYINPUT83), .A3(new_n490), .A4(new_n431), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n408), .A2(new_n267), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OR3_X1    g0294(.A1(new_n449), .A2(G1), .A3(G274), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n215), .B1(new_n449), .B2(G1), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n284), .A2(new_n495), .A3(new_n289), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(G238), .A2(G1698), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n213), .B2(G1698), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n335), .A2(new_n499), .B1(G33), .B2(G116), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(new_n355), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n354), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G179), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(G200), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n293), .B2(new_n501), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n268), .A2(G87), .A3(new_n431), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n486), .A2(new_n493), .A3(new_n506), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n494), .A2(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n474), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n267), .A2(new_n207), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT25), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n207), .B2(new_n488), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G20), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n230), .B2(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n230), .A2(KEYINPUT22), .A3(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n230), .A2(G87), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n461), .A2(new_n523), .ZN(new_n524));
  OAI221_X1 g0324(.A(new_n521), .B1(new_n328), .B2(new_n522), .C1(new_n524), .C2(KEYINPUT22), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT84), .A2(KEYINPUT24), .ZN(new_n526));
  OR2_X1    g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n255), .B1(new_n525), .B2(new_n526), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n514), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n457), .A2(G264), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G250), .A2(G1698), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n219), .B2(G1698), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n335), .A2(new_n532), .B1(G33), .B2(G294), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n456), .B(new_n530), .C1(new_n355), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT85), .B1(new_n534), .B2(G169), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n534), .A2(new_n361), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(KEYINPUT85), .A3(G169), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n529), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n534), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(KEYINPUT86), .A3(new_n293), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n534), .A2(new_n372), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT86), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n534), .B2(G190), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n529), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n457), .A2(G257), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n456), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n276), .A2(G244), .A3(new_n277), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n213), .A2(KEYINPUT4), .A3(G1698), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n551), .A2(KEYINPUT4), .B1(new_n335), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G250), .A2(G1698), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n438), .B1(new_n461), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT81), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n355), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n553), .A2(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT81), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n550), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n361), .ZN(new_n562));
  INV_X1    g0362(.A(new_n550), .ZN(new_n563));
  INV_X1    g0363(.A(new_n560), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n282), .B1(new_n559), .B2(KEYINPUT81), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n354), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n568));
  XOR2_X1   g0368(.A(G97), .B(G107), .Z(new_n569));
  OAI22_X1  g0369(.A1(new_n441), .A2(new_n568), .B1(new_n569), .B2(KEYINPUT6), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n322), .B2(new_n207), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n254), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n267), .A2(new_n206), .ZN(new_n574));
  XOR2_X1   g0374(.A(new_n574), .B(KEYINPUT79), .Z(new_n575));
  NOR2_X1   g0375(.A1(new_n488), .A2(new_n206), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n562), .A2(new_n567), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n573), .A2(new_n577), .ZN(new_n580));
  OAI211_X1 g0380(.A(G190), .B(new_n563), .C1(new_n564), .C2(new_n565), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n561), .C2(new_n372), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n510), .A2(new_n548), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n429), .A2(new_n584), .ZN(G372));
  INV_X1    g0385(.A(KEYINPUT90), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n300), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT90), .B1(new_n297), .B2(new_n299), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT17), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n381), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g0390(.A(new_n424), .B(KEYINPUT89), .Z(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n406), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n590), .B1(new_n592), .B2(new_n404), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n371), .A2(new_n380), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT88), .ZN(new_n595));
  INV_X1    g0395(.A(new_n363), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT88), .B1(new_n342), .B2(new_n363), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT18), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT18), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n587), .A2(new_n588), .B1(new_n593), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n429), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n580), .B1(new_n354), .B2(new_n566), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n505), .A2(new_n507), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(KEYINPUT26), .A3(new_n562), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(new_n502), .C1(G179), .C2(new_n501), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n605), .A2(KEYINPUT87), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n508), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n582), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n473), .A2(new_n465), .A3(new_n471), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n547), .B1(new_n539), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n579), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n606), .B1(new_n615), .B2(KEYINPUT26), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(new_n608), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n602), .B(new_n427), .C1(new_n603), .C2(new_n617), .ZN(G369));
  NAND3_X1  g0418(.A1(new_n269), .A2(new_n230), .A3(G13), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(G213), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n470), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n474), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n473), .A2(new_n465), .A3(new_n471), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n625), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(G330), .ZN(new_n629));
  INV_X1    g0429(.A(new_n624), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n529), .A2(new_n630), .ZN(new_n631));
  OAI22_X1  g0431(.A1(new_n548), .A2(new_n631), .B1(new_n540), .B2(new_n630), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n547), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n539), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n627), .A2(new_n624), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n635), .A2(new_n636), .B1(new_n539), .B2(new_n630), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(G399));
  INV_X1    g0438(.A(new_n226), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G41), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G1), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n483), .A2(G116), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n642), .A2(new_n643), .B1(new_n232), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT28), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n508), .A2(KEYINPUT26), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n608), .B1(new_n646), .B2(new_n579), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n604), .A2(new_n562), .A3(new_n609), .A4(new_n611), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(KEYINPUT26), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n539), .A2(new_n613), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT93), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n611), .A2(new_n547), .A3(new_n609), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n583), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n630), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT29), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n624), .B1(new_n616), .B2(new_n608), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT29), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT30), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n533), .A2(new_n355), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n530), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(new_n501), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(G179), .A3(new_n466), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n661), .B1(new_n665), .B2(new_n566), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n472), .A2(new_n361), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n561), .A2(KEYINPUT30), .A3(new_n667), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT92), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n561), .A2(new_n667), .A3(new_n664), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT92), .B1(new_n671), .B2(new_n661), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT91), .B1(new_n561), .B2(new_n541), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n566), .A2(new_n675), .A3(new_n534), .ZN(new_n676));
  INV_X1    g0476(.A(new_n501), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n466), .A2(G179), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n670), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n624), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n583), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n627), .A2(new_n509), .A3(new_n468), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n635), .A4(new_n630), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n679), .A2(new_n666), .A3(new_n668), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n630), .A2(new_n682), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n660), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n645), .B1(new_n693), .B2(G1), .ZN(G364));
  NOR2_X1   g0494(.A1(new_n266), .A2(G20), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n269), .B1(new_n695), .B2(G45), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n640), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n629), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(G330), .B2(new_n628), .ZN(new_n700));
  INV_X1    g0500(.A(new_n698), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n229), .B1(G20), .B2(new_n354), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n230), .A2(new_n361), .A3(new_n372), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n376), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n230), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n705), .A2(new_n201), .B1(new_n206), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n372), .A2(G179), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n710), .A2(new_n230), .A3(new_n293), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n461), .B1(new_n711), .B2(G87), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n230), .A2(new_n361), .A3(G200), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n376), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n293), .A2(G20), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT96), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n710), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n712), .B1(new_n714), .B2(new_n202), .C1(new_n718), .C2(new_n207), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n713), .A2(new_n293), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n708), .B(new_n719), .C1(G77), .C2(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n716), .A2(G179), .A3(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G159), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT32), .Z(new_n724));
  AND3_X1   g0524(.A1(new_n704), .A2(KEYINPUT97), .A3(new_n293), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT97), .B1(new_n704), .B2(new_n293), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n721), .B(new_n724), .C1(new_n203), .C2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n705), .ZN(new_n729));
  INV_X1    g0529(.A(new_n707), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n729), .A2(G326), .B1(G294), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G322), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n714), .ZN(new_n733));
  INV_X1    g0533(.A(new_n727), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT33), .B(G317), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n722), .A2(G329), .ZN(new_n737));
  INV_X1    g0537(.A(new_n720), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  INV_X1    g0539(.A(G303), .ZN(new_n740));
  INV_X1    g0540(.A(new_n711), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n461), .B1(new_n738), .B2(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(G283), .B2(new_n717), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n736), .A2(new_n737), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n703), .B1(new_n728), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n266), .A2(new_n311), .A3(KEYINPUT95), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G13), .B2(G33), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n702), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n335), .A2(new_n639), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n233), .A2(new_n449), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n753), .B(new_n754), .C1(new_n248), .C2(new_n449), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G355), .A2(KEYINPUT94), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n461), .A2(new_n639), .ZN(new_n757));
  NAND2_X1  g0557(.A1(G355), .A2(KEYINPUT94), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n755), .B1(G116), .B2(new_n226), .C1(new_n756), .C2(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n701), .B(new_n745), .C1(new_n752), .C2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT98), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n751), .B(KEYINPUT99), .Z(new_n763));
  NOR2_X1   g0563(.A1(new_n628), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n700), .B1(new_n762), .B2(new_n764), .ZN(G396));
  NAND2_X1  g0565(.A1(new_n416), .A2(new_n624), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n591), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n425), .A2(KEYINPUT102), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n422), .A2(new_n424), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n766), .B1(new_n770), .B2(KEYINPUT102), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n657), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n701), .B1(new_n773), .B2(new_n691), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(KEYINPUT103), .B1(new_n691), .B2(new_n773), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(KEYINPUT103), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n749), .A2(new_n702), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n701), .B1(new_n212), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n714), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G143), .B1(G159), .B2(new_n720), .ZN(new_n780));
  INV_X1    g0580(.A(G137), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n780), .B1(new_n781), .B2(new_n705), .C1(new_n258), .C2(new_n727), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT34), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n335), .B1(new_n202), .B2(new_n707), .C1(new_n741), .C2(new_n201), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n718), .A2(new_n203), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(G132), .C2(new_n722), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n717), .A2(G87), .ZN(new_n788));
  INV_X1    g0588(.A(new_n722), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n739), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT100), .Z(new_n791));
  INV_X1    g0591(.A(G294), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n433), .A2(new_n738), .B1(new_n714), .B2(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n461), .B1(new_n206), .B2(new_n707), .C1(new_n741), .C2(new_n207), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(G303), .C2(new_n729), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n727), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n787), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n799), .A2(KEYINPUT101), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n702), .B1(new_n799), .B2(KEYINPUT101), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n778), .B1(new_n800), .B2(new_n801), .C1(new_n772), .C2(new_n750), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n776), .A2(new_n802), .ZN(G384));
  OR2_X1    g0603(.A1(new_n570), .A2(KEYINPUT35), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n570), .A2(KEYINPUT35), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n804), .A2(G116), .A3(new_n231), .A4(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT36), .Z(new_n807));
  INV_X1    g0607(.A(new_n232), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n808), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n201), .A2(G68), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n269), .B(G13), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n341), .A2(new_n254), .ZN(new_n813));
  AOI21_X1  g0613(.A(KEYINPUT16), .B1(new_n340), .B2(new_n307), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n380), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n596), .ZN(new_n816));
  INV_X1    g0616(.A(new_n622), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n816), .A2(new_n818), .A3(new_n381), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT37), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n364), .A2(KEYINPUT37), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n594), .A2(new_n817), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n821), .A2(new_n381), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n818), .B1(new_n365), .B2(new_n382), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT39), .B1(new_n827), .B2(KEYINPUT38), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT106), .ZN(new_n829));
  XNOR2_X1  g0629(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n382), .B1(new_n599), .B2(new_n600), .ZN(new_n831));
  INV_X1    g0631(.A(new_n822), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n381), .B1(new_n342), .B2(new_n622), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n598), .B2(new_n597), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n823), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n829), .B(new_n830), .C1(new_n833), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT18), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n595), .B1(new_n594), .B2(new_n596), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n342), .A2(KEYINPUT88), .A3(new_n363), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT18), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n590), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n837), .B1(new_n844), .B2(new_n822), .ZN(new_n845));
  INV_X1    g0645(.A(new_n830), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT106), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n828), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT107), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT107), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n828), .B(new_n850), .C1(new_n838), .C2(new_n847), .ZN(new_n851));
  INV_X1    g0651(.A(new_n818), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n383), .A2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n853), .A2(KEYINPUT38), .A3(new_n824), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT38), .B1(new_n853), .B2(new_n824), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT39), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n849), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n404), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n630), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n424), .A2(new_n624), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n657), .B2(new_n772), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n854), .A2(new_n855), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n404), .B(new_n406), .C1(new_n392), .C2(new_n630), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n393), .B(new_n624), .C1(new_n402), .C2(new_n403), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT104), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n863), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n601), .B2(new_n622), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n603), .B1(new_n656), .B2(new_n659), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n602), .A2(new_n427), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n873), .B(new_n876), .Z(new_n877));
  INV_X1    g0677(.A(new_n854), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n838), .B2(new_n847), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n868), .A2(new_n869), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n680), .A2(new_n688), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT92), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n666), .B2(new_n668), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(new_n672), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n630), .B1(new_n884), .B2(new_n679), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n881), .B(new_n686), .C1(new_n885), .C2(KEYINPUT31), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n880), .A2(new_n886), .A3(KEYINPUT40), .A4(new_n772), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n879), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n880), .A2(new_n886), .A3(new_n772), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n864), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n429), .A2(new_n886), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(G330), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n877), .A2(KEYINPUT108), .A3(new_n897), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n898), .B1(new_n269), .B2(new_n695), .C1(new_n877), .C2(new_n897), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT108), .B1(new_n877), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n812), .B1(new_n899), .B2(new_n900), .ZN(G367));
  AND2_X1   g0701(.A1(new_n507), .A2(new_n624), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n609), .A2(new_n611), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n608), .B2(new_n903), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT110), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n579), .B(new_n582), .C1(new_n580), .C2(new_n630), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n579), .B2(new_n630), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n635), .A3(new_n636), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n909), .A2(new_n540), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n624), .B1(new_n914), .B2(new_n579), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT109), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n908), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n633), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n910), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n906), .A2(new_n907), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n640), .B(KEYINPUT41), .Z(new_n925));
  NAND2_X1  g0725(.A1(new_n635), .A2(new_n636), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n632), .B2(new_n636), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n629), .B(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n660), .A2(new_n691), .A3(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT112), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n910), .A2(new_n637), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT45), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n910), .A2(new_n637), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT44), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n910), .A2(new_n637), .A3(KEYINPUT44), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n633), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT111), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n937), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n920), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n929), .A2(KEYINPUT112), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n939), .A3(new_n920), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n930), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n925), .B1(new_n946), .B2(new_n693), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n924), .B1(new_n947), .B2(new_n697), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n752), .B1(new_n226), .B2(new_n408), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n244), .B2(new_n753), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n741), .A2(new_n433), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n951), .A2(KEYINPUT46), .B1(G107), .B2(new_n730), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n740), .B2(new_n714), .C1(new_n727), .C2(new_n792), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n729), .A2(G311), .B1(new_n720), .B2(G283), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n439), .A2(new_n440), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n722), .A2(G317), .B1(new_n717), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n954), .A2(new_n328), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n276), .B1(new_n741), .B2(new_n202), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G50), .B2(new_n720), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n717), .A2(G77), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n781), .C2(new_n789), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n729), .A2(G143), .B1(G68), .B2(new_n730), .ZN(new_n963));
  INV_X1    g0763(.A(G159), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n963), .B1(new_n258), .B2(new_n714), .C1(new_n727), .C2(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n953), .A2(new_n958), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n701), .B(new_n950), .C1(new_n967), .C2(new_n702), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n905), .B2(new_n763), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n948), .A2(new_n969), .ZN(G387));
  NOR2_X1   g0770(.A1(new_n632), .A2(new_n763), .ZN(new_n971));
  INV_X1    g0771(.A(new_n753), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n241), .B2(G45), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n643), .B2(new_n757), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n303), .A2(new_n201), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n449), .B1(new_n203), .B2(new_n212), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n976), .A2(new_n643), .A3(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n974), .A2(new_n978), .B1(G107), .B2(new_n226), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n752), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n698), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n707), .A2(new_n408), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n203), .A2(new_n738), .B1(new_n705), .B2(new_n964), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G50), .C2(new_n779), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n722), .A2(G150), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n335), .B1(new_n741), .B2(new_n212), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G97), .B2(new_n717), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n734), .A2(new_n303), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G317), .A2(new_n779), .B1(new_n729), .B2(G322), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n740), .B2(new_n738), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G311), .B2(new_n734), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT113), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT48), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n741), .A2(new_n792), .B1(new_n796), .B2(new_n707), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n335), .B1(new_n722), .B2(G326), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n433), .C2(new_n718), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n998), .A2(KEYINPUT49), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n989), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n971), .B(new_n981), .C1(new_n1003), .C2(new_n702), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(new_n697), .B2(new_n928), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n930), .A2(new_n944), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n640), .B1(new_n693), .B2(new_n928), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(G393));
  AND2_X1   g0808(.A1(new_n942), .A2(new_n938), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n640), .B(new_n946), .C1(new_n1006), .C2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n909), .B(new_n751), .C1(new_n579), .C2(new_n630), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n752), .B1(new_n226), .B2(new_n441), .C1(new_n251), .C2(new_n972), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n698), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n461), .B1(new_n738), .B2(new_n792), .C1(new_n796), .C2(new_n741), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G116), .B2(new_n730), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n722), .A2(G322), .B1(new_n717), .B2(G107), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n740), .C2(new_n727), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G311), .A2(new_n779), .B1(new_n729), .B2(G317), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n722), .A2(G143), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G77), .A2(new_n730), .B1(new_n720), .B2(new_n303), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n328), .B1(new_n711), .B2(G68), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n788), .A4(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n258), .A2(new_n705), .B1(new_n714), .B2(new_n964), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1025), .A2(new_n1027), .B1(new_n734), .B2(G50), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1017), .A2(new_n1020), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1013), .B1(new_n1030), .B2(new_n702), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1009), .A2(new_n697), .B1(new_n1011), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1010), .A2(new_n1032), .ZN(G390));
  NOR2_X1   g0833(.A1(new_n857), .A2(new_n750), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n276), .B1(new_n711), .B2(G87), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n212), .B2(new_n707), .C1(new_n718), .C2(new_n203), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n779), .A2(G116), .B1(new_n956), .B2(new_n720), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n796), .B2(new_n705), .C1(new_n207), .C2(new_n727), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1036), .B(new_n1038), .C1(G294), .C2(new_n722), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT121), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n707), .A2(new_n964), .ZN(new_n1043));
  INV_X1    g0843(.A(G128), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n276), .B1(new_n705), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(G132), .C2(new_n779), .ZN(new_n1046));
  XOR2_X1   g0846(.A(KEYINPUT54), .B(G143), .Z(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT120), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1048), .A2(new_n720), .B1(new_n717), .B2(G50), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT53), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n741), .B2(new_n258), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n711), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1051), .A2(new_n1052), .B1(G125), .B2(new_n722), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n734), .A2(G137), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1046), .A2(new_n1049), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1041), .A2(new_n1042), .A3(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(new_n702), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n701), .B1(new_n256), .B2(new_n777), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT119), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1034), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n880), .A2(new_n886), .A3(G330), .A4(new_n772), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n859), .B1(new_n863), .B2(new_n870), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n849), .A2(new_n851), .A3(new_n856), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n654), .A2(new_n772), .A3(new_n630), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n862), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n860), .B1(new_n1067), .B2(new_n880), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n879), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1062), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n690), .A2(G330), .A3(new_n772), .A4(new_n880), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1068), .B2(new_n879), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1064), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1064), .A2(KEYINPUT116), .A3(new_n1073), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1070), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1061), .B1(new_n1078), .B2(new_n697), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT117), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT31), .B1(new_n680), .B2(new_n624), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n686), .A2(new_n689), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n772), .B(G330), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1066), .B(new_n1065), .C1(new_n1083), .C2(new_n870), .ZN(new_n1084));
  INV_X1    g0884(.A(G330), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n584), .A2(new_n630), .B1(new_n680), .B2(new_n688), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n683), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n880), .B1(new_n1087), .B2(new_n772), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1080), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1067), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n886), .A2(G330), .A3(new_n772), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n870), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1090), .A2(new_n1092), .A3(KEYINPUT117), .A4(new_n1071), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1083), .A2(new_n870), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1062), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n863), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1089), .A2(new_n1093), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1087), .A2(new_n429), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n874), .A2(new_n1100), .A3(new_n875), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(KEYINPUT118), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n640), .B1(new_n1078), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1062), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT116), .B1(new_n1064), .B2(new_n1073), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1064), .A2(KEYINPUT116), .A3(new_n1073), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1103), .B(new_n1107), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1079), .B1(new_n1104), .B2(new_n1111), .ZN(G378));
  INV_X1    g0912(.A(new_n847), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n845), .A2(KEYINPUT106), .A3(new_n846), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n854), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n892), .B(G330), .C1(new_n1115), .C2(new_n887), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n427), .B1(new_n587), .B2(new_n588), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1120), .A2(new_n1121), .B1(new_n274), .B2(new_n622), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n274), .A2(new_n622), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1116), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1128), .A2(new_n889), .A3(G330), .A4(new_n892), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n873), .A2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n861), .A2(new_n872), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n697), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n779), .A2(G107), .B1(new_n490), .B2(new_n720), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n729), .A2(G116), .B1(G68), .B2(new_n730), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n206), .C2(new_n727), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n718), .A2(new_n202), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(G41), .B1(new_n711), .B2(G77), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n328), .A3(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1136), .B(new_n1140), .C1(G283), .C2(new_n722), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(KEYINPUT58), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(KEYINPUT58), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G41), .B1(new_n335), .B2(G33), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1143), .C1(G50), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n734), .A2(G132), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n729), .A2(G125), .B1(G150), .B2(new_n730), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n779), .A2(G128), .B1(G137), .B2(new_n720), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1048), .A2(new_n711), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1150), .A2(KEYINPUT59), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(KEYINPUT59), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n311), .B(new_n451), .C1(new_n718), .C2(new_n964), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G124), .B2(new_n722), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n702), .B1(new_n1145), .B2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT122), .Z(new_n1157));
  AOI21_X1  g0957(.A(new_n701), .B1(new_n201), .B2(new_n777), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n1128), .C2(new_n750), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1133), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1101), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1078), .B2(new_n1098), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT57), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n640), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1107), .B(new_n1098), .C1(new_n1109), .C2(new_n1108), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1101), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n873), .B(new_n1130), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1161), .B1(new_n1165), .B2(new_n1169), .ZN(G375));
  NAND2_X1  g0970(.A1(new_n1098), .A2(new_n697), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n870), .A2(new_n749), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n328), .B1(new_n711), .B2(G159), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1138), .B(new_n1173), .C1(new_n1044), .C2(new_n789), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G132), .A2(new_n729), .B1(new_n779), .B2(G137), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n734), .A2(new_n1048), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G50), .A2(new_n730), .B1(new_n720), .B2(G150), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n779), .A2(G283), .B1(G107), .B2(new_n720), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n792), .B2(new_n705), .C1(new_n433), .C2(new_n727), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n722), .A2(G303), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n982), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n276), .B1(new_n711), .B2(G97), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1181), .A2(new_n961), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1174), .A2(new_n1178), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n703), .B1(new_n1185), .B2(KEYINPUT123), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(KEYINPUT123), .B2(new_n1185), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n777), .A2(new_n203), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1172), .A2(new_n698), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1171), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT124), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1171), .A2(KEYINPUT124), .A3(new_n1189), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n925), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1102), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT125), .ZN(G381));
  OR2_X1    g0999(.A1(G393), .A2(G396), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(G381), .A2(G384), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1107), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1202), .A2(new_n696), .B1(new_n1034), .B2(new_n1060), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1103), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n641), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n1110), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(G375), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1010), .A2(new_n1032), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n948), .A3(new_n969), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1201), .A2(new_n1206), .A3(new_n1207), .A4(new_n1210), .ZN(G407));
  NAND2_X1  g1011(.A1(new_n623), .A2(G213), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1207), .A2(new_n1206), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT126), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G213), .B(G407), .C1(new_n1216), .C2(new_n1217), .ZN(G409));
  NAND2_X1  g1018(.A1(new_n1195), .A2(KEYINPUT60), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT60), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n640), .A3(new_n1221), .A4(new_n1102), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1194), .A2(G384), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(G384), .B1(new_n1194), .B2(new_n1222), .ZN(new_n1225));
  INV_X1    g1025(.A(G2897), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1224), .A2(new_n1225), .B1(new_n1226), .B2(new_n1212), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1225), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1212), .A2(new_n1226), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1223), .A3(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1227), .A2(new_n1230), .A3(KEYINPUT127), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT127), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G378), .B(new_n1161), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1167), .A2(new_n1168), .A3(new_n1196), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1206), .B1(new_n1235), .B2(new_n1160), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1212), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1238), .B2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(G396), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1208), .B1(new_n948), .B2(new_n969), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1210), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G387), .A2(G390), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1209), .A3(new_n1244), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(KEYINPUT61), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1213), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1241), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1239), .A2(new_n1243), .A3(new_n1251), .A4(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1252), .A2(new_n1255), .A3(new_n1241), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1252), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1255), .B1(new_n1252), .B2(new_n1241), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1256), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1254), .B1(new_n1261), .B2(new_n1262), .ZN(G405));
  NAND2_X1  g1063(.A1(G375), .A2(new_n1206), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1234), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1250), .A2(new_n1234), .A3(new_n1264), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1242), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1241), .A3(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G402));
endmodule


