//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(KEYINPUT74), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(G125), .A3(G140), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n193), .A3(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT75), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AOI211_X1 g015(.A(KEYINPUT75), .B(new_n192), .C1(new_n195), .C2(new_n197), .ZN(new_n202));
  OAI21_X1  g016(.A(G146), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n204), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT68), .A2(G128), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(KEYINPUT68), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT68), .A2(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n206), .B1(new_n215), .B2(G119), .ZN(new_n216));
  XOR2_X1   g030(.A(KEYINPUT24), .B(G110), .Z(new_n217));
  OAI22_X1  g031(.A1(new_n212), .A2(G110), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n193), .A2(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n194), .A2(G140), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G125), .B(G140), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT76), .A3(new_n221), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n203), .A2(new_n218), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n212), .A2(G110), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n216), .A2(new_n217), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n196), .A2(G125), .A3(G140), .ZN(new_n232));
  AOI21_X1  g046(.A(G140), .B1(new_n196), .B2(G125), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT16), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n200), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n198), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n221), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n231), .B1(new_n239), .B2(new_n203), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n191), .B1(new_n228), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n203), .A2(new_n239), .ZN(new_n243));
  INV_X1    g057(.A(new_n231), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n203), .A2(new_n218), .A3(new_n227), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n190), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n241), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT77), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G234), .ZN(new_n254));
  OAI21_X1  g068(.A(G217), .B1(new_n254), .B2(G902), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(KEYINPUT73), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(KEYINPUT78), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT25), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT78), .B1(new_n248), .B2(new_n249), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n253), .B(new_n256), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n256), .A2(G902), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n241), .A2(new_n247), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n260), .A2(KEYINPUT80), .A3(new_n266), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT11), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(G137), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT11), .A3(G134), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n275), .A2(new_n277), .A3(new_n281), .A4(new_n278), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(G131), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G131), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n275), .A2(new_n277), .A3(new_n284), .A4(new_n278), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  INV_X1    g102(.A(G143), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(G146), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n221), .A2(KEYINPUT65), .A3(G143), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(G146), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT64), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n294), .B(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n221), .A2(G143), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n292), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n293), .A2(new_n295), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n280), .A2(new_n302), .A3(G131), .A4(new_n282), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n290), .A2(new_n291), .A3(new_n305), .A4(new_n292), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n209), .A2(new_n210), .B1(new_n299), .B2(KEYINPUT1), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n299), .A2(new_n292), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n278), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n274), .A2(G137), .ZN(new_n311));
  OAI21_X1  g125(.A(G131), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n285), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n304), .A2(KEYINPUT30), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n304), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n313), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT30), .B1(new_n304), .B2(new_n313), .ZN(new_n319));
  XOR2_X1   g133(.A(G116), .B(G119), .Z(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT2), .B(G113), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT2), .B(G113), .Z(new_n323));
  XNOR2_X1  g137(.A(G116), .B(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n318), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n326), .B(KEYINPUT70), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n304), .A2(new_n330), .A3(new_n313), .ZN(new_n331));
  NOR2_X1   g145(.A1(G237), .A2(G953), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G210), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT27), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G101), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n272), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g153(.A(KEYINPUT31), .B(new_n337), .C1(new_n318), .C2(new_n328), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n304), .A2(new_n313), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n326), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n304), .A2(new_n330), .A3(KEYINPUT28), .A4(new_n313), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n331), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n336), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n339), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT71), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n327), .B(new_n319), .C1(new_n316), .C2(new_n317), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT31), .B1(new_n353), .B2(new_n337), .ZN(new_n354));
  INV_X1    g168(.A(new_n347), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n329), .A2(new_n272), .A3(new_n338), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT71), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n349), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n339), .A2(new_n340), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n350), .B1(new_n361), .B2(new_n355), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n346), .A2(new_n363), .A3(new_n342), .A4(new_n343), .ZN(new_n364));
  INV_X1    g178(.A(new_n330), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n341), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n345), .B1(new_n366), .B2(new_n331), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT72), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n331), .A2(new_n368), .A3(new_n345), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n331), .B2(new_n345), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n336), .B(new_n364), .C1(new_n371), .C2(new_n363), .ZN(new_n372));
  INV_X1    g186(.A(new_n336), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n329), .A2(new_n363), .A3(new_n373), .A4(new_n331), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n242), .A3(new_n374), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n362), .A2(KEYINPUT32), .B1(new_n375), .B2(G472), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n271), .B1(new_n360), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G478), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT15), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT9), .B(G234), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G217), .A3(new_n188), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n209), .A2(G143), .A3(new_n210), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n204), .A2(G143), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n274), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G116), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G122), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n388), .A3(G122), .ZN(new_n391));
  INV_X1    g205(.A(G122), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT91), .B1(new_n392), .B2(G116), .ZN(new_n393));
  AOI211_X1 g207(.A(G107), .B(new_n389), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n391), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(G116), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n387), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n213), .A2(new_n214), .A3(new_n289), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT13), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n204), .B2(G143), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n289), .A2(KEYINPUT13), .A3(G128), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n400), .B(G134), .C1(new_n401), .C2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G134), .B1(new_n401), .B2(new_n405), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT92), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n399), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n397), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n395), .B1(new_n397), .B2(KEYINPUT14), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n396), .B(new_n397), .C1(KEYINPUT14), .C2(new_n395), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n384), .A2(new_n274), .A3(new_n386), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n274), .B1(new_n384), .B2(new_n386), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G134), .B1(new_n401), .B2(new_n385), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(KEYINPUT93), .A3(new_n387), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n414), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n383), .B1(new_n409), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n412), .A2(new_n413), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n416), .A2(new_n417), .A3(new_n415), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT93), .B1(new_n419), .B2(new_n387), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n408), .A2(new_n406), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n410), .A2(G107), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n389), .B1(new_n393), .B2(new_n391), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n395), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n416), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n383), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n426), .A2(new_n432), .A3(KEYINPUT94), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n422), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n418), .A2(new_n420), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n436), .A2(new_n423), .B1(new_n427), .B2(new_n431), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT94), .B1(new_n437), .B2(new_n433), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n242), .B(new_n380), .C1(new_n435), .C2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n426), .A2(new_n432), .A3(new_n433), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT94), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n422), .A3(new_n434), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n380), .B1(new_n444), .B2(new_n242), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT90), .B(G475), .Z(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n188), .A3(G214), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n289), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n332), .A2(G143), .A3(G214), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n284), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT17), .ZN(new_n455));
  AND4_X1   g269(.A1(G143), .A2(new_n450), .A3(new_n188), .A4(G214), .ZN(new_n456));
  AOI21_X1  g270(.A(G143), .B1(new_n332), .B2(G214), .ZN(new_n457));
  OAI21_X1  g271(.A(G131), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(new_n284), .A3(new_n453), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n203), .A2(new_n239), .A3(new_n455), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n452), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n195), .A2(G146), .A3(new_n197), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT76), .B1(new_n225), .B2(new_n221), .ZN(new_n468));
  AND4_X1   g282(.A1(KEYINPUT76), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n456), .A2(new_n457), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT88), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n473));
  NOR4_X1   g287(.A1(new_n456), .A2(new_n457), .A3(new_n473), .A4(new_n465), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n466), .B(new_n470), .C1(new_n472), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  INV_X1    g291(.A(G104), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n462), .A2(new_n479), .A3(new_n475), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n449), .B1(new_n483), .B2(new_n242), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(G475), .A2(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n452), .A2(new_n453), .A3(new_n464), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT88), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n470), .A2(new_n466), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n221), .B1(new_n236), .B2(new_n238), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n195), .A2(KEYINPUT19), .A3(new_n197), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT19), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n219), .A2(new_n220), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n221), .A3(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n456), .A2(new_n457), .A3(G131), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n454), .ZN(new_n497));
  OAI22_X1  g311(.A1(new_n489), .A2(new_n490), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n492), .A2(new_n494), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n501), .A2(new_n221), .B1(new_n458), .B2(new_n460), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n203), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n475), .A3(KEYINPUT89), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n480), .A3(new_n504), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT20), .B(new_n487), .C1(new_n505), .C2(new_n482), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n480), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT89), .B1(new_n503), .B2(new_n475), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n482), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n510), .B2(new_n486), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n485), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n447), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G214), .B1(G237), .B2(G902), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT85), .ZN(new_n515));
  OAI21_X1  g329(.A(G210), .B1(G237), .B2(G902), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G224), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT7), .B1(new_n518), .B2(G953), .ZN(new_n519));
  INV_X1    g333(.A(new_n301), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G125), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n194), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT87), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(KEYINPUT87), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT3), .B1(new_n478), .B2(G107), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT3), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n395), .A3(G104), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n478), .A2(G107), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G101), .ZN(new_n532));
  INV_X1    g346(.A(G101), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n527), .A2(new_n529), .A3(new_n533), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(KEYINPUT4), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n536), .A3(G101), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n326), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n478), .A2(G107), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n395), .A2(G104), .ZN(new_n540));
  OAI21_X1  g354(.A(G101), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n543));
  OR3_X1    g357(.A1(new_n388), .A2(KEYINPUT5), .A3(G119), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(G113), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n325), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G122), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n538), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n522), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n520), .B2(G125), .ZN(new_n550));
  INV_X1    g364(.A(new_n519), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n547), .B(KEYINPUT8), .ZN(new_n553));
  INV_X1    g367(.A(new_n546), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n542), .B1(new_n325), .B2(new_n545), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n526), .A2(new_n548), .A3(new_n552), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n242), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n518), .A2(G953), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n550), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n548), .A2(KEYINPUT6), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n538), .A2(new_n546), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n547), .A2(KEYINPUT86), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(KEYINPUT6), .A3(new_n563), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n517), .B1(new_n558), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n560), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n571), .A2(new_n242), .A3(new_n516), .A4(new_n557), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n515), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(G234), .A2(G237), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(G952), .A3(new_n188), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(G902), .A3(G953), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT21), .B(G898), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT10), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n204), .B1(new_n299), .B2(KEYINPUT1), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n306), .B1(new_n293), .B2(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n585), .A2(new_n542), .A3(KEYINPUT81), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT81), .B1(new_n585), .B2(new_n542), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n535), .A2(new_n301), .A3(new_n537), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n542), .A2(new_n309), .A3(KEYINPUT10), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n287), .A2(new_n303), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G140), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n188), .A2(G227), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT84), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT12), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n542), .A2(new_n309), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n585), .A2(new_n542), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n585), .A2(new_n542), .A3(KEYINPUT81), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n600), .B1(new_n606), .B2(new_n592), .ZN(new_n607));
  INV_X1    g421(.A(new_n592), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n586), .A2(new_n587), .ZN(new_n609));
  OAI211_X1 g423(.A(KEYINPUT12), .B(new_n608), .C1(new_n609), .C2(new_n601), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT84), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n593), .A2(new_n612), .A3(new_n597), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n599), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT10), .B1(new_n604), .B2(new_n605), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n589), .A2(new_n590), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n608), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n597), .B1(new_n617), .B2(new_n593), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT83), .B(G469), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n242), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n597), .B1(new_n611), .B2(new_n593), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n617), .A2(new_n593), .A3(new_n597), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT82), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT82), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n615), .A2(new_n608), .A3(new_n616), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n610), .B2(new_n607), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n625), .B(new_n628), .C1(new_n630), .C2(new_n597), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G469), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n623), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(G221), .B1(new_n381), .B2(G902), .ZN(new_n635));
  AND4_X1   g449(.A1(new_n513), .A2(new_n582), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n377), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G101), .ZN(G3));
  INV_X1    g452(.A(G472), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n357), .B2(new_n242), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n641), .A2(new_n351), .A3(new_n359), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n271), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n634), .A2(new_n635), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n582), .ZN(new_n647));
  INV_X1    g461(.A(new_n482), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n488), .B(new_n473), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n227), .A2(new_n467), .B1(new_n463), .B2(new_n465), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n649), .A2(new_n650), .B1(new_n502), .B2(new_n203), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n479), .B1(new_n651), .B2(KEYINPUT89), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n648), .B1(new_n652), .B2(new_n500), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT20), .B1(new_n653), .B2(new_n487), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n510), .A2(new_n507), .A3(new_n486), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n484), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n422), .A2(KEYINPUT33), .A3(new_n441), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n378), .A2(G902), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT95), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n659), .B(new_n660), .C1(new_n435), .C2(new_n438), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n659), .B1(new_n444), .B2(new_n660), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n657), .B(new_n658), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n242), .B1(new_n435), .B2(new_n438), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n378), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n656), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT96), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT96), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n647), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n644), .A2(new_n646), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT34), .B(G104), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G6));
  NAND2_X1  g487(.A1(new_n447), .A2(new_n656), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n647), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n644), .A2(new_n646), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n228), .A2(new_n240), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT97), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n261), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n260), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n636), .A2(new_n642), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT98), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G12));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n360), .A2(new_n376), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n579), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n576), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n440), .B2(new_n445), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT100), .B1(new_n696), .B2(new_n512), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n665), .A2(new_n379), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n698), .A2(new_n439), .B1(new_n576), .B2(new_n694), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n656), .A3(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n697), .A2(new_n573), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n635), .A3(new_n634), .A4(new_n684), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n689), .B1(new_n690), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n360), .A2(new_n376), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n634), .A2(new_n635), .A3(new_n684), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT101), .A4(new_n702), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  NAND3_X1  g523(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n329), .A2(new_n331), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n336), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n366), .A2(new_n331), .ZN(new_n713));
  AOI21_X1  g527(.A(G902), .B1(new_n713), .B2(new_n373), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G472), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n360), .A2(new_n710), .A3(new_n716), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n695), .B(KEYINPUT39), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n646), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n722), .A2(KEYINPUT40), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n568), .A2(new_n572), .ZN(new_n725));
  XOR2_X1   g539(.A(new_n725), .B(KEYINPUT38), .Z(new_n726));
  INV_X1    g540(.A(new_n259), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT25), .A3(new_n257), .ZN(new_n728));
  INV_X1    g542(.A(new_n256), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n259), .B2(new_n252), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n261), .A2(new_n682), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n515), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n656), .A2(new_n446), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n720), .A2(new_n723), .A3(new_n724), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  NAND2_X1  g551(.A1(new_n664), .A2(new_n666), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n512), .A3(new_n573), .A4(new_n695), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n667), .A2(KEYINPUT103), .A3(new_n573), .A4(new_n695), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n705), .A3(new_n706), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT104), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n743), .A2(new_n705), .A3(new_n706), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G146), .ZN(G48));
  INV_X1    g563(.A(new_n635), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n598), .A2(KEYINPUT84), .B1(new_n607), .B2(new_n610), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n618), .B1(new_n751), .B2(new_n613), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n752), .B2(G902), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n623), .A3(KEYINPUT105), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(G469), .C1(new_n752), .C2(G902), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n750), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n670), .A2(new_n377), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT41), .B(G113), .Z(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT106), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n758), .B(new_n760), .ZN(G15));
  NAND3_X1  g575(.A1(new_n377), .A2(new_n675), .A3(new_n757), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G116), .ZN(G18));
  NAND2_X1  g577(.A1(new_n684), .A2(new_n513), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n360), .B2(new_n376), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n582), .A3(new_n757), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  OR2_X1    g581(.A1(new_n371), .A2(new_n336), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n350), .B1(new_n361), .B2(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n640), .A2(new_n769), .A3(new_n267), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(new_n757), .A3(new_n582), .A4(new_n733), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  NOR2_X1   g586(.A1(new_n640), .A2(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n684), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT107), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT107), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n776), .A3(new_n684), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n738), .A2(new_n512), .A3(new_n695), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n667), .A2(new_n781), .A3(new_n695), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n754), .A2(new_n756), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n635), .A3(new_n573), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  NOR3_X1   g602(.A1(new_n752), .A2(G902), .A3(new_n621), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n625), .B1(new_n630), .B2(new_n597), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n633), .B1(new_n790), .B2(new_n242), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT109), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n790), .A2(new_n242), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n623), .B(new_n793), .C1(new_n794), .C2(new_n633), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n568), .A2(new_n572), .A3(new_n732), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n750), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n780), .A2(new_n796), .A3(new_n782), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n267), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n375), .A2(G472), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n710), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT42), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n667), .A2(new_n781), .A3(new_n695), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n781), .B1(new_n667), .B2(new_n695), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT42), .ZN(new_n809));
  INV_X1    g623(.A(new_n798), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n795), .B2(new_n792), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n377), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n805), .A2(new_n812), .A3(KEYINPUT110), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT110), .B1(new_n805), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G131), .ZN(G33));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n697), .A2(new_n701), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n697), .A2(new_n701), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT111), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n377), .A2(new_n811), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G134), .ZN(G36));
  INV_X1    g636(.A(new_n721), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n633), .A2(new_n242), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT45), .B1(new_n627), .B2(new_n631), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n827));
  OAI21_X1  g641(.A(G469), .B1(new_n790), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(KEYINPUT46), .B(new_n825), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(KEYINPUT112), .A3(new_n623), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n826), .A2(new_n828), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n824), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(KEYINPUT46), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT112), .B1(new_n829), .B2(new_n623), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n635), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n738), .A2(new_n656), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT43), .B1(new_n656), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n738), .B(new_n656), .C1(new_n837), .C2(KEYINPUT43), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT114), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT114), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n643), .A3(new_n684), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT44), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n823), .B(new_n835), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n797), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(KEYINPUT115), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(KEYINPUT115), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G137), .ZN(G39));
  INV_X1    g666(.A(KEYINPUT47), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n835), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n835), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n271), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n705), .A2(new_n857), .A3(new_n779), .A4(new_n797), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(G140), .ZN(G42));
  AND3_X1   g674(.A1(new_n754), .A2(KEYINPUT49), .A3(new_n756), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT49), .B1(new_n754), .B2(new_n756), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n267), .A2(new_n750), .A3(new_n515), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n726), .A2(new_n656), .A3(new_n863), .A4(new_n738), .ZN(new_n864));
  OR4_X1    g678(.A1(new_n720), .A2(new_n861), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n640), .A2(new_n731), .A3(new_n769), .A4(KEYINPUT107), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n776), .B1(new_n773), .B2(new_n684), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n808), .B(new_n811), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n656), .A2(new_n446), .A3(new_n695), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT117), .B1(new_n869), .B2(new_n797), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n869), .A2(KEYINPUT117), .A3(new_n797), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n705), .A2(new_n706), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n821), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n805), .A2(new_n812), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT110), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n805), .A2(new_n812), .A3(KEYINPUT110), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n645), .A2(new_n647), .ZN(new_n879));
  INV_X1    g693(.A(new_n667), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n674), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n857), .A3(new_n642), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n685), .A3(new_n637), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n874), .A2(new_n877), .A3(new_n878), .A4(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n758), .A2(new_n762), .A3(new_n766), .A4(new_n771), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n770), .A2(new_n733), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n582), .B(new_n757), .C1(new_n888), .C2(new_n765), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n890), .A3(new_n758), .A4(new_n762), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n704), .A2(new_n707), .B1(new_n778), .B2(new_n786), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n733), .A2(new_n732), .A3(new_n725), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n695), .A2(new_n635), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n684), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n717), .A2(new_n796), .A3(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n894), .A2(new_n748), .A3(new_n895), .A4(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n748), .A3(new_n899), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT52), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n894), .B2(new_n895), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n893), .A2(new_n900), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n900), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n873), .A2(new_n883), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n815), .A2(new_n887), .A3(new_n891), .A4(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT54), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n576), .B1(new_n839), .B2(new_n840), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n770), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT50), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n757), .A2(new_n515), .A3(new_n726), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n757), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(new_n797), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n778), .A2(new_n912), .A3(new_n920), .ZN(new_n921));
  NOR4_X1   g735(.A1(new_n919), .A2(new_n271), .A3(new_n576), .A4(new_n797), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n738), .A2(new_n512), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n718), .A3(new_n719), .A4(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n784), .A2(new_n750), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n854), .A2(new_n855), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n913), .A2(new_n797), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT118), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n913), .A2(new_n785), .ZN(new_n931));
  INV_X1    g745(.A(G952), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(G953), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n668), .A2(new_n669), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n922), .A2(new_n718), .A3(new_n934), .A4(new_n719), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n804), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n920), .A2(new_n937), .A3(new_n912), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT48), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT48), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n920), .A2(new_n937), .A3(new_n940), .A4(new_n912), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n930), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n930), .A2(new_n942), .A3(new_n935), .A4(new_n933), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n929), .A2(KEYINPUT51), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n925), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n927), .A2(new_n928), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT51), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT119), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT54), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n894), .A2(new_n895), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n886), .ZN(new_n954));
  NOR4_X1   g768(.A1(new_n873), .A2(new_n875), .A3(new_n883), .A4(new_n903), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n954), .A2(new_n955), .A3(new_n902), .A4(new_n900), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n909), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n948), .A2(new_n949), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n929), .A2(KEYINPUT51), .ZN(new_n959));
  INV_X1    g773(.A(new_n944), .ZN(new_n960));
  INV_X1    g774(.A(new_n942), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n933), .A2(new_n935), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT118), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT119), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n958), .A2(new_n959), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n911), .A2(new_n951), .A3(new_n957), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(G952), .A2(G953), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n865), .B1(new_n967), .B2(new_n968), .ZN(G75));
  NOR2_X1   g783(.A1(new_n188), .A2(G952), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n909), .A2(new_n956), .ZN(new_n971));
  NAND2_X1  g785(.A1(G210), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n570), .B(new_n560), .ZN(new_n973));
  XOR2_X1   g787(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT121), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI22_X1  g792(.A1(new_n971), .A2(new_n972), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT56), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n909), .A2(new_n956), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(new_n976), .A3(G210), .A4(G902), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n971), .A2(new_n972), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n977), .A2(new_n980), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n975), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n970), .B1(new_n983), .B2(new_n986), .ZN(G51));
  AND4_X1   g801(.A1(KEYINPUT124), .A2(new_n981), .A3(G902), .A4(new_n831), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n242), .B1(new_n909), .B2(new_n956), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT124), .B1(new_n989), .B2(new_n831), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n824), .B(KEYINPUT123), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT57), .Z(new_n993));
  AND3_X1   g807(.A1(new_n909), .A2(new_n952), .A3(new_n956), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n952), .B1(new_n909), .B2(new_n956), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n620), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n970), .B1(new_n991), .B2(new_n997), .ZN(G54));
  AND2_X1   g812(.A1(KEYINPUT58), .A2(G475), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n989), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n970), .B1(new_n1000), .B2(new_n653), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n989), .A2(new_n1002), .A3(new_n510), .A4(new_n999), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n989), .A2(new_n510), .A3(new_n999), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT125), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(G60));
  INV_X1    g820(.A(new_n657), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n660), .B1(new_n435), .B2(new_n438), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(KEYINPUT95), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1007), .B1(new_n1009), .B2(new_n661), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n911), .A2(new_n957), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G478), .A2(G902), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT59), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1010), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n994), .B2(new_n995), .ZN(new_n1016));
  INV_X1    g830(.A(new_n970), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1014), .A2(new_n1018), .ZN(G63));
  INV_X1    g833(.A(KEYINPUT61), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G217), .A2(G902), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT60), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n909), .B2(new_n956), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n682), .B(KEYINPUT126), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  OR2_X1    g840(.A1(new_n264), .A2(new_n265), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1017), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1020), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  OR2_X1    g843(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1030), .A2(KEYINPUT61), .A3(new_n1017), .A4(new_n1025), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1031), .ZN(G66));
  INV_X1    g846(.A(new_n580), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n188), .B1(new_n1033), .B2(G224), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n887), .A2(new_n891), .A3(new_n884), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(new_n188), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n565), .B(new_n566), .C1(G898), .C2(new_n188), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1036), .B(new_n1037), .Z(G69));
  AOI21_X1  g852(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(KEYINPUT127), .ZN(new_n1040));
  OR2_X1    g854(.A1(new_n1039), .A2(KEYINPUT127), .ZN(new_n1041));
  OR4_X1    g855(.A1(new_n823), .A2(new_n835), .A3(new_n804), .A4(new_n896), .ZN(new_n1042));
  AND4_X1   g856(.A1(new_n748), .A2(new_n1042), .A3(new_n821), .A4(new_n894), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n859), .A2(new_n815), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1043), .A2(new_n1044), .A3(new_n188), .A4(new_n851), .ZN(new_n1045));
  INV_X1    g859(.A(new_n341), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n318), .B1(KEYINPUT30), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(new_n501), .Z(new_n1048));
  INV_X1    g862(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1049), .B1(G900), .B2(G953), .ZN(new_n1050));
  AND2_X1   g864(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n736), .A2(new_n748), .A3(new_n894), .ZN(new_n1052));
  OR2_X1    g866(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1053));
  AOI211_X1 g867(.A(new_n797), .B(new_n722), .C1(new_n880), .C2(new_n674), .ZN(new_n1054));
  AOI22_X1  g868(.A1(new_n856), .A2(new_n858), .B1(new_n377), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1056));
  NAND4_X1  g870(.A1(new_n851), .A2(new_n1053), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1048), .B1(new_n1057), .B2(new_n188), .ZN(new_n1058));
  OAI211_X1 g872(.A(new_n1040), .B(new_n1041), .C1(new_n1051), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1057), .A2(new_n188), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(new_n1049), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1062));
  NAND4_X1  g876(.A1(new_n1061), .A2(KEYINPUT127), .A3(new_n1062), .A4(new_n1039), .ZN(new_n1063));
  AND2_X1   g877(.A1(new_n1059), .A2(new_n1063), .ZN(G72));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  OAI21_X1  g880(.A(new_n1066), .B1(new_n1057), .B2(new_n1035), .ZN(new_n1067));
  INV_X1    g881(.A(new_n712), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n970), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1043), .A2(new_n1044), .A3(new_n851), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1066), .B1(new_n1070), .B2(new_n1035), .ZN(new_n1071));
  NOR2_X1   g885(.A1(new_n711), .A2(new_n336), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g887(.A(new_n1066), .ZN(new_n1074));
  NOR3_X1   g888(.A1(new_n1068), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n910), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g890(.A1(new_n1069), .A2(new_n1073), .A3(new_n1076), .ZN(G57));
endmodule


