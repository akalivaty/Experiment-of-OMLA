//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT66), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n470), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n470), .A2(new_n462), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT67), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n478), .B(new_n481), .C1(new_n483), .C2(G124), .ZN(G162));
  NAND2_X1  g059(.A1(new_n461), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G126), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n462), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(KEYINPUT69), .C1(new_n469), .C2(new_n468), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n462), .A2(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT69), .A3(KEYINPUT4), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n470), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n461), .B2(new_n492), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n490), .A2(new_n495), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n506), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n508), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n515), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n507), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT70), .B(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n514), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n521), .B1(new_n522), .B2(new_n523), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n507), .A2(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n514), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n517), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(new_n507), .A2(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n539), .B2(new_n514), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n517), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT72), .Z(G188));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  AND2_X1   g125(.A1(KEYINPUT5), .A2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(KEYINPUT5), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G65), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n550), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n553), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT73), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n561), .A2(KEYINPUT74), .A3(G651), .A4(new_n556), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n507), .B2(G53), .ZN(new_n565));
  AND2_X1   g140(.A1(KEYINPUT6), .A2(G651), .ZN(new_n566));
  NOR2_X1   g141(.A1(KEYINPUT6), .A2(G651), .ZN(new_n567));
  OAI211_X1 g142(.A(G53), .B(G543), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n565), .A2(new_n569), .B1(new_n570), .B2(new_n514), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n563), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(new_n514), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n507), .A2(G49), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n507), .A2(G48), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n514), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n512), .B2(G61), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n517), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n517), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n522), .A2(new_n592), .B1(new_n514), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n596));
  OAI221_X1 g171(.A(new_n596), .B1(new_n514), .B2(new_n593), .C1(new_n592), .C2(new_n522), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n591), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n576), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n514), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n512), .A2(G66), .ZN(new_n606));
  INV_X1    g181(.A(G79), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n504), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n600), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n600), .B1(new_n610), .B2(G868), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n571), .B1(new_n559), .B2(new_n562), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(G868), .B2(new_n614), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g197(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G123), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n476), .A2(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n462), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n627), .B1(new_n632), .B2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n626), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G2096), .C2(new_n632), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT76), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n648), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT77), .ZN(G401));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n626), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(G2096), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n668), .B2(new_n673), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n671), .A2(KEYINPUT78), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(KEYINPUT78), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n668), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT79), .B(KEYINPUT20), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n675), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  XNOR2_X1  g263(.A(KEYINPUT31), .B(G11), .ZN(new_n689));
  INV_X1    g264(.A(G28), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(KEYINPUT30), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT30), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(G28), .ZN(new_n694));
  OAI221_X1 g269(.A(new_n689), .B1(new_n691), .B2(new_n694), .C1(new_n632), .C2(new_n692), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G19), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n543), .B2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(G1341), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n483), .A2(G129), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n476), .A2(G141), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT26), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n699), .A2(new_n700), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  INV_X1    g280(.A(G32), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(G29), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT27), .B(G1996), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n692), .A2(G27), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G164), .B2(new_n692), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n707), .A2(new_n709), .B1(G2078), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n698), .B(new_n712), .C1(G2078), .C2(new_n711), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n692), .A2(G35), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT89), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n692), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT29), .B(G2090), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G5), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G171), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n718), .B(new_n723), .C1(G1341), .C2(new_n697), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n692), .A2(G26), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT85), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n483), .A2(G128), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n729));
  INV_X1    g304(.A(G116), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G2105), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n476), .B2(G140), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT86), .B(G2067), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n719), .A2(G4), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n610), .B2(new_n719), .ZN(new_n738));
  INV_X1    g313(.A(G1348), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n692), .B1(KEYINPUT24), .B2(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(KEYINPUT24), .B2(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n474), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n719), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n719), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G1966), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n736), .A2(new_n740), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n713), .A2(new_n724), .A3(new_n749), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n705), .B(new_n708), .C1(G29), .C2(new_n706), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n692), .A2(G33), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n461), .A2(G127), .ZN(new_n753));
  NAND2_X1  g328(.A1(G115), .A2(G2104), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(G2105), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT25), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n476), .A2(G139), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n752), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2072), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n751), .B(new_n764), .C1(new_n744), .C2(new_n743), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(KEYINPUT87), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n747), .A2(G1966), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT88), .Z(new_n768));
  NOR2_X1   g343(.A1(new_n765), .A2(KEYINPUT87), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n719), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n614), .B2(new_n719), .ZN(new_n773));
  INV_X1    g348(.A(G1956), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n750), .A2(new_n766), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT90), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n719), .A2(G23), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n580), .B2(new_n719), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT83), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT84), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n719), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n719), .ZN(new_n786));
  INV_X1    g361(.A(G1971), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G6), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n588), .B2(G16), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n783), .A2(new_n784), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT82), .B(KEYINPUT34), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n692), .A2(G25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n483), .A2(G119), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n476), .A2(G131), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n462), .A2(G107), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT80), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(G29), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n719), .A2(G24), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n808));
  OAI21_X1  g383(.A(G16), .B1(new_n598), .B2(KEYINPUT81), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G1986), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n795), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT36), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n777), .A2(new_n815), .ZN(G311));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n817));
  XNOR2_X1  g392(.A(G311), .B(new_n817), .ZN(G150));
  NAND2_X1  g393(.A1(new_n610), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n507), .A2(G55), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n514), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n517), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n543), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n543), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n820), .B(new_n829), .Z(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n826), .A2(new_n832), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT93), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT92), .B(KEYINPUT37), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n801), .B(KEYINPUT95), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n624), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT94), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT68), .B1(new_n470), .B2(new_n496), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n497), .A2(KEYINPUT69), .A3(KEYINPUT4), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n461), .A2(new_n492), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n847));
  NAND2_X1  g422(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n496), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(KEYINPUT4), .B1(new_n849), .B2(KEYINPUT69), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n842), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n495), .A2(new_n843), .A3(KEYINPUT94), .A4(new_n845), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n489), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n762), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n841), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n704), .B(new_n733), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n476), .A2(G142), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n462), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n483), .B2(G130), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n856), .B(new_n861), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n855), .B(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n632), .B(new_n474), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G162), .ZN(new_n865));
  AOI21_X1  g440(.A(G37), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n863), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g443(.A(new_n598), .B(G288), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(G290), .A2(G288), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n598), .A2(new_n580), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT99), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G303), .B(new_n588), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n869), .A2(new_n877), .A3(new_n870), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n879), .A2(KEYINPUT100), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n829), .B(new_n619), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n605), .A2(new_n609), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n614), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n883), .B1(new_n614), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n888));
  NAND3_X1  g463(.A1(G299), .A2(new_n888), .A3(new_n610), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT96), .B1(new_n614), .B2(new_n884), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT98), .Z(new_n894));
  INV_X1    g469(.A(new_n882), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n886), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n614), .A2(new_n883), .A3(new_n884), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n894), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n881), .B(new_n902), .Z(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G868), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n826), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n826), .ZN(G331));
  AND3_X1   g481(.A1(new_n876), .A2(KEYINPUT102), .A3(new_n878), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT102), .B1(new_n876), .B2(new_n878), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n910));
  XNOR2_X1  g485(.A(G171), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n829), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G171), .B(KEYINPUT101), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n827), .A3(new_n828), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(G286), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n914), .A3(G168), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n892), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n900), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n897), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n892), .A2(new_n920), .A3(new_n896), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n917), .ZN(new_n927));
  AOI21_X1  g502(.A(G168), .B1(new_n912), .B2(new_n914), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT41), .B1(new_n887), .B2(new_n891), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n920), .B2(new_n900), .ZN(new_n931));
  INV_X1    g506(.A(new_n923), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n925), .B(new_n929), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n909), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n901), .A2(new_n929), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n879), .A3(new_n919), .ZN(new_n937));
  INV_X1    g512(.A(G37), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n919), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n909), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n938), .A3(new_n937), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT104), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n919), .A3(new_n933), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT43), .B(new_n939), .C1(new_n952), .C2(new_n909), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n945), .B1(new_n940), .B2(new_n943), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n948), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n949), .B1(new_n941), .B2(new_n946), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n935), .A2(new_n945), .A3(new_n940), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT44), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT105), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n957), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  INV_X1    g539(.A(G1966), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT94), .B1(new_n501), .B2(new_n495), .ZN(new_n966));
  INV_X1    g541(.A(new_n852), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n490), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT106), .B1(new_n853), .B2(G1384), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT45), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n464), .A2(G40), .A3(new_n473), .A4(new_n465), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n495), .A2(new_n845), .A3(new_n843), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n970), .B1(new_n977), .B2(new_n489), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n965), .B1(new_n973), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n971), .A2(new_n972), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n974), .B1(KEYINPUT50), .B2(new_n978), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n744), .A3(new_n983), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n964), .B(G286), .C1(new_n980), .C2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G2090), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n968), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n974), .B1(new_n976), .B2(new_n978), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n787), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G303), .A2(G8), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT55), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(G8), .A3(new_n995), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n985), .A2(KEYINPUT63), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n580), .A2(G1976), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(G8), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(KEYINPUT52), .ZN(new_n1003));
  INV_X1    g578(.A(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(G288), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1000), .A2(G8), .A3(new_n1001), .A4(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n586), .A2(new_n517), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n576), .A2(G86), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT107), .B(G1981), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1007), .A2(new_n1008), .A3(new_n582), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(G1981), .B1(new_n584), .B2(new_n587), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT108), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1000), .A2(G8), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1006), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n999), .B1(new_n1003), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1002), .A2(KEYINPUT52), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(KEYINPUT109), .A3(new_n1006), .A4(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n995), .B1(new_n992), .B2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n998), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  AOI211_X1 g599(.A(KEYINPUT112), .B(new_n1022), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n997), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g603(.A(KEYINPUT113), .B(new_n997), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n981), .B1(new_n971), .B2(new_n972), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n978), .B2(KEYINPUT50), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n502), .A2(KEYINPUT110), .A3(new_n981), .A4(new_n970), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n974), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1030), .A2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1036), .A2(new_n986), .B1(new_n787), .B2(new_n990), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n994), .B1(new_n1037), .B2(new_n964), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1003), .A2(new_n1017), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n996), .A4(new_n985), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT63), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1040), .A2(KEYINPUT111), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT111), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1028), .A2(new_n1029), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1348), .B1(new_n982), .B2(new_n983), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1000), .A2(G2067), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n610), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n1051), .B2(new_n610), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n610), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT120), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1052), .A3(new_n610), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1049), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n543), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT58), .B(G1341), .Z(new_n1062));
  NAND2_X1  g637(.A1(new_n1000), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1996), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n988), .A2(new_n989), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT59), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n507), .A2(new_n564), .A3(G53), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(KEYINPUT115), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(KEYINPUT115), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n514), .A2(new_n570), .ZN(new_n1074));
  NOR4_X1   g649(.A1(new_n1072), .A2(new_n1073), .A3(KEYINPUT57), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1075), .A2(new_n563), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n774), .C1(new_n1030), .C2(new_n1035), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT116), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n988), .A2(new_n989), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT117), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n988), .A2(new_n989), .A3(new_n1084), .A4(new_n1081), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n853), .A2(KEYINPUT106), .A3(G1384), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT50), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1034), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1078), .B1(new_n1091), .B2(new_n774), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1077), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT114), .B1(new_n1036), .B2(G1956), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1094), .A2(new_n1076), .A3(new_n1079), .A4(new_n1086), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1067), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1095), .A2(KEYINPUT61), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT119), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1094), .A2(new_n1101), .A3(new_n1079), .A4(new_n1086), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1077), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1060), .A2(new_n1098), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n610), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1106));
  XOR2_X1   g681(.A(new_n1106), .B(KEYINPUT118), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1095), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1038), .A2(new_n1039), .A3(new_n996), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n980), .A2(G168), .A3(new_n984), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  AOI21_X1  g689(.A(G168), .B1(new_n980), .B2(new_n984), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1117), .A3(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n990), .A2(G2078), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n973), .A2(new_n979), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(G2078), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n982), .A2(new_n983), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n722), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT45), .B1(new_n968), .B2(new_n970), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n853), .A2(new_n976), .A3(G1384), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n462), .B1(new_n472), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1133), .B2(new_n472), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n466), .A2(G40), .A3(new_n1135), .A4(new_n1125), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1131), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1127), .B2(new_n722), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT122), .B(G1961), .C1(new_n982), .C2(new_n983), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1138), .B(G301), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1130), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1112), .B(new_n1119), .C1(new_n1143), .C2(KEYINPUT54), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n1129), .B2(G171), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT124), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1138), .B(new_n1148), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1145), .B1(new_n1150), .B2(G171), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1144), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1110), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1016), .A2(new_n1004), .A3(new_n580), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1010), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1155), .A2(G8), .A3(new_n1000), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1021), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(new_n996), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1130), .B(new_n1111), .C1(new_n1119), .C2(KEYINPUT62), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1045), .A2(new_n1153), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1131), .A2(new_n975), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n704), .B(new_n1064), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n733), .A2(G2067), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n733), .A2(G2067), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n801), .B(new_n805), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n598), .B(new_n811), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1164), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1164), .A2(new_n1064), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT46), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1167), .A2(new_n1166), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1164), .B1(new_n704), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT125), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT47), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1178), .B(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT47), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1168), .A2(new_n802), .A3(new_n805), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1163), .B1(new_n1185), .B2(new_n1167), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1164), .A2(new_n811), .A3(new_n598), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT126), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT48), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1188), .A2(new_n1189), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1181), .A2(new_n1184), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1193), .B(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1173), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g771(.A1(G227), .A2(new_n459), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n652), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1199), .A2(G229), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n867), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n953), .A2(new_n954), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n1201), .A2(new_n1202), .ZN(G308));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(G225));
endmodule


