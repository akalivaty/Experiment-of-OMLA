//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n201), .B(new_n206), .C1(new_n202), .C2(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n204), .A2(new_n210), .A3(new_n205), .A4(new_n207), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n209), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT69), .B1(new_n209), .B2(new_n211), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n200), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT2), .B(G113), .Z(new_n215));
  XNOR2_X1  g029(.A(G116), .B(G119), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  AOI21_X1  g035(.A(G128), .B1(new_n194), .B2(new_n196), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n195), .A2(KEYINPUT1), .A3(G146), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n223), .B(KEYINPUT68), .C1(new_n190), .C2(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n190), .A2(new_n228), .A3(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n202), .A2(G137), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT67), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n205), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n232), .B(G131), .C1(new_n234), .C2(new_n231), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(new_n235), .A3(new_n211), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n214), .A2(new_n220), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT70), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n214), .A2(new_n239), .A3(new_n220), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n214), .A2(KEYINPUT30), .A3(new_n236), .ZN(new_n242));
  INV_X1    g056(.A(new_n229), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n225), .B2(new_n226), .ZN(new_n244));
  INV_X1    g058(.A(new_n235), .ZN(new_n245));
  INV_X1    g059(.A(new_n211), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI221_X4 g061(.A(KEYINPUT66), .B1(new_n199), .B2(new_n192), .C1(new_n209), .C2(new_n211), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n209), .A2(new_n211), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(new_n200), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n247), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n219), .B(new_n242), .C1(new_n252), .C2(KEYINPUT30), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G210), .ZN(new_n255));
  INV_X1    g069(.A(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n257), .B(new_n258), .Z(new_n259));
  NAND3_X1  g073(.A1(new_n241), .A2(new_n253), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n241), .A2(new_n253), .A3(KEYINPUT31), .A4(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n237), .A2(new_n265), .ZN(new_n266));
  OR3_X1    g080(.A1(new_n247), .A2(new_n248), .A3(new_n251), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n238), .A2(new_n240), .B1(new_n267), .B2(new_n219), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n268), .B2(new_n265), .ZN(new_n269));
  INV_X1    g083(.A(new_n259), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n188), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n273), .ZN(new_n275));
  AOI211_X1 g089(.A(KEYINPUT71), .B(new_n275), .C1(new_n264), .C2(new_n271), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n187), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(KEYINPUT32), .A3(new_n273), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n269), .A2(new_n270), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n241), .A2(new_n253), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n270), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n220), .B1(new_n214), .B2(new_n236), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n238), .B2(new_n240), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n266), .B1(new_n286), .B2(new_n265), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G472), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n278), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G128), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n197), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n229), .A2(new_n294), .A3(new_n223), .ZN(new_n295));
  INV_X1    g109(.A(G107), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G104), .ZN(new_n297));
  INV_X1    g111(.A(G104), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G107), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n256), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(new_n298), .B2(G107), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n296), .A3(G104), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n302), .A2(new_n304), .A3(new_n256), .A4(new_n299), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n295), .B(new_n301), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n296), .A2(G104), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(KEYINPUT3), .B2(new_n297), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n256), .A4(new_n304), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n300), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n308), .B1(new_n230), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n250), .ZN(new_n316));
  INV_X1    g130(.A(new_n213), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n209), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT12), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n316), .A2(KEYINPUT12), .B1(new_n319), .B2(new_n315), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n302), .A2(new_n304), .A3(new_n299), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G101), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n321), .A2(KEYINPUT79), .A3(new_n322), .A4(G101), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n325), .A2(new_n326), .B1(new_n199), .B2(new_n192), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n322), .B1(new_n321), .B2(G101), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT78), .B(new_n328), .C1(new_n306), .C2(new_n307), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n312), .A2(new_n313), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT78), .B1(new_n331), .B2(new_n328), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n327), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n212), .A2(new_n213), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n227), .B2(new_n229), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n314), .A2(new_n336), .B1(new_n308), .B2(new_n335), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n320), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G140), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G227), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n340), .B(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n317), .A2(new_n318), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n325), .A2(new_n326), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n200), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n331), .A2(new_n328), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n351), .B2(new_n329), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n336), .A2(new_n314), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n308), .A2(new_n335), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n346), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n338), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n345), .B1(new_n357), .B2(new_n344), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n292), .B1(new_n358), .B2(new_n284), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT81), .B1(new_n357), .B2(new_n344), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n361), .B(new_n343), .C1(new_n356), .C2(new_n338), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n316), .A2(KEYINPUT12), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n319), .A2(new_n315), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n338), .A2(new_n364), .A3(new_n343), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n320), .A2(KEYINPUT80), .A3(new_n338), .A4(new_n343), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n292), .B(new_n284), .C1(new_n363), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT82), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n334), .B1(new_n333), .B2(new_n337), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n344), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n361), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n357), .A2(KEYINPUT81), .A3(new_n344), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n368), .A2(new_n369), .ZN(new_n379));
  AOI21_X1  g193(.A(G902), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n292), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n359), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(KEYINPUT9), .B(G234), .Z(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT75), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n284), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G221), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(KEYINPUT76), .Z(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G217), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(G234), .B2(new_n284), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n394));
  INV_X1    g208(.A(G119), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G128), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n293), .A2(G119), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT24), .B(G110), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT72), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n397), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT23), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n396), .A2(KEYINPUT23), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n404), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n401), .B(new_n403), .C1(new_n407), .C2(G110), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(KEYINPUT73), .ZN(new_n409));
  XNOR2_X1  g223(.A(G125), .B(G140), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n193), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n413));
  INV_X1    g227(.A(G125), .ZN(new_n414));
  OR3_X1    g228(.A1(new_n414), .A2(KEYINPUT16), .A3(G140), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(G146), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT74), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n409), .A2(new_n411), .A3(new_n412), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n415), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(G146), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(G110), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n398), .B2(new_n399), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G137), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n341), .A2(G221), .A3(G234), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n418), .A2(new_n423), .A3(new_n427), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n394), .B1(new_n431), .B2(G902), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n429), .A2(KEYINPUT25), .A3(new_n284), .A4(new_n430), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n393), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n431), .A2(G902), .A3(new_n392), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(G110), .B(G122), .Z(new_n437));
  NAND2_X1  g251(.A1(new_n347), .A2(new_n219), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n351), .B2(new_n329), .ZN(new_n439));
  INV_X1    g253(.A(G116), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n440), .A2(KEYINPUT5), .A3(G119), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n216), .B2(KEYINPUT5), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n217), .B1(G113), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n314), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n437), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n437), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n330), .A2(new_n332), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n444), .B(new_n447), .C1(new_n448), .C2(new_n438), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n200), .A2(G125), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n244), .B2(G125), .ZN(new_n452));
  INV_X1    g266(.A(G224), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G953), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n452), .B(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(new_n437), .C1(new_n439), .C2(new_n445), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n456), .B1(KEYINPUT7), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n437), .B(KEYINPUT8), .Z(new_n461));
  NOR2_X1   g275(.A1(new_n314), .A2(new_n443), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n445), .B2(new_n462), .ZN(new_n463));
  OR3_X1    g277(.A1(new_n452), .A2(KEYINPUT7), .A3(new_n454), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n463), .A3(new_n449), .A4(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n284), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT83), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n466), .B(new_n469), .Z(new_n470));
  OAI21_X1  g284(.A(G214), .B1(G237), .B2(G902), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G237), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n341), .A3(G214), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n475), .A3(new_n195), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n254), .B(G214), .C1(KEYINPUT84), .C2(G143), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n210), .A3(new_n477), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT89), .B1(new_n479), .B2(new_n480), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n478), .A2(new_n484), .A3(KEYINPUT17), .A4(G131), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n420), .A2(new_n482), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n478), .A2(new_n487), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT18), .A2(G131), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n410), .B(new_n193), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n491), .B(new_n492), .C1(new_n488), .C2(new_n490), .ZN(new_n493));
  XNOR2_X1  g307(.A(G113), .B(G122), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT88), .B(G104), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n486), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n479), .A2(new_n481), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT19), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n410), .B1(KEYINPUT87), .B2(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n410), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n193), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n481), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n417), .A2(new_n501), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(new_n493), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n498), .B1(new_n509), .B2(new_n497), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT20), .ZN(new_n511));
  INV_X1    g325(.A(G475), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n284), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n515));
  INV_X1    g329(.A(new_n498), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n497), .B1(new_n508), .B2(new_n493), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n512), .B(new_n284), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n515), .B1(new_n518), .B2(KEYINPUT20), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n518), .A2(new_n515), .A3(KEYINPUT20), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G952), .ZN(new_n523));
  AOI211_X1 g337(.A(G953), .B(new_n523), .C1(G234), .C2(G237), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT21), .B(G898), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI211_X1 g340(.A(new_n284), .B(new_n341), .C1(G234), .C2(G237), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G478), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(KEYINPUT15), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G122), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G116), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT91), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n535), .A2(KEYINPUT14), .A3(G107), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n440), .A2(G122), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT92), .B1(new_n293), .B2(G143), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n195), .A3(G128), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(G128), .B2(new_n195), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n543), .A2(G134), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n543), .A2(G134), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n537), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n296), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n535), .A2(G107), .A3(new_n537), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI221_X1 g364(.A(new_n538), .B1(new_n545), .B2(new_n546), .C1(new_n550), .C2(new_n536), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT93), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n542), .A2(new_n552), .B1(G128), .B2(new_n195), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n202), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n544), .A2(new_n548), .A3(new_n549), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n558), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n553), .B(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G134), .B1(new_n563), .B2(new_n555), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT94), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n551), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n385), .A2(G217), .A3(new_n341), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n564), .A3(KEYINPUT94), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n567), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n551), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n532), .B1(new_n574), .B2(new_n284), .ZN(new_n575));
  AOI211_X1 g389(.A(G902), .B(new_n531), .C1(new_n568), .C2(new_n573), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n486), .A2(new_n493), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n496), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n498), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n512), .B1(new_n580), .B2(new_n284), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n522), .A2(new_n529), .A3(new_n577), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n472), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n291), .A2(new_n390), .A3(new_n436), .A4(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  AOI22_X1  g400(.A1(new_n262), .A2(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n587));
  OAI21_X1  g401(.A(G472), .B1(new_n587), .B2(G902), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n436), .B(new_n588), .C1(new_n274), .C2(new_n276), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n466), .A2(new_n468), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT95), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n466), .A2(new_n468), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n466), .A2(new_n594), .A3(new_n468), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n471), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n590), .A2(new_n390), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n530), .A2(new_n284), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n574), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n568), .A2(KEYINPUT33), .A3(new_n573), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n600), .B1(new_n604), .B2(G478), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n574), .A2(new_n530), .A3(new_n284), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n582), .B1(new_n520), .B2(new_n521), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n599), .A2(new_n528), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT34), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  INV_X1    g427(.A(new_n577), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n518), .A2(KEYINPUT20), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n581), .B1(new_n615), .B2(new_n513), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n528), .B(KEYINPUT96), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n599), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G107), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NOR2_X1   g436(.A1(new_n428), .A2(KEYINPUT36), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT97), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n424), .B(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n625), .A2(new_n284), .A3(new_n393), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n434), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n628), .B(new_n588), .C1(new_n274), .C2(new_n276), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n390), .A4(new_n584), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G110), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G12));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n527), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n524), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n616), .B(new_n640), .C1(new_n575), .C2(new_n576), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n596), .A2(new_n642), .A3(new_n471), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n596), .A2(new_n642), .A3(KEYINPUT100), .A4(new_n471), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n647), .A2(new_n291), .A3(new_n390), .A4(new_n628), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  INV_X1    g463(.A(new_n609), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n577), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n471), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n640), .B(KEYINPUT39), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n390), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n628), .B(new_n652), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n470), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n286), .A2(new_n270), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n284), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n270), .B1(new_n241), .B2(new_n253), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n277), .A2(new_n278), .A3(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n654), .A2(new_n655), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n656), .A2(new_n658), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT102), .B(G143), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G45));
  NAND4_X1  g481(.A1(new_n605), .A2(new_n609), .A3(new_n606), .A4(new_n640), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n383), .A2(new_n668), .A3(new_n389), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n291), .A3(new_n598), .A4(new_n628), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  AOI22_X1  g485(.A1(new_n376), .A2(new_n377), .B1(new_n368), .B2(new_n369), .ZN(new_n672));
  OAI21_X1  g486(.A(G469), .B1(new_n672), .B2(G902), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n381), .B1(new_n380), .B2(new_n292), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n672), .A2(KEYINPUT82), .A3(G469), .A4(G902), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n387), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n597), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n607), .A2(new_n650), .A3(new_n528), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n291), .A2(new_n677), .A3(new_n436), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  INV_X1    g495(.A(new_n619), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n291), .A2(new_n677), .A3(new_n682), .A4(new_n436), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  INV_X1    g498(.A(new_n583), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n291), .A2(new_n677), .A3(new_n685), .A4(new_n628), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  NAND2_X1  g501(.A1(new_n287), .A2(new_n270), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n275), .B1(new_n264), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n272), .A2(new_n284), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(G472), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n436), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n677), .A2(new_n692), .A3(new_n618), .A4(new_n651), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT103), .B(G122), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G24));
  AND2_X1   g509(.A1(new_n691), .A2(new_n628), .ZN(new_n696));
  INV_X1    g510(.A(new_n668), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n677), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  INV_X1    g513(.A(new_n359), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n674), .B2(new_n675), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n372), .A2(new_n382), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n700), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n387), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT105), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n187), .B1(new_n587), .B2(new_n275), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n290), .A2(new_n278), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n471), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n470), .A2(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n709), .A2(new_n436), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n702), .A2(new_n705), .A3(new_n713), .A4(new_n387), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n707), .A2(new_n712), .A3(new_n697), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT42), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n291), .A2(new_n436), .A3(new_n711), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n707), .A2(new_n718), .A3(new_n697), .A4(new_n714), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n210), .ZN(G33));
  INV_X1    g535(.A(new_n717), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n707), .A3(new_n642), .A4(new_n714), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  XNOR2_X1  g538(.A(new_n358), .B(KEYINPUT45), .ZN(new_n725));
  OAI21_X1  g539(.A(G469), .B1(new_n725), .B2(G902), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT46), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(G469), .C1(new_n725), .C2(G902), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(new_n703), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n387), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n653), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n607), .B2(new_n609), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n607), .A2(new_n609), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT43), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n739), .B(new_n734), .C1(new_n607), .C2(new_n609), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n588), .B1(new_n274), .B2(new_n276), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n628), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n733), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(new_n711), .C1(new_n744), .C2(new_n743), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT108), .B(G137), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G39));
  AND3_X1   g562(.A1(new_n730), .A2(KEYINPUT47), .A3(new_n387), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT47), .B1(new_n730), .B2(new_n387), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n751), .A2(new_n291), .A3(new_n710), .A4(new_n470), .ZN(new_n752));
  INV_X1    g566(.A(new_n436), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n697), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n638), .A2(KEYINPUT112), .A3(new_n639), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT112), .B1(new_n638), .B2(new_n639), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n628), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n702), .A2(new_n705), .A3(new_n760), .A4(new_n387), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT113), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n663), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n597), .A2(new_n577), .A3(new_n650), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n761), .B2(KEYINPUT113), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n648), .A2(new_n670), .A3(new_n698), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n718), .A2(new_n707), .A3(new_n697), .A4(new_n714), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n769), .A2(new_n722), .B1(KEYINPUT42), .B2(new_n715), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n648), .A2(new_n670), .A3(new_n698), .ZN(new_n771));
  INV_X1    g585(.A(new_n663), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n761), .B2(KEYINPUT113), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n383), .A2(new_n704), .ZN(new_n774));
  AOI211_X1 g588(.A(KEYINPUT104), .B(new_n359), .C1(new_n372), .C2(new_n382), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n387), .A4(new_n760), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n773), .A2(new_n778), .A3(new_n764), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n771), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n577), .B(KEYINPUT111), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(new_n609), .ZN(new_n783));
  INV_X1    g597(.A(new_n472), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n590), .A2(new_n390), .A3(new_n784), .A4(new_n618), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n633), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n585), .B1(new_n785), .B2(new_n610), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT110), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n585), .B(new_n789), .C1(new_n785), .C2(new_n610), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n786), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n768), .A2(new_n770), .A3(new_n781), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n707), .A2(new_n697), .A3(new_n691), .A4(new_n714), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n782), .A2(new_n616), .A3(new_n640), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n291), .A3(new_n390), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n627), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n711), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n679), .A2(new_n683), .A3(new_n686), .A4(new_n693), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n723), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n757), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n791), .A2(new_n781), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n780), .B1(new_n771), .B2(new_n779), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n720), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n798), .A2(new_n723), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n711), .B2(new_n796), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n801), .A2(new_n803), .A3(KEYINPUT53), .A4(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n800), .A2(new_n806), .A3(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT54), .B1(new_n800), .B2(new_n806), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n756), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n800), .A2(new_n806), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n800), .A2(new_n806), .A3(KEYINPUT54), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(KEYINPUT114), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  INV_X1    g629(.A(new_n676), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n741), .A2(new_n524), .A3(new_n816), .A4(new_n692), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n658), .A2(new_n471), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n818), .B1(new_n817), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n741), .A2(new_n524), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n824), .A2(new_n816), .A3(new_n711), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n696), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n772), .A2(new_n436), .A3(new_n524), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n816), .A2(new_n711), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n827), .A2(new_n828), .A3(new_n609), .A4(new_n608), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n751), .A2(KEYINPUT115), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n749), .B2(new_n750), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n703), .A2(new_n673), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT116), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n389), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n832), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n824), .A2(new_n692), .A3(new_n711), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n815), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n829), .B1(new_n821), .B2(new_n822), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n751), .A2(new_n837), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(KEYINPUT51), .A3(new_n826), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n523), .A2(G953), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n824), .A2(new_n677), .A3(new_n692), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n841), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n709), .A2(new_n436), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n825), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT48), .Z(new_n851));
  NOR3_X1   g665(.A1(new_n827), .A2(new_n610), .A3(new_n828), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n809), .A2(new_n814), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n523), .A2(new_n341), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n737), .A2(new_n436), .A3(new_n388), .A4(new_n471), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT109), .Z(new_n858));
  OR2_X1    g672(.A1(new_n835), .A2(KEYINPUT49), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n658), .B1(KEYINPUT49), .B2(new_n835), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n858), .A2(new_n772), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(G75));
  AOI21_X1  g680(.A(new_n284), .B1(new_n800), .B2(new_n806), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(G210), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(KEYINPUT118), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n450), .A2(new_n458), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n456), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT55), .Z(new_n873));
  AND2_X1   g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n870), .A2(new_n873), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT118), .B1(new_n868), .B2(new_n869), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n341), .A2(G952), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(G51));
  OAI21_X1  g692(.A(KEYINPUT57), .B1(new_n292), .B2(new_n284), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n812), .A2(new_n813), .A3(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n292), .A2(new_n284), .A3(KEYINPUT57), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n880), .A2(new_n881), .B1(new_n363), .B2(new_n370), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n867), .A2(G469), .A3(new_n725), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(G54));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT119), .B1(new_n885), .B2(new_n512), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n885), .A2(new_n512), .A3(KEYINPUT119), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n867), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n510), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT120), .Z(new_n891));
  INV_X1    g705(.A(new_n877), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n888), .B2(new_n889), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(G60));
  INV_X1    g708(.A(new_n604), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n600), .B(KEYINPUT59), .Z(new_n896));
  NAND4_X1  g710(.A1(new_n812), .A2(new_n895), .A3(new_n813), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n892), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n809), .A2(new_n814), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n895), .B1(new_n900), .B2(new_n896), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(G63));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n391), .A2(new_n284), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n810), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n877), .B1(new_n907), .B2(new_n625), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n431), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n908), .A2(new_n909), .B1(new_n910), .B2(KEYINPUT61), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(G66));
  AOI21_X1  g727(.A(new_n341), .B1(new_n525), .B2(G224), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n791), .A2(new_n798), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT124), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n917), .B2(new_n341), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n871), .B1(G898), .B2(new_n341), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n918), .B(new_n919), .Z(G69));
  XNOR2_X1  g734(.A(new_n771), .B(KEYINPUT125), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n732), .A2(new_n653), .A3(new_n849), .A4(new_n764), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n754), .A2(new_n746), .ZN(new_n924));
  INV_X1    g738(.A(new_n723), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n720), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n341), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n242), .B1(new_n252), .B2(KEYINPUT30), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n505), .Z(new_n929));
  OAI211_X1 g743(.A(new_n927), .B(new_n929), .C1(new_n637), .C2(new_n341), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n921), .A2(new_n665), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n783), .A2(new_n610), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n722), .A2(new_n654), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n924), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(G953), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n930), .B(new_n931), .C1(new_n938), .C2(new_n929), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n341), .B1(G227), .B2(G900), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G72));
  NAND2_X1  g755(.A1(new_n926), .A2(new_n916), .ZN(new_n942));
  NAND2_X1  g756(.A1(G472), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT63), .Z(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT127), .Z(new_n945));
  AOI21_X1  g759(.A(new_n281), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n877), .B1(new_n946), .B2(new_n270), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n282), .A2(new_n260), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n810), .A2(new_n944), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n934), .A2(new_n916), .A3(new_n937), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n945), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n661), .B2(new_n952), .ZN(G57));
endmodule


