//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OR2_X1    g0004(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n205), .A2(G50), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT64), .B(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR3_X1   g0013(.A1(new_n212), .A2(new_n213), .A3(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT0), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n207), .A2(new_n211), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n223), .B(new_n229), .C1(G97), .C2(G257), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(G1), .B2(G20), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n217), .B(new_n232), .C1(new_n216), .C2(new_n215), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  OAI211_X1 g0050(.A(new_n212), .B(G274), .C1(G41), .C2(G45), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT68), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n252), .B1(new_n258), .B2(new_n226), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G222), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n266), .B(new_n268), .C1(new_n269), .C2(new_n267), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(new_n253), .C1(G77), .C2(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n259), .A2(new_n260), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n261), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n259), .B(KEYINPUT69), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n271), .ZN(new_n277));
  OAI21_X1  g0077(.A(G190), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT74), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n209), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G1), .B2(new_n213), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G13), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n285), .A2(new_n213), .A3(G1), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n225), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n284), .A2(KEYINPUT72), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT72), .B1(new_n284), .B2(new_n288), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT64), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n294), .A2(new_n300), .B1(G150), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n282), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n279), .B1(new_n292), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n281), .ZN(new_n307));
  INV_X1    g0107(.A(new_n291), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n289), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT74), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n278), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n276), .A2(new_n275), .A3(new_n271), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n305), .A2(new_n310), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT9), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n313), .A2(new_n314), .A3(new_n317), .A4(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(new_n278), .A3(new_n317), .A4(new_n312), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n315), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n304), .B2(new_n292), .ZN(new_n326));
  AOI21_X1  g0126(.A(G179), .B1(new_n315), .B2(new_n316), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n264), .A2(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(G232), .B2(new_n267), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n228), .B2(new_n267), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(new_n253), .C1(G107), .C2(new_n266), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n257), .A2(G244), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n335), .A2(new_n252), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G200), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT15), .B(G87), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n300), .A2(new_n341), .B1(G77), .B2(new_n208), .ZN(new_n342));
  INV_X1    g0142(.A(new_n301), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n293), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n281), .B1(new_n219), .B2(new_n286), .ZN(new_n345));
  INV_X1    g0145(.A(new_n283), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G77), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n337), .A2(KEYINPUT73), .A3(G190), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT73), .B1(new_n337), .B2(G190), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n339), .B(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n323), .A2(new_n329), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n262), .ZN(new_n355));
  NAND2_X1  g0155(.A1(KEYINPUT76), .A2(G33), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(KEYINPUT3), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n226), .A2(G1698), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n269), .A2(new_n267), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n357), .A2(new_n330), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n253), .ZN(new_n363));
  INV_X1    g0163(.A(G232), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n253), .A2(new_n256), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n252), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(KEYINPUT78), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT68), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n251), .B(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n362), .B2(new_n253), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n366), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n368), .B1(new_n375), .B2(new_n324), .ZN(new_n376));
  INV_X1    g0176(.A(G58), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n227), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n201), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n301), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(KEYINPUT76), .A2(G33), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT76), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n263), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n298), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G68), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n357), .A2(new_n330), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n390), .B2(new_n213), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n382), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT3), .B1(new_n355), .B2(new_n356), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT7), .B(new_n298), .C1(new_n393), .C2(new_n265), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n387), .B1(new_n266), .B2(G20), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n381), .B1(new_n396), .B2(G68), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n281), .B(new_n392), .C1(new_n397), .C2(KEYINPUT16), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n294), .A2(new_n346), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT71), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n293), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n286), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n398), .A2(KEYINPUT77), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT77), .B1(new_n398), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n376), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT18), .ZN(new_n408));
  INV_X1    g0208(.A(G200), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n373), .B1(new_n372), .B2(new_n366), .ZN(new_n410));
  INV_X1    g0210(.A(new_n253), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n360), .B2(new_n361), .ZN(new_n412));
  NOR4_X1   g0212(.A1(new_n412), .A2(KEYINPUT78), .A3(new_n371), .A4(new_n365), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n367), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n398), .A2(new_n404), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n398), .A2(new_n404), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n414), .B2(new_n417), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n376), .B(new_n426), .C1(new_n405), .C2(new_n406), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n408), .A2(new_n422), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT14), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n371), .B1(G238), .B2(new_n257), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n364), .A2(G1698), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n266), .B(new_n433), .C1(G226), .C2(G1698), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n431), .B(new_n432), .C1(new_n436), .C2(new_n411), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n411), .B1(new_n434), .B2(new_n435), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n252), .B1(new_n258), .B2(new_n228), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT13), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n430), .B1(new_n441), .B2(G169), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G179), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT75), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n432), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n431), .B(new_n446), .C1(new_n436), .C2(new_n411), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n438), .A2(new_n439), .B1(new_n445), .B2(new_n432), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n441), .A2(new_n430), .A3(G169), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n443), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI22_X1  g0252(.A1(new_n299), .A2(new_n219), .B1(new_n225), .B2(new_n343), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n213), .A2(G68), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n281), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT11), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n455), .A2(new_n456), .B1(new_n227), .B2(new_n283), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n455), .A2(new_n456), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n212), .A3(G13), .ZN(new_n459));
  XOR2_X1   g0259(.A(new_n459), .B(KEYINPUT12), .Z(new_n460));
  NOR3_X1   g0260(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n452), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n441), .A2(G200), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n447), .A2(new_n448), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G190), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n338), .A2(new_n324), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n337), .A2(new_n444), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n348), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n429), .A2(new_n463), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n353), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT7), .B1(new_n332), .B2(new_n213), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n264), .B1(new_n383), .B2(new_n384), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n208), .B1(new_n474), .B2(new_n331), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n475), .B2(KEYINPUT7), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT79), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n396), .A2(new_n479), .A3(G107), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  XOR2_X1   g0281(.A(G97), .B(G107), .Z(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(KEYINPUT6), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n208), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n301), .A2(G77), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n478), .A2(new_n480), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n212), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n287), .A2(new_n282), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n486), .A2(new_n281), .B1(G97), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G97), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n286), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT80), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n255), .A2(G1), .ZN(new_n495));
  AND2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  NOR2_X1   g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n411), .A2(new_n498), .A3(G257), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n499), .B(KEYINPUT81), .ZN(new_n500));
  INV_X1    g0300(.A(G274), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G250), .A2(G1698), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n332), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n386), .A2(G244), .A3(new_n267), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT4), .ZN(new_n509));
  AOI211_X1 g0309(.A(new_n504), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n500), .B(new_n502), .C1(new_n510), .C2(new_n411), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n324), .ZN(new_n512));
  INV_X1    g0312(.A(new_n511), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n444), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n494), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(G200), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n503), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n253), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(G190), .A3(new_n502), .A4(new_n500), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n490), .A2(new_n516), .A3(new_n520), .A4(new_n493), .ZN(new_n521));
  INV_X1    g0321(.A(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n222), .A2(new_n267), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n357), .A2(new_n330), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G294), .B1(new_n383), .B2(new_n384), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n411), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n502), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n411), .A2(G264), .A3(new_n498), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(KEYINPUT84), .A3(new_n409), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n530), .B2(new_n416), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n530), .A2(G200), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(G116), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n355), .B2(new_n356), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n213), .B1(new_n538), .B2(KEYINPUT23), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n330), .A2(new_n331), .A3(G87), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n540), .A2(new_n541), .B1(new_n208), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n357), .A2(new_n298), .A3(KEYINPUT22), .A4(new_n330), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n545), .A2(new_n221), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT83), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n477), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n544), .A2(new_n546), .A3(new_n547), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n539), .B(new_n543), .C1(new_n545), .C2(new_n221), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT83), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT24), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  OAI211_X1 g0355(.A(KEYINPUT83), .B(new_n555), .C1(new_n552), .C2(new_n549), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n281), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT25), .B1(new_n287), .B2(G107), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n287), .A2(KEYINPUT25), .A3(G107), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n489), .B2(G107), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n536), .A2(new_n557), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n411), .A2(G270), .A3(new_n498), .ZN(new_n562));
  INV_X1    g0362(.A(G264), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G1698), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n522), .A2(new_n267), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n357), .A2(new_n330), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G303), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n266), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n562), .B1(new_n568), .B2(new_n253), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n502), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n489), .A2(G116), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n286), .A2(new_n537), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n298), .B(new_n503), .C1(G33), .C2(new_n491), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n280), .A2(new_n209), .B1(G20), .B2(new_n537), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n572), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n571), .B(new_n579), .C1(new_n416), .C2(new_n570), .ZN(new_n580));
  AND4_X1   g0380(.A1(new_n515), .A2(new_n521), .A3(new_n561), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n530), .A2(G169), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n444), .B2(new_n530), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g0385(.A1(KEYINPUT82), .A2(KEYINPUT21), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n570), .A2(new_n578), .A3(G169), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(KEYINPUT82), .A2(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n570), .A2(new_n444), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n578), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n324), .B1(new_n569), .B2(new_n502), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(KEYINPUT82), .A3(KEYINPUT21), .A4(new_n578), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n495), .A2(G274), .ZN(new_n596));
  OR3_X1    g0396(.A1(new_n253), .A2(new_n222), .A3(new_n495), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G238), .A2(G1698), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n220), .B2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n538), .B1(new_n386), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n596), .B(new_n597), .C1(new_n600), .C2(new_n411), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G190), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n386), .A2(G68), .A3(new_n298), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n299), .B2(new_n491), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n221), .A2(new_n491), .A3(new_n477), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n435), .A2(new_n605), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n208), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n604), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n281), .B1(new_n286), .B2(new_n340), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n489), .A2(G87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n601), .A2(G200), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n603), .A2(new_n611), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n489), .A2(new_n341), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n602), .A2(new_n444), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n601), .A2(new_n324), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n585), .A2(new_n595), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n472), .A2(new_n581), .A3(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n470), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n452), .A2(new_n462), .B1(new_n467), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n425), .A2(new_n422), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT18), .B1(new_n376), .B2(new_n423), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n324), .B1(new_n410), .B2(new_n413), .ZN(new_n627));
  INV_X1    g0427(.A(new_n368), .ZN(new_n628));
  AND4_X1   g0428(.A1(KEYINPUT18), .A2(new_n423), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n328), .B1(new_n630), .B2(new_n323), .ZN(new_n631));
  INV_X1    g0431(.A(new_n472), .ZN(new_n632));
  INV_X1    g0432(.A(new_n521), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT86), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT85), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n618), .B(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n616), .A2(new_n617), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n614), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n637), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(KEYINPUT86), .A3(new_n614), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n633), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n585), .A2(new_n595), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n561), .ZN(new_n646));
  INV_X1    g0446(.A(new_n515), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n643), .B(new_n644), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n620), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n638), .B1(new_n649), .B2(KEYINPUT26), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n631), .B1(new_n632), .B2(new_n651), .ZN(G369));
  NOR2_X1   g0452(.A1(new_n208), .A2(new_n285), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n212), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n653), .A2(KEYINPUT87), .A3(new_n654), .A4(new_n212), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n654), .B1(new_n653), .B2(new_n212), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n662), .A2(KEYINPUT88), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT88), .ZN(new_n665));
  INV_X1    g0465(.A(G213), .ZN(new_n666));
  AOI211_X1 g0466(.A(new_n666), .B(new_n660), .C1(new_n657), .C2(new_n658), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n667), .B2(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n579), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(new_n594), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n580), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n669), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n582), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n561), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n585), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n582), .A2(new_n669), .A3(new_n584), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n595), .A2(new_n674), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n678), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0486(.A(new_n214), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n607), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n207), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n674), .B1(new_n648), .B2(new_n650), .ZN(new_n694));
  OR3_X1    g0494(.A1(new_n694), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n640), .A2(new_n642), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n638), .B1(new_n697), .B2(KEYINPUT26), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n647), .A2(new_n644), .A3(new_n620), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT26), .B1(new_n643), .B2(new_n646), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n647), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .A3(new_n669), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT91), .B1(new_n694), .B2(KEYINPUT29), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n695), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n511), .A2(new_n570), .A3(new_n531), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n444), .A3(new_n601), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n527), .A2(new_n529), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n570), .A2(new_n444), .A3(new_n601), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n513), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n513), .A2(KEYINPUT30), .A3(new_n708), .A4(new_n707), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n706), .A2(new_n711), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n674), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n581), .A2(new_n621), .A3(new_n669), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n704), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n693), .B1(new_n725), .B2(G1), .ZN(G364));
  NAND2_X1  g0526(.A1(new_n653), .A2(G45), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n689), .A2(G1), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n673), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n672), .A2(G330), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n209), .B1(G20), .B2(new_n324), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n298), .A2(new_n444), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n416), .A2(new_n409), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n298), .A2(G190), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G179), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(G326), .A2(new_n735), .B1(new_n739), .B2(G329), .ZN(new_n740));
  INV_X1    g0540(.A(G322), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n732), .A2(G190), .A3(new_n409), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n732), .A2(new_n416), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n409), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G317), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(KEYINPUT33), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(KEYINPUT33), .B2(new_n747), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n744), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G311), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n736), .A2(new_n444), .A3(G200), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G283), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n737), .A2(G190), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n208), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n266), .B1(new_n757), .B2(G294), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n749), .A2(new_n751), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n733), .A2(G20), .A3(new_n444), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n743), .B(new_n759), .C1(G303), .C2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n756), .B(KEYINPUT96), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n491), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(G68), .B2(new_n745), .ZN(new_n766));
  INV_X1    g0566(.A(new_n750), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n219), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT95), .B(G159), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n739), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT32), .Z(new_n771));
  AOI22_X1  g0571(.A1(new_n753), .A2(G107), .B1(new_n735), .B2(G50), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n742), .B(KEYINPUT94), .Z(new_n773));
  OAI211_X1 g0573(.A(new_n771), .B(new_n772), .C1(new_n377), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n760), .A2(new_n221), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n768), .A2(new_n774), .A3(new_n332), .A4(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n731), .B1(new_n762), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT92), .B1(G13), .B2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(KEYINPUT92), .A2(G13), .A3(G33), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n777), .B1(new_n672), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n246), .A2(G45), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n386), .A2(new_n687), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n785), .B(new_n786), .C1(G45), .C2(new_n207), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n266), .A2(new_n214), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(G116), .B2(new_n214), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n782), .A2(new_n731), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n728), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT93), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n729), .A2(new_n730), .B1(new_n784), .B2(new_n793), .ZN(G396));
  INV_X1    g0594(.A(KEYINPUT100), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n669), .B2(new_n349), .ZN(new_n796));
  OAI211_X1 g0596(.A(KEYINPUT100), .B(new_n348), .C1(new_n664), .C2(new_n668), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n796), .A2(new_n352), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n470), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n623), .A2(new_n669), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n694), .B(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n802), .A2(new_n724), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT101), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n802), .A2(new_n724), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(KEYINPUT101), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n804), .A2(new_n805), .A3(new_n728), .A4(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G150), .A2(new_n745), .B1(new_n750), .B2(new_n769), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  INV_X1    g0609(.A(G143), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n734), .C1(new_n773), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT34), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n386), .B1(new_n738), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(KEYINPUT99), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n814), .A2(KEYINPUT99), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(G58), .C2(new_n757), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n752), .A2(new_n227), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G50), .B2(new_n761), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n812), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n760), .A2(new_n477), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n266), .B(new_n765), .C1(G303), .C2(new_n735), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n221), .A2(new_n752), .B1(new_n742), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G311), .B2(new_n739), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G116), .A2(new_n750), .B1(new_n745), .B2(G283), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n821), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n781), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n731), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT97), .Z(new_n832));
  AOI22_X1  g0632(.A1(new_n829), .A2(new_n731), .B1(new_n219), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n728), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n833), .B(new_n834), .C1(new_n801), .C2(new_n781), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n807), .A2(new_n835), .ZN(G384));
  NOR2_X1   g0636(.A1(new_n463), .A2(new_n674), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n392), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n382), .B1(new_n389), .B2(new_n391), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT16), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n282), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT103), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT7), .B1(new_n386), .B2(G20), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n227), .B1(new_n390), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n381), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n281), .B1(new_n848), .B2(KEYINPUT16), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT103), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n403), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT104), .B1(new_n851), .B2(new_n662), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n843), .B(new_n281), .C1(new_n848), .C2(KEYINPUT16), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n392), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n840), .A2(new_n841), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n843), .B1(new_n855), .B2(new_n281), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n404), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n667), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT77), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n423), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n398), .A2(KEYINPUT77), .A3(new_n404), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n426), .B1(new_n864), .B2(new_n376), .ZN(new_n865));
  INV_X1    g0665(.A(new_n427), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n625), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n860), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n857), .A2(new_n376), .B1(new_n418), .B2(new_n419), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n852), .A2(new_n870), .A3(new_n859), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n662), .B1(new_n862), .B2(new_n863), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n424), .B1(new_n864), .B2(new_n376), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n871), .A2(KEYINPUT37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n869), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n871), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n874), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n852), .A2(new_n859), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n428), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT39), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n667), .B1(new_n405), .B2(new_n406), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n376), .A2(new_n423), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n420), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n626), .A2(new_n629), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n872), .B1(new_n625), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n869), .A2(new_n875), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT39), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n876), .B1(new_n869), .B2(new_n875), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT105), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT39), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n885), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT106), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n885), .A2(new_n905), .A3(new_n897), .A4(new_n902), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n838), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n694), .A2(new_n801), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n800), .ZN(new_n909));
  INV_X1    g0709(.A(new_n467), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n462), .B(new_n674), .C1(new_n452), .C2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n462), .B1(new_n664), .B2(new_n668), .ZN(new_n912));
  AOI211_X1 g0712(.A(KEYINPUT14), .B(new_n324), .C1(new_n437), .C2(new_n440), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n442), .A2(new_n913), .A3(new_n449), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n467), .B(new_n912), .C1(new_n914), .C2(new_n461), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n900), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n891), .A2(new_n662), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n907), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n695), .A2(new_n472), .A3(new_n703), .A4(new_n702), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n631), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n722), .A2(new_n721), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n916), .A2(new_n799), .A3(new_n800), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT107), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT40), .B1(new_n895), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n898), .A2(new_n929), .A3(new_n899), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n925), .A2(new_n926), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n929), .A2(KEYINPUT107), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n928), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n472), .A2(new_n925), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n934), .B(new_n935), .Z(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(G330), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n923), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n212), .B2(new_n653), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n210), .B(new_n208), .C1(new_n483), .C2(KEYINPUT35), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n537), .B(new_n940), .C1(KEYINPUT35), .C2(new_n483), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT102), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT36), .Z(new_n943));
  OAI21_X1  g0743(.A(G77), .B1(new_n377), .B2(new_n227), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n207), .A2(new_n944), .B1(G50), .B2(new_n227), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(G1), .A3(new_n285), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n943), .A3(new_n946), .ZN(G367));
  NOR2_X1   g0747(.A1(new_n764), .A2(new_n227), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G50), .B2(new_n750), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n761), .A2(G58), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n753), .A2(G77), .B1(new_n739), .B2(G137), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n810), .B2(new_n734), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(G150), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n266), .B1(new_n742), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n745), .B2(new_n769), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n949), .A2(new_n950), .A3(new_n953), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n760), .B2(new_n537), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n960), .C1(new_n746), .C2(new_n824), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT112), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n390), .B1(new_n738), .B2(new_n747), .ZN(new_n963));
  XOR2_X1   g0763(.A(KEYINPUT111), .B(G311), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n752), .A2(new_n491), .B1(new_n734), .B2(new_n965), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n963), .B(new_n966), .C1(G283), .C2(new_n750), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n962), .B(new_n967), .C1(new_n567), .C2(new_n773), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n756), .A2(new_n477), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n957), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n728), .B1(new_n971), .B2(new_n731), .ZN(new_n972));
  INV_X1    g0772(.A(new_n786), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n791), .B1(new_n214), .B2(new_n340), .C1(new_n973), .C2(new_n240), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n669), .B1(new_n611), .B2(new_n612), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n638), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n697), .B2(new_n975), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n972), .B(new_n974), .C1(new_n783), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n727), .A2(G1), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n647), .A2(new_n674), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n674), .A2(new_n494), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n515), .A3(new_n521), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n684), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT45), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT109), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n684), .A2(new_n988), .A3(new_n984), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n684), .B2(new_n984), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n991), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n993), .A2(KEYINPUT44), .A3(new_n989), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n986), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n681), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n683), .A2(KEYINPUT110), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(new_n673), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n679), .A2(new_n682), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n681), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n986), .A2(new_n992), .A3(new_n994), .A4(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n996), .A2(new_n725), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n725), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n688), .B(KEYINPUT41), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n979), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n683), .A2(KEYINPUT42), .A3(new_n984), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT108), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT42), .B1(new_n683), .B2(new_n984), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(KEYINPUT108), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n515), .B1(new_n982), .B2(new_n585), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n669), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n681), .A2(new_n983), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1014), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n978), .B1(new_n1006), .B2(new_n1022), .ZN(G387));
  NOR2_X1   g0823(.A1(new_n679), .A2(new_n783), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n786), .B1(new_n237), .B2(new_n255), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n690), .B2(new_n789), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n227), .A2(new_n219), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n293), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n225), .ZN(new_n1029));
  AOI211_X1 g0829(.A(G116), .B(new_n607), .C1(new_n1029), .C2(KEYINPUT50), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1030), .B(new_n255), .C1(KEYINPUT50), .C2(new_n1029), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1026), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n687), .A2(new_n477), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n782), .B(new_n731), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G303), .A2(new_n750), .B1(new_n745), .B2(new_n964), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n741), .B2(new_n734), .C1(new_n773), .C2(new_n747), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n824), .B2(new_n760), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G283), .B2(new_n757), .ZN(new_n1039));
  XOR2_X1   g0839(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n386), .B1(new_n739), .B2(G326), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n537), .C2(new_n752), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n746), .A2(new_n401), .B1(new_n491), .B2(new_n752), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n764), .A2(new_n340), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G68), .C2(new_n750), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n761), .A2(G77), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n742), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1048), .A2(G50), .B1(new_n735), .B2(G159), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n954), .B2(new_n738), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1046), .A2(new_n1047), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1043), .B1(new_n390), .B2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1024), .B(new_n1034), .C1(new_n1053), .C2(new_n731), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(new_n834), .B1(new_n1000), .B2(new_n979), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1000), .A2(new_n725), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n688), .B(KEYINPUT114), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1000), .A2(new_n725), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1055), .B1(new_n1059), .B2(new_n1060), .ZN(G393));
  INV_X1    g0861(.A(KEYINPUT115), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n996), .A2(new_n1062), .A3(new_n1002), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1062), .B2(new_n1002), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1056), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1003), .B(new_n1058), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n984), .A2(new_n782), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n791), .B1(new_n491), .B2(new_n214), .C1(new_n973), .C2(new_n249), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n266), .B1(new_n761), .B2(G283), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n738), .B2(new_n741), .C1(new_n477), .C2(new_n752), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT117), .Z(new_n1071));
  OAI22_X1  g0871(.A1(new_n824), .A2(new_n767), .B1(new_n746), .B2(new_n567), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G116), .B2(new_n757), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1048), .A2(G311), .B1(new_n735), .B2(G317), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1071), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1048), .A2(G159), .B1(new_n735), .B2(G150), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(KEYINPUT51), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n390), .B(new_n1079), .C1(G68), .C2(new_n761), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n764), .A2(new_n219), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1028), .B2(new_n750), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n752), .A2(new_n221), .B1(new_n738), .B2(new_n810), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1078), .B2(KEYINPUT51), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n746), .A2(new_n225), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1077), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n728), .B1(new_n1087), .B2(new_n731), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1067), .A2(new_n1068), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1064), .B2(new_n979), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1066), .A2(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n935), .A2(G330), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n921), .A2(new_n1093), .A3(new_n631), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n801), .A2(G330), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n916), .A3(new_n925), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n723), .A2(new_n1096), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n916), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n909), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n916), .B1(new_n1096), .B2(new_n925), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1098), .B2(new_n916), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n701), .A2(new_n669), .A3(new_n799), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1103), .A2(new_n800), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1092), .B1(new_n1095), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n909), .A2(new_n916), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n838), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n904), .A2(new_n906), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n895), .A2(new_n837), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n916), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1098), .A2(new_n916), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1097), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1107), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1097), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n909), .A2(new_n1099), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT118), .B1(new_n1122), .B2(new_n1094), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1117), .A2(new_n1124), .A3(new_n1058), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n904), .A2(new_n830), .A3(new_n906), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1081), .A2(new_n266), .A3(new_n775), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n739), .A2(G294), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1048), .A2(G116), .B1(new_n735), .B2(G283), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n491), .A2(new_n767), .B1(new_n746), .B2(new_n477), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n818), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n266), .B1(new_n752), .B2(new_n225), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1136));
  INV_X1    g0936(.A(G125), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1137), .A2(new_n738), .B1(new_n734), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n761), .A2(G150), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n742), .A2(new_n813), .B1(new_n1140), .B2(KEYINPUT53), .ZN(new_n1141));
  NOR4_X1   g0941(.A1(new_n1135), .A2(new_n1136), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT54), .B(G143), .Z(new_n1143));
  AOI22_X1  g0943(.A1(new_n763), .A2(G159), .B1(new_n750), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(new_n809), .C2(new_n746), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1140), .A2(KEYINPUT53), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1132), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1147), .A2(new_n731), .B1(new_n401), .B2(new_n832), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1126), .A2(new_n834), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n979), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1125), .A2(new_n1151), .ZN(G378));
  AOI21_X1  g0952(.A(new_n901), .B1(new_n900), .B2(KEYINPUT39), .ZN(new_n1153));
  AOI211_X1 g0953(.A(KEYINPUT105), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n905), .B1(new_n1155), .B2(new_n897), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n906), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n837), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n934), .A2(G330), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n305), .A2(new_n310), .A3(new_n667), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT56), .Z(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT55), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n323), .B2(new_n329), .ZN(new_n1164));
  AOI211_X1 g0964(.A(KEYINPUT55), .B(new_n328), .C1(new_n320), .C2(new_n322), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n329), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(KEYINPUT55), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n323), .A2(new_n1163), .A3(new_n329), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1171), .A3(new_n1161), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1159), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n934), .A2(G330), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n919), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1158), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1175), .B1(new_n934), .B2(G330), .ZN(new_n1180));
  INV_X1    g0980(.A(G330), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1181), .B(new_n1173), .C1(new_n928), .C2(new_n933), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n907), .B2(new_n919), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT121), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1179), .A2(new_n1184), .A3(KEYINPUT121), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1058), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1120), .A2(new_n1121), .A3(new_n1106), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n1095), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1189), .B1(new_n1193), .B2(new_n979), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1057), .A2(new_n1190), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1094), .B1(new_n1150), .B2(new_n1106), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT122), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1179), .A2(new_n1184), .A3(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1183), .B(KEYINPUT122), .C1(new_n907), .C2(new_n919), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1195), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n948), .B1(new_n341), .B2(new_n750), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n491), .B2(new_n746), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n739), .A2(G283), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1047), .A2(new_n254), .A3(new_n390), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT120), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n753), .A2(G58), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n477), .B2(new_n742), .C1(new_n537), .C2(new_n734), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT58), .Z(new_n1210));
  NAND2_X1  g1010(.A1(new_n761), .A2(new_n1143), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n734), .B2(new_n1137), .C1(new_n1138), .C2(new_n742), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n764), .A2(new_n954), .B1(new_n809), .B2(new_n767), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G132), .C2(new_n745), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT59), .ZN(new_n1215));
  AOI21_X1  g1015(.A(G41), .B1(new_n739), .B2(G124), .ZN(new_n1216));
  AOI21_X1  g1016(.A(G33), .B1(new_n753), .B2(new_n769), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G41), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1210), .B(new_n1218), .C1(G50), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n728), .B1(new_n1220), .B2(new_n731), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n831), .A2(new_n225), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n1173), .C2(new_n781), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1194), .A2(new_n1201), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(G375));
  NAND2_X1  g1025(.A1(new_n1095), .A2(new_n1106), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1122), .A2(new_n1094), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1005), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1112), .A2(new_n830), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n746), .A2(new_n537), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1230), .B(new_n1045), .C1(G107), .C2(new_n750), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1048), .A2(G283), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n738), .A2(new_n567), .B1(new_n491), .B2(new_n760), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT123), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n332), .B1(new_n734), .B2(new_n824), .C1(new_n219), .C2(new_n752), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1234), .B2(new_n1233), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1231), .A2(new_n1232), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n767), .A2(new_n954), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n734), .A2(new_n813), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n764), .A2(new_n225), .B1(new_n1240), .B2(KEYINPUT124), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(KEYINPUT124), .B2(new_n1240), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n390), .B1(new_n761), .B2(G159), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1207), .B(new_n1243), .C1(new_n1138), .C2(new_n738), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n745), .B2(new_n1143), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1242), .B(new_n1245), .C1(new_n809), .C2(new_n773), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1238), .B1(new_n1239), .B2(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1247), .A2(new_n731), .B1(new_n227), .B2(new_n832), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1229), .A2(new_n834), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1106), .B2(new_n979), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1228), .A2(new_n1250), .ZN(G381));
  NAND2_X1  g1051(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1125), .A2(new_n1151), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(G375), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1005), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1003), .B2(new_n725), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1020), .B(new_n1021), .C1(new_n1259), .C2(new_n979), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1260), .A2(new_n978), .A3(new_n1090), .A4(new_n1066), .ZN(new_n1261));
  INV_X1    g1061(.A(G384), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1250), .A3(new_n1228), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(new_n1261), .A2(G396), .A3(G393), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1257), .A2(new_n1264), .ZN(G407));
  OAI21_X1  g1065(.A(new_n1257), .B1(new_n663), .B2(new_n1264), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(G213), .ZN(G409));
  INV_X1    g1067(.A(KEYINPUT127), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(G390), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(G396), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1261), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1269), .B2(new_n1261), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1268), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1261), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1270), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1269), .A2(new_n1270), .A3(new_n1261), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(KEYINPUT127), .A3(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1273), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1192), .A2(new_n1095), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT121), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1179), .A2(new_n1184), .A3(KEYINPUT121), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1281), .B(new_n1005), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1198), .A2(new_n979), .A3(new_n1199), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1223), .A3(new_n1285), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1224), .A2(G378), .B1(new_n1255), .B2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n666), .A2(G343), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT126), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1253), .B1(new_n1125), .B2(new_n1151), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1254), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1286), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1194), .A2(new_n1201), .A3(G378), .A4(new_n1223), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1288), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1289), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1227), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1122), .A2(KEYINPUT60), .A3(new_n1094), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(new_n1058), .A3(new_n1226), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1250), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1262), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1280), .B1(new_n1297), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1288), .A2(G2897), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1303), .B(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1289), .A2(new_n1296), .A3(new_n1308), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1303), .B(new_n1288), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1310), .B2(new_n1280), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1279), .B1(new_n1305), .B2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1304), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1310), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT63), .B1(new_n1294), .B2(new_n1307), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1314), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1313), .A2(new_n1320), .ZN(G405));
  NAND2_X1  g1121(.A1(new_n1273), .A2(new_n1278), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1322), .B(new_n1293), .C1(new_n1224), .C2(new_n1256), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1293), .B1(new_n1256), .B2(new_n1224), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1279), .A2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1323), .A2(new_n1325), .A3(new_n1304), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1304), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


