//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n463), .B1(new_n470), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AOI211_X1 g047(.A(KEYINPUT68), .B(new_n472), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT3), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT70), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(new_n464), .A3(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(G137), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n476), .A2(new_n477), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G101), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n474), .A2(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n478), .A2(new_n482), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(new_n472), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n488), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  OAI21_X1  g071(.A(G2104), .B1(new_n472), .B2(G114), .ZN(new_n497));
  NOR2_X1   g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n498), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(G2104), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n472), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n499), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n478), .A2(G126), .A3(G2105), .A4(new_n482), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT4), .A2(G138), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n478), .A2(new_n472), .A3(new_n482), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(G543), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n521), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n514), .A2(new_n516), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n529), .B1(new_n525), .B2(new_n530), .C1(new_n531), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n519), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n522), .A2(new_n537), .B1(new_n538), .B2(new_n525), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  INV_X1    g115(.A(new_n525), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n522), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n519), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(KEYINPUT73), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n525), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n556), .ZN(new_n559));
  NAND4_X1  g134(.A1(new_n521), .A2(new_n559), .A3(G53), .A4(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n522), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n532), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n566), .A2(KEYINPUT74), .A3(G651), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT74), .B1(new_n566), .B2(G651), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n561), .B(new_n563), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n570), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G299));
  OR2_X1    g148(.A1(new_n536), .A2(new_n539), .ZN(G301));
  OR2_X1    g149(.A1(new_n520), .A2(new_n526), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT76), .ZN(G303));
  NAND2_X1  g151(.A1(new_n562), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n541), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n562), .A2(G86), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n541), .A2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n517), .A2(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT77), .Z(new_n585));
  AND2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n581), .B(new_n582), .C1(new_n586), .C2(new_n519), .ZN(G305));
  AOI22_X1  g162(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n519), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n522), .A2(new_n590), .B1(new_n591), .B2(new_n525), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n589), .A2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n522), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n532), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(G54), .A2(new_n541), .B1(new_n598), .B2(G651), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT10), .B1(new_n522), .B2(new_n594), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  XNOR2_X1  g181(.A(G299), .B(KEYINPUT78), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(new_n601), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  OAI221_X1 g187(.A(new_n542), .B1(new_n543), .B2(new_n522), .C1(new_n519), .C2(new_n545), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n602), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n601), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n489), .A2(G123), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n491), .A2(G135), .ZN(new_n620));
  OR2_X1    g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n489), .A2(new_n623), .A3(G123), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n619), .A2(new_n620), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT80), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT3), .B(G2104), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n484), .A2(new_n628), .A3(new_n472), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT13), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n627), .A2(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2438), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2430), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  AOI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n650), .B(KEYINPUT17), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n652), .B1(new_n654), .B2(new_n651), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  INV_X1    g231(.A(new_n650), .ZN(new_n657));
  INV_X1    g232(.A(new_n651), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(new_n649), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n649), .A3(new_n651), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n656), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT83), .B(G2096), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT19), .Z(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n672), .A2(new_n673), .B1(new_n668), .B2(new_n674), .ZN(new_n675));
  OR3_X1    g250(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n675), .B(new_n676), .C1(new_n673), .C2(new_n672), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT85), .B(G1986), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(KEYINPUT23), .A3(G20), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT23), .ZN(new_n688));
  INV_X1    g263(.A(G20), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(G16), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n571), .A2(new_n572), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n687), .B(new_n690), .C1(new_n691), .C2(new_n686), .ZN(new_n692));
  INV_X1    g267(.A(G1956), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n610), .A2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G4), .B2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G1348), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G19), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n547), .B2(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G1341), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT31), .B(G11), .Z(new_n702));
  OR2_X1    g277(.A1(G29), .A2(G33), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT25), .Z(new_n705));
  AOI22_X1  g280(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n478), .A2(new_n482), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(new_n472), .ZN(new_n708));
  INV_X1    g283(.A(G139), .ZN(new_n709));
  OAI221_X1 g284(.A(new_n705), .B1(new_n472), .B2(new_n706), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n703), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G2072), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n702), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n696), .A2(new_n697), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  NAND2_X1  g291(.A1(G164), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G27), .B2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G2078), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND4_X1   g295(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n694), .A2(new_n698), .A3(new_n701), .A4(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT92), .B1(G29), .B2(G32), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n489), .A2(G129), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT26), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n707), .A2(G141), .B1(G105), .B2(new_n484), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n725), .B(new_n728), .C1(new_n729), .C2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(new_n711), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n730), .B(KEYINPUT91), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n734), .A2(KEYINPUT92), .A3(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT27), .B(G1996), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G5), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G171), .B2(G16), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G1961), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G34), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n742), .A2(new_n743), .A3(new_n711), .ZN(new_n744));
  INV_X1    g319(.A(G160), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n711), .ZN(new_n746));
  INV_X1    g321(.A(G2084), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n740), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n737), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n733), .A2(new_n735), .ZN(new_n752));
  INV_X1    g327(.A(new_n736), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n754));
  INV_X1    g329(.A(G26), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G29), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(G29), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT89), .ZN(new_n758));
  INV_X1    g333(.A(G140), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n708), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n489), .A2(G128), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n491), .A2(KEYINPUT89), .A3(G140), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n760), .A2(new_n761), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n757), .B1(new_n765), .B2(G29), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n756), .B1(new_n766), .B2(new_n754), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n752), .A2(new_n753), .B1(G2067), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n711), .A2(G35), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n495), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT29), .B(G2090), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n770), .B(new_n771), .Z(new_n772));
  NAND2_X1  g347(.A1(G168), .A2(G16), .ZN(new_n773));
  OR2_X1    g348(.A1(G16), .A2(G21), .ZN(new_n774));
  AOI21_X1  g349(.A(G1966), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n719), .B2(new_n718), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G28), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G28), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n780), .A2(new_n781), .A3(new_n711), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n782), .B1(new_n625), .B2(new_n711), .C1(new_n775), .C2(new_n776), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n773), .A2(G1966), .A3(new_n774), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n772), .A2(new_n778), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n767), .A2(G2067), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n768), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n723), .A2(new_n751), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n520), .A2(new_n526), .A3(new_n686), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G22), .ZN(new_n792));
  OAI21_X1  g367(.A(KEYINPUT86), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n791), .A2(KEYINPUT86), .A3(new_n792), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n791), .A2(KEYINPUT86), .A3(new_n792), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n797), .A2(G1971), .A3(new_n793), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT34), .ZN(new_n800));
  OR2_X1    g375(.A1(G16), .A2(G23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G288), .B2(new_n686), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G305), .A2(G16), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n686), .A2(G6), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  AND3_X1   g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n805), .B2(new_n806), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n799), .A2(new_n800), .A3(new_n804), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n686), .A2(G24), .ZN(new_n812));
  INV_X1    g387(.A(G290), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n686), .ZN(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n711), .A2(G25), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n489), .A2(G119), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n491), .A2(G131), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n817), .B1(new_n822), .B2(new_n711), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n811), .A2(new_n816), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT87), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n811), .A2(KEYINPUT87), .A3(new_n816), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n794), .A2(new_n795), .A3(new_n790), .ZN(new_n832));
  AOI21_X1  g407(.A(G1971), .B1(new_n797), .B2(new_n793), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n810), .B(new_n804), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT88), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT36), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT36), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n831), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n789), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n739), .A2(G1961), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n746), .A2(new_n747), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n700), .A2(G1341), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(G311));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT95), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n749), .B(KEYINPUT94), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n848), .A2(new_n787), .A3(new_n722), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n831), .A2(new_n839), .A3(new_n836), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n839), .B1(new_n831), .B2(new_n836), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n849), .B(new_n844), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n842), .A4(new_n843), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n847), .A2(new_n855), .ZN(G150));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  INV_X1    g432(.A(G67), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n532), .B2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(KEYINPUT96), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(KEYINPUT96), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(G651), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  INV_X1    g439(.A(G55), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n522), .A2(new_n864), .B1(new_n865), .B2(new_n525), .ZN(new_n866));
  OAI21_X1  g441(.A(G860), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NOR2_X1   g443(.A1(new_n601), .A2(new_n611), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT39), .ZN(new_n872));
  INV_X1    g447(.A(new_n866), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n613), .A2(new_n873), .A3(new_n862), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n613), .B1(new_n862), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n868), .B1(new_n878), .B2(G860), .ZN(G145));
  XNOR2_X1  g454(.A(new_n745), .B(new_n495), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n511), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n507), .A2(new_n508), .A3(new_n510), .A4(KEYINPUT98), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n734), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n732), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n710), .A2(KEYINPUT99), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n710), .A2(KEYINPUT100), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n765), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  INV_X1    g468(.A(new_n765), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n892), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n886), .A3(new_n888), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n489), .A2(G130), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n491), .A2(G142), .ZN(new_n901));
  NOR2_X1   g476(.A1(G106), .A2(G2105), .ZN(new_n902));
  OAI21_X1  g477(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n900), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(new_n630), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n630), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(new_n822), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n822), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n899), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n896), .A2(new_n898), .A3(new_n911), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n625), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n625), .B1(new_n913), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n881), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n915), .A3(new_n880), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  NAND2_X1  g500(.A1(G299), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n571), .A2(KEYINPUT102), .A3(new_n572), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n610), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n610), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n877), .B(new_n615), .ZN(new_n932));
  INV_X1    g507(.A(new_n926), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n927), .A2(new_n610), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(KEYINPUT41), .A3(new_n928), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n934), .B(new_n926), .ZN(new_n938));
  INV_X1    g513(.A(new_n932), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT103), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n575), .B(G288), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(G305), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G290), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n945), .A2(G305), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(G305), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n813), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT42), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n942), .A2(new_n944), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n942), .B2(new_n944), .ZN(new_n954));
  OAI21_X1  g529(.A(G868), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n602), .B1(new_n863), .B2(new_n866), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(G295));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n956), .ZN(G331));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n951), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n947), .A2(KEYINPUT105), .A3(new_n950), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G301), .A2(G168), .ZN(new_n965));
  NAND2_X1  g540(.A1(G171), .A2(G286), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n875), .B2(new_n876), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n547), .B1(new_n863), .B2(new_n866), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(new_n874), .A3(new_n965), .A4(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n967), .B(KEYINPUT104), .C1(new_n875), .C2(new_n876), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(new_n935), .A3(new_n928), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n938), .A2(KEYINPUT106), .A3(new_n974), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n968), .A2(new_n970), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n931), .A2(new_n936), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n964), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n974), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n931), .A2(new_n936), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n938), .A2(new_n968), .A3(new_n970), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n951), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n921), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n960), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n963), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT105), .B1(new_n947), .B2(new_n950), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n981), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n977), .A2(new_n978), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(KEYINPUT107), .A3(new_n921), .A4(new_n986), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n959), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n964), .B1(new_n984), .B2(new_n985), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(new_n987), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT44), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT43), .B1(new_n997), .B2(new_n987), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n994), .A2(new_n921), .A3(new_n986), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(KEYINPUT43), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(new_n1005), .ZN(G397));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n885), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n483), .A2(new_n485), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n472), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n628), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT68), .B1(new_n1013), .B2(new_n472), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n470), .A2(new_n463), .A3(G2105), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT108), .B(G40), .Z(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1010), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1010), .A2(KEYINPUT109), .A3(new_n1019), .ZN(new_n1023));
  INV_X1    g598(.A(G1996), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n734), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n765), .B(G2067), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1022), .A2(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(new_n1024), .A3(new_n734), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(KEYINPUT110), .A3(new_n1028), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n822), .B(new_n825), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(G290), .B(G1986), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1020), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1031), .A2(new_n1032), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1039), .B(KEYINPUT111), .Z(new_n1040));
  AOI211_X1 g615(.A(new_n1009), .B(G1384), .C1(new_n883), .C2(new_n884), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n511), .A2(new_n1007), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1009), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n474), .A2(new_n486), .A3(new_n1017), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(G1971), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n511), .A2(new_n1049), .A3(new_n1007), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT113), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n511), .A2(new_n1053), .A3(new_n1049), .A4(new_n1007), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(new_n1052), .A3(new_n1044), .A4(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1055), .A2(G2090), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1047), .A2(KEYINPUT112), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1048), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1059), .B(KEYINPUT55), .Z(new_n1060));
  NAND3_X1  g635(.A1(new_n1058), .A2(G8), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1060), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1052), .A2(new_n1044), .A3(new_n1050), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G2090), .ZN(new_n1064));
  OAI21_X1  g639(.A(G8), .B1(new_n1047), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G8), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1042), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1044), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1976), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(G288), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  INV_X1    g647(.A(G288), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(G1976), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1071), .A2(KEYINPUT52), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(G305), .B(G1981), .ZN(new_n1076));
  NOR2_X1   g651(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n1077));
  XOR2_X1   g652(.A(new_n1076), .B(new_n1077), .Z(new_n1078));
  AOI211_X1 g653(.A(new_n1072), .B(new_n1075), .C1(new_n1078), .C2(new_n1069), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1061), .A2(new_n1066), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1055), .A2(new_n697), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1044), .A2(new_n1068), .A3(KEYINPUT117), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1019), .B2(new_n1042), .ZN(new_n1084));
  INV_X1    g659(.A(G2067), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n610), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n569), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n569), .B2(KEYINPUT116), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1019), .B1(new_n1009), .B2(new_n1042), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1063), .A2(new_n693), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI211_X1 g674(.A(KEYINPUT118), .B(new_n1091), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1088), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1095), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1041), .A2(new_n1045), .A3(G1996), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT119), .B(G1341), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT58), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT120), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT117), .B1(new_n1044), .B2(new_n1068), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1019), .A2(new_n1083), .A3(new_n1042), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1092), .A2(new_n1093), .A3(new_n1024), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n547), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT59), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1109), .A2(new_n1115), .A3(new_n1118), .A4(new_n547), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1102), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1097), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT121), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(new_n1121), .C1(new_n1122), .C2(new_n1097), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n610), .B1(new_n1087), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1081), .A2(new_n1086), .A3(KEYINPUT60), .A4(new_n601), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1087), .A2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1120), .A2(new_n1124), .A3(new_n1126), .A4(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1102), .A2(KEYINPUT61), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT122), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1137), .B(new_n1134), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1103), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(G171), .B(KEYINPUT54), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT53), .B1(new_n1046), .B2(new_n719), .ZN(new_n1142));
  INV_X1    g717(.A(G1961), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1055), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1045), .B1(KEYINPUT45), .B2(new_n1068), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(KEYINPUT53), .A3(new_n719), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n1148));
  OAI21_X1  g723(.A(G2105), .B1(new_n470), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1013), .A2(KEYINPUT125), .ZN(new_n1150));
  OAI21_X1  g725(.A(G40), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1041), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT53), .B(new_n719), .C1(new_n486), .C2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1153), .B2(new_n486), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1010), .A3(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1144), .A2(new_n1141), .A3(new_n1156), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1145), .A2(G1966), .B1(G2084), .B2(new_n1055), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G8), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT51), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(G286), .A2(G8), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1159), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1166));
  OAI211_X1 g741(.A(G8), .B(new_n1162), .C1(new_n1158), .C2(G286), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1158), .A2(G8), .A3(G286), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1147), .B(new_n1157), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1140), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT62), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1168), .A2(new_n1175), .A3(new_n1169), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1173), .A2(G171), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1080), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1159), .A2(G286), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1080), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1058), .A2(G8), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1179), .B1(new_n1183), .B2(new_n1062), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1184), .A2(new_n1061), .A3(new_n1079), .A4(new_n1180), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g761(.A(G1976), .B(G288), .C1(new_n1078), .C2(new_n1069), .ZN(new_n1187));
  NOR2_X1   g762(.A1(G305), .A2(G1981), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT115), .Z(new_n1189));
  OR2_X1    g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1061), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1069), .A2(new_n1190), .B1(new_n1191), .B2(new_n1079), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1186), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1040), .B1(new_n1178), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n822), .A2(new_n825), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT126), .Z(new_n1196));
  NAND3_X1  g771(.A1(new_n1031), .A2(new_n1032), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n894), .A2(new_n1085), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT127), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1197), .A2(new_n1201), .A3(new_n1198), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1200), .A2(new_n1034), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT46), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1026), .A2(new_n732), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1205), .B1(new_n1033), .B2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT47), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1020), .A2(new_n815), .A3(new_n813), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT48), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1031), .A2(new_n1032), .A3(new_n1036), .A4(new_n1210), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1203), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1194), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g788(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1215));
  NAND4_X1  g789(.A1(new_n1003), .A2(new_n922), .A3(new_n684), .A4(new_n1215), .ZN(G225));
  INV_X1    g790(.A(G225), .ZN(G308));
endmodule


