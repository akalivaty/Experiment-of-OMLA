

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n370), .B(n331), .ZN(n335) );
  XNOR2_X1 U324 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U325 ( .A(n346), .B(n345), .Z(n556) );
  XOR2_X1 U326 ( .A(KEYINPUT25), .B(n463), .Z(n291) );
  INV_X1 U327 ( .A(KEYINPUT54), .ZN(n432) );
  INV_X1 U328 ( .A(KEYINPUT71), .ZN(n401) );
  XNOR2_X1 U329 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U330 ( .A(n335), .B(n334), .ZN(n339) );
  INV_X1 U331 ( .A(KEYINPUT64), .ZN(n435) );
  XNOR2_X1 U332 ( .A(n404), .B(n403), .ZN(n405) );
  NOR2_X1 U333 ( .A1(n476), .A2(n583), .ZN(n477) );
  NOR2_X1 U334 ( .A1(n473), .A2(n472), .ZN(n486) );
  NOR2_X1 U335 ( .A1(n464), .A2(n451), .ZN(n565) );
  XNOR2_X1 U336 ( .A(KEYINPUT38), .B(n479), .ZN(n499) );
  XNOR2_X1 U337 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U338 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n480) );
  XNOR2_X1 U339 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(G15GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n292), .B(G113GAT), .ZN(n400) );
  XOR2_X1 U343 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n294) );
  XNOR2_X1 U344 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U346 ( .A(n295), .B(G183GAT), .Z(n297) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(G176GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n426) );
  XNOR2_X1 U349 ( .A(n400), .B(n426), .ZN(n306) );
  XOR2_X1 U350 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n299) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U353 ( .A(n300), .B(KEYINPUT65), .Z(n304) );
  XNOR2_X1 U354 ( .A(G99GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n301), .B(G120GAT), .ZN(n369) );
  XNOR2_X1 U356 ( .A(G134GAT), .B(G127GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n302), .B(KEYINPUT0), .ZN(n320) );
  XNOR2_X1 U358 ( .A(n369), .B(n320), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X2 U360 ( .A(n306), .B(n305), .Z(n525) );
  INV_X1 U361 ( .A(n525), .ZN(n464) );
  XOR2_X1 U362 ( .A(G148GAT), .B(G120GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(G141GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U365 ( .A(G29GAT), .B(G85GAT), .Z(n309) );
  XNOR2_X1 U366 ( .A(n310), .B(n309), .ZN(n326) );
  XOR2_X1 U367 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n312) );
  XNOR2_X1 U368 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U370 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n314) );
  XNOR2_X1 U371 ( .A(G1GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n324) );
  XOR2_X1 U374 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n322) );
  XOR2_X1 U375 ( .A(KEYINPUT2), .B(G162GAT), .Z(n318) );
  XNOR2_X1 U376 ( .A(KEYINPUT91), .B(G155GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U378 ( .A(KEYINPUT3), .B(n319), .Z(n445) );
  XNOR2_X1 U379 ( .A(n320), .B(n445), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n328) );
  NAND2_X1 U383 ( .A1(G225GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n513) );
  XOR2_X1 U385 ( .A(KEYINPUT82), .B(KEYINPUT9), .Z(n330) );
  XNOR2_X1 U386 ( .A(G190GAT), .B(G162GAT), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n346) );
  XOR2_X1 U388 ( .A(G85GAT), .B(G92GAT), .Z(n370) );
  XOR2_X1 U389 ( .A(G43GAT), .B(G134GAT), .Z(n331) );
  XOR2_X1 U390 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n333) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G218GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U393 ( .A(KEYINPUT66), .B(KEYINPUT81), .Z(n337) );
  NAND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  XOR2_X1 U395 ( .A(n337), .B(n336), .Z(n338) );
  XNOR2_X1 U396 ( .A(n339), .B(n338), .ZN(n344) );
  XOR2_X1 U397 ( .A(KEYINPUT8), .B(G50GAT), .Z(n341) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(G29GAT), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U400 ( .A(KEYINPUT7), .B(n342), .Z(n397) );
  XNOR2_X1 U401 ( .A(n397), .B(G106GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  INV_X1 U403 ( .A(n556), .ZN(n410) );
  XNOR2_X1 U404 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n347) );
  XOR2_X1 U405 ( .A(n410), .B(n347), .Z(n583) );
  XOR2_X1 U406 ( .A(G78GAT), .B(G211GAT), .Z(n349) );
  XNOR2_X1 U407 ( .A(G183GAT), .B(G71GAT), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U409 ( .A(n350), .B(G155GAT), .Z(n352) );
  XOR2_X1 U410 ( .A(G1GAT), .B(G8GAT), .Z(n393) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(n393), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n357) );
  XNOR2_X1 U413 ( .A(G57GAT), .B(G64GAT), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n353), .B(KEYINPUT13), .ZN(n371) );
  XOR2_X1 U415 ( .A(n371), .B(KEYINPUT12), .Z(n355) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U418 ( .A(n357), .B(n356), .Z(n365) );
  XOR2_X1 U419 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n359) );
  XNOR2_X1 U420 ( .A(G15GAT), .B(G127GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U422 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n361) );
  XNOR2_X1 U423 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U426 ( .A(n365), .B(n364), .Z(n533) );
  NOR2_X1 U427 ( .A1(n583), .A2(n533), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n366), .B(KEYINPUT45), .ZN(n385) );
  XNOR2_X1 U429 ( .A(G106GAT), .B(G78GAT), .ZN(n367) );
  XOR2_X1 U430 ( .A(n367), .B(G148GAT), .Z(n437) );
  INV_X1 U431 ( .A(n437), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n384) );
  XOR2_X1 U433 ( .A(n371), .B(n370), .Z(n373) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U436 ( .A(KEYINPUT32), .B(KEYINPUT80), .Z(n375) );
  NAND2_X1 U437 ( .A1(G230GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U439 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U440 ( .A(KEYINPUT33), .B(KEYINPUT77), .Z(n379) );
  XNOR2_X1 U441 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n380), .B(KEYINPUT31), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n454) );
  NAND2_X1 U446 ( .A1(n385), .A2(n454), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n386), .B(KEYINPUT111), .ZN(n407) );
  XOR2_X1 U448 ( .A(KEYINPUT74), .B(KEYINPUT29), .Z(n388) );
  XNOR2_X1 U449 ( .A(KEYINPUT75), .B(KEYINPUT70), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U451 ( .A(KEYINPUT72), .B(KEYINPUT68), .Z(n390) );
  XNOR2_X1 U452 ( .A(KEYINPUT73), .B(KEYINPUT69), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n406) );
  XOR2_X1 U455 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XOR2_X1 U456 ( .A(n438), .B(n393), .Z(n395) );
  NAND2_X1 U457 ( .A1(G229GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U459 ( .A(n396), .B(G197GAT), .Z(n399) );
  XNOR2_X1 U460 ( .A(G169GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n400), .B(KEYINPUT30), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n570) );
  XNOR2_X1 U464 ( .A(KEYINPUT76), .B(n570), .ZN(n559) );
  INV_X1 U465 ( .A(n559), .ZN(n527) );
  NAND2_X1 U466 ( .A1(n407), .A2(n527), .ZN(n415) );
  XOR2_X1 U467 ( .A(KEYINPUT47), .B(KEYINPUT110), .Z(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT41), .B(n454), .ZN(n564) );
  AND2_X1 U469 ( .A1(n564), .A2(n570), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n408), .B(KEYINPUT46), .ZN(n409) );
  INV_X1 U471 ( .A(n533), .ZN(n578) );
  NOR2_X1 U472 ( .A1(n409), .A2(n578), .ZN(n411) );
  NAND2_X1 U473 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  NAND2_X1 U475 ( .A1(n415), .A2(n414), .ZN(n416) );
  XOR2_X1 U476 ( .A(KEYINPUT48), .B(n416), .Z(n543) );
  XOR2_X1 U477 ( .A(KEYINPUT98), .B(G64GAT), .Z(n418) );
  NAND2_X1 U478 ( .A1(G226GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U480 ( .A(n419), .B(G92GAT), .Z(n424) );
  XOR2_X1 U481 ( .A(KEYINPUT83), .B(KEYINPUT97), .Z(n421) );
  XNOR2_X1 U482 ( .A(G8GAT), .B(KEYINPUT96), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U484 ( .A(G36GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n431) );
  XOR2_X1 U487 ( .A(KEYINPUT90), .B(G204GAT), .Z(n428) );
  XNOR2_X1 U488 ( .A(G197GAT), .B(G211GAT), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U490 ( .A(G218GAT), .B(KEYINPUT21), .Z(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n448) );
  XOR2_X2 U492 ( .A(n431), .B(n448), .Z(n515) );
  INV_X1 U493 ( .A(n515), .ZN(n460) );
  NOR2_X1 U494 ( .A1(n543), .A2(n460), .ZN(n433) );
  NOR2_X1 U495 ( .A1(n513), .A2(n434), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n569) );
  XNOR2_X1 U497 ( .A(KEYINPUT23), .B(n437), .ZN(n440) );
  XNOR2_X1 U498 ( .A(G50GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n442) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n447) );
  XNOR2_X1 U504 ( .A(n445), .B(KEYINPUT24), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n465) );
  NOR2_X1 U507 ( .A1(n569), .A2(n465), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NAND2_X1 U509 ( .A1(n565), .A2(n556), .ZN(n453) );
  INV_X1 U510 ( .A(n454), .ZN(n575) );
  NOR2_X1 U511 ( .A1(n527), .A2(n575), .ZN(n487) );
  INV_X1 U512 ( .A(KEYINPUT104), .ZN(n475) );
  XOR2_X1 U513 ( .A(KEYINPUT27), .B(n515), .Z(n467) );
  INV_X1 U514 ( .A(n467), .ZN(n455) );
  NAND2_X1 U515 ( .A1(n455), .A2(n513), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n456), .B(KEYINPUT99), .ZN(n545) );
  XNOR2_X1 U517 ( .A(n465), .B(KEYINPUT67), .ZN(n457) );
  XOR2_X1 U518 ( .A(n457), .B(KEYINPUT28), .Z(n519) );
  INV_X1 U519 ( .A(n519), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n545), .A2(n458), .ZN(n524) );
  XNOR2_X1 U521 ( .A(n525), .B(KEYINPUT88), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n524), .A2(n459), .ZN(n473) );
  INV_X1 U523 ( .A(KEYINPUT101), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n464), .A2(n460), .ZN(n461) );
  XNOR2_X1 U525 ( .A(n461), .B(KEYINPUT100), .ZN(n462) );
  NOR2_X1 U526 ( .A1(n465), .A2(n462), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT26), .ZN(n568) );
  NOR2_X1 U529 ( .A1(n467), .A2(n568), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n291), .A2(n468), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n513), .A2(n469), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n578), .A2(n486), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT37), .B(n477), .Z(n512) );
  NAND2_X1 U536 ( .A1(n487), .A2(n512), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(KEYINPUT105), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n525), .A2(n499), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n565), .A2(n578), .ZN(n483) );
  XNOR2_X1 U540 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1350GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n489) );
  NOR2_X1 U543 ( .A1(n556), .A2(n533), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NOR2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n501) );
  AND2_X1 U546 ( .A1(n487), .A2(n501), .ZN(n494) );
  NAND2_X1 U547 ( .A1(n494), .A2(n513), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U549 ( .A(G1GAT), .B(n490), .Z(G1324GAT) );
  NAND2_X1 U550 ( .A1(n494), .A2(n515), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .Z(n493) );
  NAND2_X1 U553 ( .A1(n494), .A2(n525), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n519), .A2(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  NAND2_X1 U558 ( .A1(n513), .A2(n499), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n515), .A2(n499), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n499), .A2(n519), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U564 ( .A(n564), .ZN(n530) );
  NOR2_X1 U565 ( .A1(n570), .A2(n530), .ZN(n511) );
  AND2_X1 U566 ( .A1(n511), .A2(n501), .ZN(n508) );
  NAND2_X1 U567 ( .A1(n508), .A2(n513), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n502), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(G64GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U572 ( .A1(n508), .A2(n515), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n525), .A2(n508), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U577 ( .A1(n508), .A2(n519), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  AND2_X1 U579 ( .A1(n512), .A2(n511), .ZN(n520) );
  NAND2_X1 U580 ( .A1(n513), .A2(n520), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n515), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(KEYINPUT108), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n525), .A2(n520), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n522) );
  NAND2_X1 U588 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n543), .A2(n524), .ZN(n526) );
  NAND2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n539) );
  NOR2_X1 U593 ( .A1(n527), .A2(n539), .ZN(n528) );
  XOR2_X1 U594 ( .A(KEYINPUT112), .B(n528), .Z(n529) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n539), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n539), .ZN(n538) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(KEYINPUT113), .B(n536), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1342GAT) );
  NOR2_X1 U605 ( .A1(n410), .A2(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n543), .A2(n568), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(KEYINPUT117), .B(n546), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n557), .A2(n570), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT118), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT52), .B(n551), .Z(n553) );
  NAND2_X1 U619 ( .A1(n557), .A2(n564), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT121), .Z(n555) );
  NAND2_X1 U622 ( .A1(n557), .A2(n578), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n565), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n562) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n563), .Z(n567) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  XOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT60), .Z(n572) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  INV_X1 U646 ( .A(n581), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

