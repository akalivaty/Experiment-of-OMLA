//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT64), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n210), .B(new_n211), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n209), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n226), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n222), .A2(new_n223), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NOR2_X1   g0051(.A1(new_n202), .A2(new_n213), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G58), .A2(G68), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n254), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT16), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n228), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT7), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT73), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n262), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(KEYINPUT73), .A3(new_n264), .ZN(new_n269));
  AND4_X1   g0069(.A1(KEYINPUT74), .A2(new_n268), .A3(G68), .A4(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT7), .B1(new_n273), .B2(new_n228), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n213), .B1(new_n274), .B2(KEYINPUT73), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT74), .B1(new_n275), .B2(new_n268), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n258), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n280), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n279), .A2(new_n227), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n267), .ZN(new_n284));
  OAI21_X1  g0084(.A(G68), .B1(new_n274), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT16), .B1(new_n285), .B2(new_n256), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n277), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n227), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(KEYINPUT67), .B2(new_n278), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  INV_X1    g0091(.A(G1), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n290), .A2(new_n291), .A3(new_n293), .A4(new_n281), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n279), .A2(new_n281), .A3(new_n227), .A4(new_n293), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT68), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT8), .B(G58), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n292), .A2(G20), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT69), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n297), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n299), .A2(new_n293), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(KEYINPUT75), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT75), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n299), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(new_n294), .B2(new_n296), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n308), .B2(new_n303), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n288), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT76), .ZN(new_n313));
  OR2_X1    g0113(.A1(G223), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n314), .B1(G226), .B2(new_n315), .C1(new_n271), .C2(new_n272), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G41), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G1), .A3(G13), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n292), .B1(G41), .B2(G45), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G274), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n289), .B2(new_n321), .ZN(new_n327));
  INV_X1    g0127(.A(new_n323), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n325), .A2(G232), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n313), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n322), .B1(new_n316), .B2(new_n317), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n322), .A3(G274), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n324), .B2(new_n236), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT76), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n312), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n331), .A2(new_n333), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n311), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT18), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT18), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n311), .A2(new_n343), .A3(new_n340), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n330), .B2(new_n334), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n288), .A2(new_n310), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT17), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n305), .A2(new_n309), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n269), .A2(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n275), .A2(KEYINPUT74), .A3(new_n268), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n282), .B1(new_n359), .B2(new_n258), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n353), .B1(new_n360), .B2(new_n287), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n349), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n342), .A2(new_n344), .A3(new_n352), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n332), .B1(new_n324), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n273), .A2(new_n315), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(G223), .B1(G77), .B2(new_n273), .ZN(new_n368));
  INV_X1    g0168(.A(G222), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n261), .A2(new_n262), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n315), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n366), .B1(new_n372), .B2(new_n319), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n337), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G169), .B2(new_n373), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n297), .A2(G50), .A3(new_n301), .ZN(new_n376));
  OAI21_X1  g0176(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n377));
  INV_X1    g0177(.A(G150), .ZN(new_n378));
  INV_X1    g0178(.A(new_n255), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n228), .A2(G33), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n377), .B1(new_n378), .B2(new_n379), .C1(new_n298), .C2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n293), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n381), .A2(new_n283), .B1(new_n201), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(KEYINPUT9), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(KEYINPUT9), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n373), .A2(G190), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n373), .A2(new_n345), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n386), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT10), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(KEYINPUT10), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n385), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n236), .A2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n370), .B(new_n394), .C1(G226), .C2(G1698), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n322), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n332), .B1(new_n324), .B2(new_n214), .ZN(new_n398));
  OR3_X1    g0198(.A1(new_n397), .A2(KEYINPUT13), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT13), .B1(new_n397), .B2(new_n398), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(KEYINPUT71), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(KEYINPUT13), .C1(new_n397), .C2(new_n398), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n401), .A2(G200), .A3(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n399), .A2(G190), .A3(new_n400), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n255), .A2(G50), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT72), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n380), .A2(new_n215), .B1(new_n228), .B2(G68), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n283), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT11), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n382), .A2(new_n213), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT12), .ZN(new_n414));
  INV_X1    g0214(.A(new_n295), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(G68), .A3(new_n301), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n411), .A2(new_n412), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n404), .A2(new_n405), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n401), .A2(G169), .A3(new_n403), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n401), .A2(new_n421), .A3(G169), .A4(new_n403), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n399), .A2(G179), .A3(new_n400), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n418), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n370), .A2(G232), .A3(new_n315), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT70), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n367), .A2(G238), .B1(G107), .B2(new_n273), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n322), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n332), .B1(new_n324), .B2(new_n216), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n312), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n429), .A2(new_n430), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n337), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n415), .A2(G77), .A3(new_n301), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT15), .B(G87), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n436), .A2(new_n380), .B1(new_n228), .B2(new_n215), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n299), .B2(new_n255), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n435), .B1(G77), .B2(new_n293), .C1(new_n438), .C2(new_n282), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n432), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n431), .A2(G200), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n433), .B2(G190), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n364), .A2(new_n393), .A3(new_n425), .A4(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(G238), .B(new_n315), .C1(new_n271), .C2(new_n272), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G116), .ZN(new_n447));
  OAI21_X1  g0247(.A(G244), .B1(new_n271), .B2(new_n272), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n315), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n319), .ZN(new_n450));
  INV_X1    g0250(.A(G45), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n326), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n322), .C1(G250), .C2(new_n452), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT79), .B1(new_n455), .B2(new_n347), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n450), .A2(new_n457), .A3(G190), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(G200), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n370), .A2(new_n228), .A3(G68), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT19), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n228), .B1(new_n396), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(G87), .B2(new_n207), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n380), .B2(new_n205), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n283), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n436), .A2(new_n382), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n292), .A2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n415), .A2(G87), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n456), .A2(new_n458), .A3(new_n459), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n455), .A2(new_n312), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n295), .B1(new_n292), .B2(G33), .ZN(new_n473));
  INV_X1    g0273(.A(new_n436), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n467), .A3(new_n466), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n472), .B(new_n476), .C1(G179), .C2(new_n455), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n471), .A2(KEYINPUT80), .A3(new_n477), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n448), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n216), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n370), .A2(new_n315), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n370), .A2(G250), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n315), .B1(new_n489), .B2(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n319), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT5), .B(G41), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n452), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G257), .A3(new_n322), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n327), .A2(new_n452), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n312), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n448), .A2(new_n483), .B1(G33), .B2(G283), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n483), .B1(new_n370), .B2(G250), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n500), .B(new_n486), .C1(new_n315), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n496), .B1(new_n502), .B2(new_n319), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n337), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n505), .A2(new_n205), .A3(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(G97), .B(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n508), .A2(new_n228), .B1(new_n215), .B2(new_n379), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n206), .B1(new_n265), .B2(new_n267), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n283), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n473), .A2(G97), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n293), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n499), .A2(new_n504), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT78), .ZN(new_n517));
  INV_X1    g0317(.A(new_n515), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n503), .A2(G190), .ZN(new_n519));
  OAI21_X1  g0319(.A(G200), .B1(new_n503), .B2(KEYINPUT77), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n491), .A2(KEYINPUT77), .A3(new_n497), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT78), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n499), .A2(new_n504), .A3(new_n515), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n228), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G20), .B2(new_n447), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n228), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n370), .A2(new_n228), .A3(G87), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n531), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(KEYINPUT82), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n282), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT82), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n536), .A2(new_n538), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(new_n531), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n541), .B1(new_n539), .B2(KEYINPUT82), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n473), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n293), .A2(G107), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT25), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n370), .A2(G257), .A3(G1698), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n370), .A2(G250), .A3(new_n315), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G294), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n319), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(KEYINPUT83), .A3(new_n319), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n319), .B1(new_n452), .B2(new_n492), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G264), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n564), .A2(new_n495), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G169), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n558), .A2(new_n319), .B1(G264), .B2(new_n563), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G179), .A3(new_n495), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n554), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n552), .B1(new_n542), .B2(new_n547), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n561), .A2(new_n347), .A3(new_n565), .A4(new_n562), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n559), .A2(new_n495), .A3(new_n564), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n345), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n563), .A2(G270), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n579), .A2(new_n495), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n370), .A2(G264), .A3(G1698), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n370), .A2(G257), .A3(new_n315), .ZN(new_n582));
  INV_X1    g0382(.A(G303), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n370), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n319), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n312), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n473), .A2(G116), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n382), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(G20), .B1(G33), .B2(G283), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n260), .A2(G97), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(G20), .B2(new_n588), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n283), .A2(KEYINPUT20), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT20), .B1(new_n283), .B2(new_n592), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n587), .B(new_n589), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n580), .A2(G179), .A3(new_n585), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n596), .A2(new_n597), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n586), .A2(new_n595), .A3(KEYINPUT21), .ZN(new_n600));
  INV_X1    g0400(.A(new_n595), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n580), .A2(new_n585), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n601), .B(new_n603), .C1(new_n347), .C2(new_n602), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n599), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n578), .A2(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n445), .A2(new_n482), .A3(new_n526), .A4(new_n606), .ZN(G372));
  NAND2_X1  g0407(.A1(new_n424), .A2(new_n417), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n418), .B2(new_n440), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n362), .A2(new_n352), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n361), .A2(KEYINPUT18), .A3(new_n339), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n343), .B1(new_n311), .B2(new_n340), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n391), .A2(new_n392), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n385), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n517), .A2(new_n524), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(KEYINPUT26), .A3(new_n480), .A4(new_n481), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n470), .A2(new_n459), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n455), .A2(new_n347), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n477), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n620), .B1(new_n625), .B2(new_n516), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n574), .A2(new_n337), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(G169), .B2(new_n566), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n599), .B(new_n600), .C1(new_n629), .C2(new_n572), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n623), .B1(new_n572), .B2(new_n576), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n526), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n627), .A2(new_n632), .A3(new_n477), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n445), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n617), .A2(new_n634), .ZN(G369));
  NAND3_X1  g0435(.A1(new_n292), .A2(new_n228), .A3(G13), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT27), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT85), .ZN(new_n640));
  INV_X1    g0440(.A(G213), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n640), .A2(G343), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n601), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n599), .A2(new_n600), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n605), .B2(new_n645), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n644), .A2(new_n572), .ZN(new_n650));
  OAI22_X1  g0450(.A1(new_n578), .A2(new_n650), .B1(new_n571), .B2(new_n644), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n643), .B1(new_n599), .B2(new_n600), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n571), .A3(new_n577), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n554), .A2(new_n644), .A3(new_n570), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n224), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G1), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n230), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT28), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n633), .A2(new_n644), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT29), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n606), .A2(new_n482), .A3(new_n526), .A4(new_n644), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT30), .ZN(new_n669));
  INV_X1    g0469(.A(new_n455), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n503), .A2(new_n670), .A3(new_n568), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n580), .A2(G179), .A3(new_n585), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n568), .A2(new_n450), .A3(new_n454), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n598), .A2(new_n674), .A3(KEYINPUT30), .A4(new_n503), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n670), .A2(G179), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(new_n498), .A3(new_n574), .A4(new_n602), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n643), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT31), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n668), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n630), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n631), .A2(new_n517), .A3(new_n524), .A4(new_n522), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n477), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n618), .A2(new_n620), .A3(new_n480), .A4(new_n481), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT26), .B1(new_n625), .B2(new_n516), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n644), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT29), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n667), .A2(new_n684), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT86), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT86), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n667), .A2(new_n695), .A3(new_n684), .A4(new_n692), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n665), .B1(new_n697), .B2(G1), .ZN(G364));
  AND2_X1   g0498(.A1(new_n228), .A2(G13), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n292), .B1(new_n699), .B2(G45), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n660), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n370), .A2(new_n224), .ZN(new_n703));
  INV_X1    g0503(.A(G355), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n703), .A2(new_n704), .B1(G116), .B2(new_n224), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n247), .A2(G45), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n273), .A2(new_n224), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(new_n451), .B2(new_n231), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(G13), .A2(G33), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n227), .B1(G20), .B2(new_n312), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT87), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n702), .B1(new_n709), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT32), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n228), .A2(G179), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G190), .A2(G200), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT89), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT89), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(KEYINPUT90), .B(G159), .Z(new_n725));
  AOI21_X1  g0525(.A(new_n717), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n228), .A2(new_n337), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G200), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT88), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n347), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n726), .B1(G50), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G87), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n718), .A2(G190), .A3(G200), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n718), .A2(new_n347), .A3(G200), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n206), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n727), .A2(new_n719), .ZN(new_n737));
  INV_X1    g0537(.A(new_n727), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n345), .A2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n370), .B1(new_n215), .B2(new_n737), .C1(new_n741), .C2(new_n202), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n730), .A2(G190), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n736), .B(new_n742), .C1(G68), .C2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(G20), .B1(new_n739), .B2(G179), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT91), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G97), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n724), .A2(new_n717), .A3(new_n725), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n732), .A2(new_n744), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT92), .Z(new_n754));
  INV_X1    g0554(.A(new_n743), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT33), .B(G317), .Z(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n741), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT94), .Z(new_n759));
  INV_X1    g0559(.A(new_n731), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  INV_X1    g0561(.A(G294), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n749), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n765));
  INV_X1    g0565(.A(new_n737), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n370), .B1(new_n766), .B2(G311), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n767), .B1(new_n768), .B2(new_n735), .C1(new_n583), .C2(new_n734), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G329), .B2(new_n724), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n764), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n754), .B1(new_n759), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n716), .B1(new_n772), .B2(new_n713), .ZN(new_n773));
  INV_X1    g0573(.A(new_n712), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n648), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n649), .A2(new_n702), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G330), .B2(new_n648), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n444), .A2(new_n644), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n633), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n666), .ZN(new_n783));
  INV_X1    g0583(.A(new_n440), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n644), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n441), .A2(new_n442), .B1(new_n439), .B2(new_n643), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n782), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n684), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n702), .B1(new_n789), .B2(new_n684), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n710), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n713), .A2(new_n710), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n702), .B1(G77), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n751), .B1(new_n755), .B2(new_n768), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n273), .B1(new_n741), .B2(new_n762), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G116), .B2(new_n766), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n735), .A2(new_n733), .ZN(new_n800));
  INV_X1    g0600(.A(new_n734), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(G107), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n799), .B(new_n802), .C1(new_n803), .C2(new_n723), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n797), .B(new_n804), .C1(G303), .C2(new_n731), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT95), .B(G143), .Z(new_n806));
  AOI22_X1  g0606(.A1(new_n740), .A2(new_n806), .B1(new_n766), .B2(new_n725), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n755), .B2(new_n378), .C1(new_n808), .C2(new_n760), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT34), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n749), .A2(new_n202), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n735), .A2(new_n213), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G50), .B2(new_n801), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT96), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n370), .B1(new_n813), .B2(new_n814), .C1(new_n815), .C2(new_n723), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n811), .B(new_n816), .C1(new_n814), .C2(new_n813), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n805), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n796), .B1(new_n819), .B2(new_n713), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G384));
  INV_X1    g0622(.A(new_n508), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n823), .A2(KEYINPUT35), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(KEYINPUT35), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n824), .A2(G116), .A3(new_n229), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT36), .Z(new_n827));
  OAI211_X1 g0627(.A(new_n231), .B(G77), .C1(new_n202), .C2(new_n213), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n201), .A2(G68), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n292), .B(G13), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n256), .B1(new_n270), .B2(new_n276), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT16), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n353), .B1(new_n834), .B2(new_n360), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n640), .A2(new_n642), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n350), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n339), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT37), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT97), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(KEYINPUT97), .B(KEYINPUT37), .C1(new_n837), .C2(new_n838), .ZN(new_n842));
  INV_X1    g0642(.A(new_n836), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n257), .B1(new_n357), .B2(new_n358), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n844), .A2(new_n282), .A3(new_n286), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n353), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n341), .A2(new_n846), .A3(new_n847), .A4(new_n350), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n841), .A2(new_n842), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n835), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n363), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n851), .A3(KEYINPUT38), .ZN(new_n852));
  INV_X1    g0652(.A(new_n846), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n363), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n341), .A2(new_n350), .A3(new_n846), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n848), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n849), .A2(new_n851), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n859), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(KEYINPUT39), .A3(new_n852), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n424), .A2(new_n417), .A3(new_n644), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n614), .A2(new_n843), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n852), .ZN(new_n871));
  INV_X1    g0671(.A(new_n418), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n643), .A2(new_n417), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n608), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n417), .B(new_n643), .C1(new_n424), .C2(new_n418), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n782), .B2(new_n785), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n870), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n869), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n617), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n667), .A2(new_n692), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(new_n445), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n879), .B(new_n882), .Z(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT98), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n679), .B2(new_n680), .ZN(new_n886));
  AOI211_X1 g0686(.A(KEYINPUT98), .B(KEYINPUT31), .C1(new_n678), .C2(new_n643), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n668), .A2(new_n888), .A3(new_n682), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n787), .B1(new_n874), .B2(new_n875), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n884), .B1(new_n861), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(new_n890), .A3(new_n884), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n865), .B2(new_n852), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n445), .A2(new_n889), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n897), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(G330), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n883), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n292), .B2(new_n699), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n883), .A2(new_n900), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n831), .B1(new_n902), .B2(new_n903), .ZN(G367));
  INV_X1    g0704(.A(new_n715), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n905), .B1(new_n224), .B2(new_n436), .C1(new_n243), .C2(new_n707), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n907), .A2(new_n702), .A3(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n644), .A2(new_n470), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n477), .A3(new_n624), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT99), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n910), .A2(new_n477), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT46), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n734), .B2(new_n588), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n917), .B(new_n919), .C1(new_n755), .C2(new_n762), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT109), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(KEYINPUT109), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n370), .B1(new_n740), .B2(G303), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n923), .B1(new_n205), .B2(new_n735), .C1(new_n768), .C2(new_n737), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(G317), .B2(new_n724), .ZN(new_n925));
  AOI22_X1  g0725(.A1(G311), .A2(new_n731), .B1(new_n750), .B2(G107), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n921), .A2(new_n922), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT110), .ZN(new_n928));
  AOI22_X1  g0728(.A1(G150), .A2(new_n740), .B1(new_n766), .B2(G50), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n202), .B2(new_n734), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n723), .A2(new_n808), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(new_n731), .C2(new_n806), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n370), .B1(new_n735), .B2(new_n215), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT111), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n743), .A2(new_n725), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n750), .A2(G68), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n932), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT47), .Z(new_n939));
  INV_X1    g0739(.A(new_n713), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n909), .B1(new_n774), .B2(new_n916), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n643), .A2(new_n515), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n526), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n644), .A2(new_n516), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n945), .A2(new_n571), .A3(new_n577), .A4(new_n653), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n946), .A2(KEYINPUT102), .A3(KEYINPUT42), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT102), .B1(new_n946), .B2(KEYINPUT42), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n947), .A2(new_n948), .B1(KEYINPUT42), .B2(new_n946), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n945), .B(KEYINPUT101), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n571), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n644), .B1(new_n951), .B2(new_n618), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n949), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT103), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n950), .A2(new_n652), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT104), .Z(new_n960));
  INV_X1    g0760(.A(KEYINPUT105), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n955), .B1(KEYINPUT43), .B2(new_n916), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n949), .A2(new_n952), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n960), .A2(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n960), .A2(new_n961), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n958), .A2(new_n964), .A3(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n654), .B1(new_n651), .B2(new_n653), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n649), .B(new_n971), .Z(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n694), .B2(new_n696), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n657), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT45), .ZN(new_n975));
  INV_X1    g0775(.A(new_n945), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n975), .B1(new_n976), .B2(new_n656), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT106), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n656), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n974), .A2(new_n977), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n983), .A2(new_n652), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n652), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT107), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n973), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n973), .B2(new_n987), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n697), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n660), .B(KEYINPUT41), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n701), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n941), .B1(new_n970), .B2(new_n995), .ZN(G387));
  INV_X1    g0796(.A(new_n972), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n697), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n660), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n694), .A2(new_n696), .A3(new_n972), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n651), .A2(new_n774), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n703), .A2(new_n662), .B1(G107), .B2(new_n224), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n239), .A2(new_n451), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n662), .ZN(new_n1007));
  AOI211_X1 g0807(.A(G45), .B(new_n1007), .C1(G68), .C2(G77), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n298), .A2(G50), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n707), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1005), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n702), .B1(new_n1012), .B2(new_n715), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n723), .A2(new_n378), .B1(new_n215), .B2(new_n734), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT112), .Z(new_n1015));
  NOR2_X1   g0815(.A1(new_n735), .A2(new_n205), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n370), .B1(new_n213), .B2(new_n737), .C1(new_n741), .C2(new_n201), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n474), .C2(new_n750), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G159), .A2(new_n731), .B1(new_n743), .B2(new_n299), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1015), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n749), .A2(new_n768), .B1(new_n762), .B2(new_n734), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G317), .A2(new_n740), .B1(new_n766), .B2(G303), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n755), .B2(new_n803), .C1(new_n757), .C2(new_n760), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT49), .Z(new_n1027));
  OAI221_X1 g0827(.A(new_n273), .B1(new_n588), .B2(new_n735), .C1(new_n723), .C2(new_n761), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1013), .B1(new_n1029), .B2(new_n713), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n997), .A2(new_n701), .B1(new_n1004), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1003), .A2(new_n1031), .ZN(G393));
  OAI21_X1  g0832(.A(new_n905), .B1(new_n205), .B2(new_n224), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n250), .A2(new_n707), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n702), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT114), .Z(new_n1036));
  AOI22_X1  g0836(.A1(new_n731), .A2(G317), .B1(G311), .B2(new_n740), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT52), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G303), .A2(new_n743), .B1(new_n750), .B2(G116), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n735), .A2(new_n206), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n273), .B1(new_n737), .B2(new_n762), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G283), .C2(new_n801), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n757), .C2(new_n723), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n731), .A2(G150), .B1(G159), .B2(new_n740), .ZN(new_n1044));
  XOR2_X1   g0844(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n724), .A2(new_n806), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n743), .A2(G50), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n370), .B1(new_n737), .B2(new_n298), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n800), .B(new_n1049), .C1(G68), .C2(new_n801), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n750), .A2(G77), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1038), .A2(new_n1043), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1036), .B1(new_n713), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n950), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n774), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n987), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n700), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n973), .A2(new_n987), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT107), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n989), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n661), .B1(new_n1057), .B2(new_n998), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(G390));
  AOI21_X1  g0864(.A(KEYINPUT38), .B1(new_n854), .B2(new_n857), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n850), .A2(new_n843), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n614), .B2(new_n610), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n341), .A2(new_n350), .A3(new_n846), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n839), .A2(new_n840), .B1(new_n1068), .B2(new_n847), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1069), .B2(new_n842), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1065), .B1(new_n1070), .B2(KEYINPUT38), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n868), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n874), .A2(new_n875), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n784), .A2(new_n786), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n691), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n785), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1072), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n683), .A2(G330), .A3(new_n788), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1073), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT39), .B1(new_n852), .B2(new_n860), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n849), .A2(KEYINPUT38), .A3(new_n851), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT38), .B1(new_n849), .B2(new_n851), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1082), .B1(new_n1085), .B2(KEYINPUT39), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT116), .B1(new_n877), .B2(new_n868), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT116), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1076), .B1(new_n633), .B2(new_n781), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1088), .B(new_n867), .C1(new_n1089), .C2(new_n876), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1078), .B(new_n1081), .C1(new_n1086), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1090), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n477), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n577), .A2(new_n624), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n525), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n1096), .B2(new_n630), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n780), .B1(new_n1097), .B2(new_n627), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1073), .B1(new_n1098), .B2(new_n1076), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1088), .B1(new_n1099), .B2(new_n867), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1093), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n863), .A2(new_n866), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1101), .A2(new_n1102), .B1(new_n1077), .B2(new_n1072), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n889), .A2(new_n890), .A3(G330), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n692), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n666), .A2(KEYINPUT29), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n445), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n445), .A2(G330), .A3(new_n889), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n617), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1104), .B1(new_n1080), .B2(new_n1073), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1089), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n889), .A2(G330), .A3(new_n788), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n876), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1081), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1110), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n661), .B1(new_n1105), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1092), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n702), .B1(new_n299), .B2(new_n795), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n737), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n370), .B1(new_n741), .B2(new_n815), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n735), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1126), .C1(G50), .C2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G128), .A2(new_n731), .B1(new_n750), .B2(G159), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n808), .C2(new_n755), .ZN(new_n1130));
  OR3_X1    g0930(.A1(new_n734), .A2(KEYINPUT53), .A3(new_n378), .ZN(new_n1131));
  OAI21_X1  g0931(.A(KEYINPUT53), .B1(new_n734), .B2(new_n378), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1132), .C1(new_n723), .C2(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G107), .A2(new_n743), .B1(new_n731), .B2(G283), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n737), .A2(new_n205), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1136), .B(new_n812), .C1(G116), .C2(new_n740), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n724), .A2(G294), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1051), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n273), .B1(new_n734), .B2(new_n733), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1130), .A2(new_n1134), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1123), .B1(new_n1142), .B2(new_n713), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1086), .B2(new_n711), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n1105), .B2(new_n700), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1122), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  INV_X1    g0947(.A(KEYINPUT122), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n836), .A2(new_n384), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n393), .B(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1150), .B(new_n1151), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(G330), .B1(new_n893), .B2(new_n895), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(new_n869), .B2(new_n878), .ZN(new_n1155));
  INV_X1    g0955(.A(G330), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT40), .B1(new_n1071), .B2(new_n891), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n894), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1156), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n879), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1153), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n879), .A2(new_n1160), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1154), .A2(new_n869), .A3(new_n878), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1164), .A3(new_n1152), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1110), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1162), .A2(new_n1165), .B1(new_n1166), .B2(new_n1121), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1148), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n661), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1163), .A2(new_n1164), .A3(new_n1152), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1152), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1121), .A2(new_n1166), .ZN(new_n1174));
  OAI211_X1 g0974(.A(KEYINPUT122), .B(new_n1170), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1168), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1152), .A2(new_n710), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n702), .B1(G50), .B2(new_n795), .ZN(new_n1178));
  INV_X1    g0978(.A(G41), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G50), .B1(new_n260), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n370), .B2(G41), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n205), .A2(new_n755), .B1(new_n760), .B2(new_n588), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n724), .A2(G283), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1127), .A2(G58), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G107), .A2(new_n740), .B1(new_n766), .B2(new_n474), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1183), .A2(new_n936), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1179), .B(new_n273), .C1(new_n734), .C2(new_n215), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT118), .Z(new_n1188));
  NOR3_X1   g0988(.A1(new_n1182), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G128), .A2(new_n740), .B1(new_n766), .B2(G137), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n734), .B2(new_n1124), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n760), .A2(new_n1133), .B1(new_n378), .B2(new_n749), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT120), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(G132), .C2(new_n743), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT59), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n724), .A2(G124), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n1127), .C2(new_n725), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1181), .B(new_n1191), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n940), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1178), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1177), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1173), .B2(new_n700), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1176), .A2(new_n1210), .ZN(G375));
  NAND2_X1  g1011(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n701), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n702), .B1(G68), .B2(new_n795), .ZN(new_n1214));
  INV_X1    g1014(.A(G159), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1184), .B1(new_n1215), .B2(new_n734), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n370), .B1(new_n378), .B2(new_n737), .C1(new_n741), .C2(new_n808), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G128), .C2(new_n724), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G132), .A2(new_n731), .B1(new_n750), .B2(G50), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n755), .C2(new_n1124), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n723), .A2(new_n583), .B1(new_n205), .B2(new_n734), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT123), .Z(new_n1222));
  AOI22_X1  g1022(.A1(G116), .A2(new_n743), .B1(new_n731), .B2(G294), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n273), .B1(new_n206), .B2(new_n737), .C1(new_n741), .C2(new_n768), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G77), .B2(new_n1127), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(new_n436), .C2(new_n749), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1220), .B1(new_n1222), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1214), .B1(new_n1227), .B2(new_n713), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1073), .B2(new_n711), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1213), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1212), .A2(new_n1166), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1119), .A2(new_n994), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1231), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  NAND3_X1  g1034(.A1(new_n1003), .A2(new_n778), .A3(new_n1031), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G378), .A2(G384), .A3(new_n1235), .A4(G381), .ZN(new_n1236));
  INV_X1    g1036(.A(G375), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n941), .B(new_n1063), .C1(new_n970), .C2(new_n995), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .ZN(G407));
  NOR2_X1   g1040(.A1(new_n641), .A2(G343), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1237), .A2(new_n1146), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(new_n1242), .A3(G213), .ZN(G409));
  NAND2_X1  g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1235), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT125), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1238), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n993), .B1(new_n1061), .B2(new_n697), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n968), .B(new_n969), .C1(new_n1249), .C2(new_n701), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1063), .B1(new_n1250), .B2(new_n941), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1246), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1253), .A2(new_n1245), .A3(new_n1247), .A4(new_n1238), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1176), .A2(G378), .A3(new_n1210), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1173), .A2(new_n1174), .A3(new_n993), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1146), .B1(new_n1257), .B2(new_n1209), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1241), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1232), .A2(KEYINPUT60), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1118), .A2(new_n661), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1232), .A2(KEYINPUT60), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1232), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1263), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1269), .B2(new_n1231), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n821), .B(new_n1230), .C1(new_n1263), .C2(new_n1268), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1259), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1255), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1272), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1241), .A2(G2897), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1262), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n821), .B1(new_n1281), .B2(new_n1230), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1269), .A2(G384), .A3(new_n1231), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1283), .A3(new_n1278), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1277), .B1(new_n1259), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1275), .A2(new_n1276), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1259), .A2(new_n1289), .A3(new_n1272), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1259), .B2(new_n1272), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1290), .A2(new_n1286), .A3(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1255), .B(KEYINPUT126), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1288), .B1(new_n1292), .B2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(new_n1272), .A2(KEYINPUT127), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1252), .A2(new_n1295), .A3(new_n1254), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1295), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1237), .A2(G378), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1256), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n1299), .A2(new_n1300), .B1(KEYINPUT127), .B2(new_n1272), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1298), .B(new_n1301), .ZN(G402));
endmodule


