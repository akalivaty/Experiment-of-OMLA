

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779;

  AND2_X1 U373 ( .A1(n621), .A2(n620), .ZN(n767) );
  NOR2_X1 U374 ( .A1(n640), .A2(n630), .ZN(n631) );
  INV_X2 U375 ( .A(KEYINPUT4), .ZN(n456) );
  XNOR2_X1 U376 ( .A(n631), .B(n632), .ZN(n648) );
  NOR2_X1 U377 ( .A1(n613), .A2(n684), .ZN(n380) );
  NOR2_X2 U378 ( .A1(n460), .A2(n751), .ZN(n665) );
  NOR2_X2 U379 ( .A1(n739), .A2(n751), .ZN(n740) );
  XNOR2_X2 U380 ( .A(n469), .B(KEYINPUT35), .ZN(n776) );
  OR2_X2 U381 ( .A1(n649), .A2(n459), .ZN(n589) );
  NOR2_X2 U382 ( .A1(n464), .A2(n751), .ZN(n445) );
  INV_X2 U383 ( .A(n649), .ZN(n351) );
  XNOR2_X1 U384 ( .A(n371), .B(n370), .ZN(n590) );
  XNOR2_X1 U385 ( .A(n397), .B(n586), .ZN(n605) );
  INV_X2 U386 ( .A(G128), .ZN(n513) );
  NOR2_X1 U387 ( .A1(n369), .A2(n704), .ZN(n638) );
  XNOR2_X1 U388 ( .A(n466), .B(n454), .ZN(n606) );
  INV_X1 U389 ( .A(KEYINPUT32), .ZN(n477) );
  XNOR2_X1 U390 ( .A(n436), .B(KEYINPUT65), .ZN(n354) );
  AND2_X1 U391 ( .A1(n427), .A2(n425), .ZN(n424) );
  AND2_X1 U392 ( .A1(n647), .A2(n666), .ZN(n406) );
  NAND2_X1 U393 ( .A1(n633), .A2(n707), .ZN(n666) );
  OR2_X1 U394 ( .A1(n592), .A2(n390), .ZN(n614) );
  AND2_X1 U395 ( .A1(n493), .A2(n490), .ZN(n489) );
  NAND2_X1 U396 ( .A1(n498), .A2(n495), .ZN(n707) );
  NOR2_X1 U397 ( .A1(n488), .A2(n487), .ZN(n486) );
  XNOR2_X1 U398 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U399 ( .A(n448), .B(KEYINPUT20), .ZN(n544) );
  XNOR2_X1 U400 ( .A(n522), .B(n359), .ZN(n387) );
  XNOR2_X1 U401 ( .A(n473), .B(n472), .ZN(n522) );
  XNOR2_X1 U402 ( .A(G110), .B(G104), .ZN(n473) );
  XNOR2_X1 U403 ( .A(G119), .B(KEYINPUT72), .ZN(n509) );
  XNOR2_X1 U404 ( .A(G902), .B(KEYINPUT15), .ZN(n656) );
  XNOR2_X2 U405 ( .A(n352), .B(n353), .ZN(n649) );
  NOR2_X1 U406 ( .A1(n661), .A2(G902), .ZN(n352) );
  XNOR2_X1 U407 ( .A(G472), .B(KEYINPUT100), .ZN(n353) );
  BUF_X1 U408 ( .A(n381), .Z(n355) );
  BUF_X1 U409 ( .A(n627), .Z(n356) );
  BUF_X1 U410 ( .A(n565), .Z(n357) );
  XNOR2_X1 U411 ( .A(n436), .B(KEYINPUT65), .ZN(n388) );
  NAND2_X2 U412 ( .A1(n434), .A2(n433), .ZN(n436) );
  NOR2_X1 U413 ( .A1(n623), .A2(n559), .ZN(n593) );
  INV_X1 U414 ( .A(KEYINPUT19), .ZN(n451) );
  AND2_X1 U415 ( .A1(n495), .A2(KEYINPUT68), .ZN(n494) );
  INV_X1 U416 ( .A(G469), .ZN(n370) );
  OR2_X1 U417 ( .A1(n736), .A2(G902), .ZN(n371) );
  AND2_X1 U418 ( .A1(n723), .A2(KEYINPUT2), .ZN(n726) );
  XNOR2_X1 U419 ( .A(n635), .B(KEYINPUT33), .ZN(n729) );
  XNOR2_X1 U420 ( .A(n518), .B(n455), .ZN(n385) );
  INV_X1 U421 ( .A(KEYINPUT80), .ZN(n455) );
  XNOR2_X1 U422 ( .A(n519), .B(n529), .ZN(n386) );
  XOR2_X1 U423 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n512) );
  NAND2_X1 U424 ( .A1(n489), .A2(n486), .ZN(n704) );
  NOR2_X1 U425 ( .A1(G953), .A2(G237), .ZN(n574) );
  NAND2_X1 U426 ( .A1(n776), .A2(KEYINPUT44), .ZN(n405) );
  NOR2_X1 U427 ( .A1(n409), .A2(n776), .ZN(n408) );
  INV_X1 U428 ( .A(KEYINPUT10), .ZN(n528) );
  XOR2_X1 U429 ( .A(G137), .B(G140), .Z(n530) );
  XOR2_X1 U430 ( .A(n607), .B(KEYINPUT38), .Z(n698) );
  AND2_X1 U431 ( .A1(n634), .A2(n361), .ZN(n591) );
  OR2_X1 U432 ( .A1(n744), .A2(G902), .ZN(n397) );
  INV_X1 U433 ( .A(KEYINPUT68), .ZN(n492) );
  NAND2_X1 U434 ( .A1(n708), .A2(n492), .ZN(n491) );
  NAND2_X1 U435 ( .A1(n483), .A2(n499), .ZN(n485) );
  NAND2_X1 U436 ( .A1(n500), .A2(G902), .ZN(n499) );
  INV_X1 U437 ( .A(n546), .ZN(n500) );
  NAND2_X1 U438 ( .A1(n546), .A2(n497), .ZN(n496) );
  INV_X1 U439 ( .A(G902), .ZN(n497) );
  NOR2_X1 U440 ( .A1(n590), .A2(n564), .ZN(n599) );
  XNOR2_X1 U441 ( .A(n566), .B(n481), .ZN(n480) );
  INV_X1 U442 ( .A(KEYINPUT83), .ZN(n481) );
  XNOR2_X1 U443 ( .A(KEYINPUT13), .B(G475), .ZN(n454) );
  OR2_X1 U444 ( .A1(n743), .A2(G902), .ZN(n466) );
  XNOR2_X1 U445 ( .A(n657), .B(n658), .ZN(n659) );
  INV_X1 U446 ( .A(G953), .ZN(n755) );
  NOR2_X1 U447 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U448 ( .A1(n731), .A2(n367), .ZN(n398) );
  XNOR2_X1 U449 ( .A(n641), .B(n365), .ZN(n374) );
  NOR2_X1 U450 ( .A1(n394), .A2(n422), .ZN(n421) );
  INV_X1 U451 ( .A(KEYINPUT75), .ZN(n423) );
  INV_X1 U452 ( .A(KEYINPUT87), .ZN(n468) );
  NOR2_X1 U453 ( .A1(n431), .A2(n430), .ZN(n429) );
  INV_X1 U454 ( .A(n779), .ZN(n415) );
  INV_X1 U455 ( .A(n374), .ZN(n372) );
  OR2_X1 U456 ( .A1(G902), .A2(G237), .ZN(n567) );
  XNOR2_X1 U457 ( .A(KEYINPUT21), .B(n527), .ZN(n628) );
  XNOR2_X1 U458 ( .A(n545), .B(KEYINPUT25), .ZN(n546) );
  XOR2_X1 U459 ( .A(KEYINPUT5), .B(G116), .Z(n547) );
  XNOR2_X1 U460 ( .A(KEYINPUT90), .B(KEYINPUT48), .ZN(n501) );
  INV_X1 U461 ( .A(G134), .ZN(n517) );
  XOR2_X1 U462 ( .A(KEYINPUT105), .B(G122), .Z(n569) );
  XNOR2_X1 U463 ( .A(G104), .B(G113), .ZN(n568) );
  XOR2_X1 U464 ( .A(G140), .B(G143), .Z(n503) );
  XNOR2_X1 U465 ( .A(KEYINPUT104), .B(KEYINPUT103), .ZN(n570) );
  XOR2_X1 U466 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n571) );
  NAND2_X1 U467 ( .A1(G237), .A2(G234), .ZN(n554) );
  NOR2_X1 U468 ( .A1(n707), .A2(n628), .ZN(n561) );
  XNOR2_X1 U469 ( .A(n752), .B(n382), .ZN(n565) );
  XNOR2_X1 U470 ( .A(n383), .B(n514), .ZN(n382) );
  XNOR2_X1 U471 ( .A(n385), .B(n386), .ZN(n383) );
  INV_X1 U472 ( .A(KEYINPUT30), .ZN(n443) );
  XOR2_X1 U473 ( .A(KEYINPUT24), .B(KEYINPUT99), .Z(n533) );
  XNOR2_X1 U474 ( .A(G119), .B(KEYINPUT73), .ZN(n532) );
  XNOR2_X1 U475 ( .A(KEYINPUT98), .B(KEYINPUT78), .ZN(n537) );
  XNOR2_X1 U476 ( .A(n575), .B(n531), .ZN(n764) );
  XOR2_X1 U477 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n536) );
  INV_X1 U478 ( .A(G475), .ZN(n399) );
  INV_X1 U479 ( .A(KEYINPUT96), .ZN(n472) );
  XNOR2_X1 U480 ( .A(n450), .B(n449), .ZN(n728) );
  INV_X1 U481 ( .A(KEYINPUT41), .ZN(n449) );
  NOR2_X1 U482 ( .A1(n695), .A2(n700), .ZN(n450) );
  XNOR2_X1 U483 ( .A(n462), .B(n461), .ZN(n613) );
  INV_X1 U484 ( .A(KEYINPUT39), .ZN(n461) );
  NAND2_X1 U485 ( .A1(n391), .A2(n594), .ZN(n390) );
  XNOR2_X1 U486 ( .A(n600), .B(KEYINPUT82), .ZN(n602) );
  INV_X1 U487 ( .A(n491), .ZN(n484) );
  XNOR2_X1 U488 ( .A(n661), .B(KEYINPUT62), .ZN(n663) );
  AND2_X2 U489 ( .A1(n388), .A2(n400), .ZN(n749) );
  XNOR2_X1 U490 ( .A(n636), .B(n471), .ZN(n470) );
  XNOR2_X1 U491 ( .A(KEYINPUT81), .B(KEYINPUT34), .ZN(n471) );
  NOR2_X1 U492 ( .A1(n610), .A2(n609), .ZN(n678) );
  INV_X1 U493 ( .A(n602), .ZN(n679) );
  INV_X1 U494 ( .A(KEYINPUT108), .ZN(n453) );
  OR2_X1 U495 ( .A1(n648), .A2(n463), .ZN(n650) );
  OR2_X1 U496 ( .A1(n651), .A2(n351), .ZN(n463) );
  INV_X1 U497 ( .A(KEYINPUT92), .ZN(n392) );
  INV_X1 U498 ( .A(KEYINPUT60), .ZN(n401) );
  NAND2_X1 U499 ( .A1(n659), .A2(n403), .ZN(n447) );
  AND2_X1 U500 ( .A1(n730), .A2(n398), .ZN(n732) );
  INV_X1 U501 ( .A(n684), .ZN(n373) );
  NOR2_X1 U502 ( .A1(n726), .A2(n399), .ZN(n358) );
  XNOR2_X1 U503 ( .A(KEYINPUT16), .B(KEYINPUT74), .ZN(n359) );
  XNOR2_X1 U504 ( .A(n590), .B(KEYINPUT1), .ZN(n369) );
  INV_X1 U505 ( .A(n697), .ZN(n459) );
  INV_X1 U506 ( .A(n707), .ZN(n391) );
  XNOR2_X1 U507 ( .A(KEYINPUT9), .B(KEYINPUT106), .ZN(n360) );
  AND2_X1 U508 ( .A1(n708), .A2(n697), .ZN(n361) );
  AND2_X1 U509 ( .A1(n486), .A2(n442), .ZN(n362) );
  INV_X1 U510 ( .A(n369), .ZN(n651) );
  AND2_X1 U511 ( .A1(n651), .A2(KEYINPUT91), .ZN(n363) );
  AND2_X1 U512 ( .A1(n362), .A2(n489), .ZN(n364) );
  XOR2_X1 U513 ( .A(KEYINPUT102), .B(KEYINPUT31), .Z(n365) );
  XOR2_X1 U514 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n366) );
  AND2_X1 U515 ( .A1(n729), .A2(n728), .ZN(n367) );
  XOR2_X1 U516 ( .A(n660), .B(KEYINPUT56), .Z(n368) );
  NOR2_X1 U517 ( .A1(n769), .A2(G952), .ZN(n751) );
  INV_X1 U518 ( .A(n751), .ZN(n403) );
  XNOR2_X2 U519 ( .A(n456), .B(G101), .ZN(n519) );
  NAND2_X1 U520 ( .A1(n372), .A2(n670), .ZN(n646) );
  AND2_X1 U521 ( .A1(n374), .A2(n373), .ZN(n685) );
  AND2_X1 U522 ( .A1(n374), .A2(n675), .ZN(n688) );
  NAND2_X1 U523 ( .A1(n376), .A2(n375), .ZN(n378) );
  NAND2_X1 U524 ( .A1(n476), .A2(n742), .ZN(n375) );
  NAND2_X1 U525 ( .A1(n475), .A2(n358), .ZN(n376) );
  NAND2_X1 U526 ( .A1(n377), .A2(n403), .ZN(n402) );
  XNOR2_X1 U527 ( .A(n378), .B(n404), .ZN(n377) );
  NAND2_X1 U528 ( .A1(n379), .A2(n415), .ZN(n414) );
  INV_X1 U529 ( .A(n778), .ZN(n379) );
  XNOR2_X1 U530 ( .A(n380), .B(KEYINPUT40), .ZN(n778) );
  NOR2_X2 U531 ( .A1(n381), .A2(KEYINPUT2), .ZN(n435) );
  AND2_X1 U532 ( .A1(n767), .A2(n381), .ZN(n723) );
  NAND2_X1 U533 ( .A1(n355), .A2(n755), .ZN(n756) );
  XNOR2_X2 U534 ( .A(n389), .B(KEYINPUT45), .ZN(n381) );
  XNOR2_X2 U535 ( .A(n387), .B(n384), .ZN(n752) );
  XNOR2_X2 U536 ( .A(n548), .B(n581), .ZN(n384) );
  XNOR2_X2 U537 ( .A(n504), .B(G122), .ZN(n581) );
  XNOR2_X2 U538 ( .A(n509), .B(n510), .ZN(n548) );
  NAND2_X1 U539 ( .A1(n358), .A2(n354), .ZN(n476) );
  AND2_X1 U540 ( .A1(n354), .A2(n741), .ZN(n475) );
  NOR2_X1 U541 ( .A1(n439), .A2(n438), .ZN(n437) );
  OR2_X2 U542 ( .A1(n767), .A2(KEYINPUT2), .ZN(n433) );
  XNOR2_X1 U543 ( .A(n414), .B(KEYINPUT46), .ZN(n413) );
  XNOR2_X1 U544 ( .A(n553), .B(n552), .ZN(n661) );
  NAND2_X2 U545 ( .A1(n652), .A2(n479), .ZN(n478) );
  NAND2_X1 U546 ( .A1(n395), .A2(n410), .ZN(n389) );
  NOR2_X1 U547 ( .A1(n416), .A2(n413), .ZN(n502) );
  NOR2_X2 U548 ( .A1(n707), .A2(n650), .ZN(n673) );
  NOR2_X1 U549 ( .A1(n408), .A2(n407), .ZN(n395) );
  NAND2_X1 U550 ( .A1(n429), .A2(n428), .ZN(n418) );
  XNOR2_X1 U551 ( .A(n393), .B(n392), .ZN(n633) );
  NAND2_X1 U552 ( .A1(n652), .A2(n369), .ZN(n393) );
  NAND2_X1 U553 ( .A1(n470), .A2(n637), .ZN(n469) );
  XNOR2_X1 U554 ( .A(n411), .B(n655), .ZN(n410) );
  NOR2_X2 U555 ( .A1(n777), .A2(n673), .ZN(n654) );
  INV_X1 U556 ( .A(n394), .ZN(n432) );
  NAND2_X1 U557 ( .A1(n603), .A2(n604), .ZN(n394) );
  NAND2_X1 U558 ( .A1(n419), .A2(n424), .ZN(n417) );
  XNOR2_X2 U559 ( .A(n396), .B(n453), .ZN(n675) );
  NAND2_X1 U560 ( .A1(n596), .A2(n606), .ZN(n396) );
  XNOR2_X1 U561 ( .A(n696), .B(n468), .ZN(n644) );
  XNOR2_X1 U562 ( .A(n582), .B(n457), .ZN(n585) );
  INV_X1 U563 ( .A(n726), .ZN(n400) );
  XNOR2_X1 U564 ( .A(n402), .B(n401), .ZN(G60) );
  INV_X1 U565 ( .A(n743), .ZN(n404) );
  NOR2_X2 U566 ( .A1(n654), .A2(n653), .ZN(n411) );
  NAND2_X1 U567 ( .A1(n406), .A2(n405), .ZN(n407) );
  NAND2_X1 U568 ( .A1(n654), .A2(n653), .ZN(n409) );
  XNOR2_X2 U569 ( .A(n412), .B(n577), .ZN(n765) );
  XNOR2_X1 U570 ( .A(n412), .B(n360), .ZN(n457) );
  XNOR2_X2 U571 ( .A(n518), .B(n517), .ZN(n412) );
  NAND2_X1 U572 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U573 ( .A1(n421), .A2(n420), .ZN(n419) );
  INV_X1 U574 ( .A(n611), .ZN(n420) );
  NAND2_X1 U575 ( .A1(n612), .A2(n423), .ZN(n422) );
  NAND2_X1 U576 ( .A1(n426), .A2(KEYINPUT75), .ZN(n425) );
  NAND2_X1 U577 ( .A1(n432), .A2(n612), .ZN(n426) );
  NAND2_X1 U578 ( .A1(n611), .A2(KEYINPUT75), .ZN(n427) );
  AND2_X1 U579 ( .A1(n458), .A2(n651), .ZN(n690) );
  NAND2_X1 U580 ( .A1(n458), .A2(n363), .ZN(n428) );
  NOR2_X1 U581 ( .A1(n651), .A2(KEYINPUT91), .ZN(n430) );
  NOR2_X1 U582 ( .A1(n458), .A2(KEYINPUT91), .ZN(n431) );
  NOR2_X2 U583 ( .A1(n435), .A2(n656), .ZN(n434) );
  XNOR2_X1 U584 ( .A(n589), .B(n443), .ZN(n441) );
  NAND2_X1 U585 ( .A1(n441), .A2(n437), .ZN(n444) );
  INV_X1 U586 ( .A(n489), .ZN(n438) );
  NAND2_X1 U587 ( .A1(n440), .A2(n486), .ZN(n439) );
  NOR2_X1 U588 ( .A1(n590), .A2(n593), .ZN(n440) );
  INV_X1 U589 ( .A(n590), .ZN(n442) );
  XNOR2_X2 U590 ( .A(n444), .B(KEYINPUT77), .ZN(n608) );
  NAND2_X1 U591 ( .A1(n608), .A2(n698), .ZN(n462) );
  XNOR2_X1 U592 ( .A(n445), .B(KEYINPUT124), .ZN(G66) );
  NAND2_X1 U593 ( .A1(n565), .A2(n656), .ZN(n482) );
  INV_X2 U594 ( .A(n446), .ZN(n529) );
  XNOR2_X2 U595 ( .A(G146), .B(G125), .ZN(n446) );
  NOR2_X1 U596 ( .A1(n614), .A2(n617), .ZN(n595) );
  XNOR2_X1 U597 ( .A(n662), .B(n663), .ZN(n460) );
  XNOR2_X1 U598 ( .A(n750), .B(n748), .ZN(n464) );
  XNOR2_X1 U599 ( .A(n452), .B(n451), .ZN(n627) );
  XNOR2_X1 U600 ( .A(n447), .B(n368), .ZN(G51) );
  NAND2_X1 U601 ( .A1(n656), .A2(G234), .ZN(n448) );
  NOR2_X2 U602 ( .A1(n648), .A2(n634), .ZN(n652) );
  NOR2_X2 U603 ( .A1(n617), .A2(n459), .ZN(n452) );
  NOR2_X2 U604 ( .A1(n675), .A2(n680), .ZN(n696) );
  NOR2_X1 U605 ( .A1(n644), .A2(n597), .ZN(n598) );
  XOR2_X2 U606 ( .A(KEYINPUT71), .B(G131), .Z(n577) );
  XNOR2_X1 U607 ( .A(n578), .B(n576), .ZN(n467) );
  XNOR2_X1 U608 ( .A(n575), .B(n467), .ZN(n579) );
  XOR2_X2 U609 ( .A(n351), .B(KEYINPUT6), .Z(n634) );
  INV_X2 U610 ( .A(n557), .ZN(n769) );
  XNOR2_X1 U611 ( .A(n595), .B(KEYINPUT36), .ZN(n458) );
  XNOR2_X2 U612 ( .A(n765), .B(n520), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n749), .A2(G472), .ZN(n662) );
  NAND2_X1 U614 ( .A1(n465), .A2(n679), .ZN(n612) );
  XNOR2_X1 U615 ( .A(n598), .B(KEYINPUT76), .ZN(n465) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n621) );
  NAND2_X1 U617 ( .A1(n749), .A2(G217), .ZN(n750) );
  XNOR2_X2 U618 ( .A(n474), .B(n366), .ZN(n640) );
  NAND2_X1 U619 ( .A1(n627), .A2(n626), .ZN(n474) );
  XNOR2_X2 U620 ( .A(n478), .B(n477), .ZN(n777) );
  AND2_X1 U621 ( .A1(n651), .A2(n391), .ZN(n479) );
  XNOR2_X2 U622 ( .A(n482), .B(n480), .ZN(n617) );
  NAND2_X1 U623 ( .A1(n748), .A2(n500), .ZN(n483) );
  INV_X1 U624 ( .A(n485), .ZN(n498) );
  NAND2_X1 U625 ( .A1(n485), .A2(n484), .ZN(n490) );
  NOR2_X1 U626 ( .A1(n708), .A2(n492), .ZN(n487) );
  NOR2_X1 U627 ( .A1(n495), .A2(n491), .ZN(n488) );
  NAND2_X1 U628 ( .A1(n494), .A2(n498), .ZN(n493) );
  OR2_X1 U629 ( .A1(n748), .A2(n496), .ZN(n495) );
  XNOR2_X2 U630 ( .A(G953), .B(KEYINPUT64), .ZN(n557) );
  XNOR2_X1 U631 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U632 ( .A(n547), .B(G137), .ZN(n549) );
  NAND2_X1 U633 ( .A1(n629), .A2(n708), .ZN(n630) );
  XNOR2_X1 U634 ( .A(n548), .B(n549), .ZN(n550) );
  XNOR2_X1 U635 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U636 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U637 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n562) );
  XNOR2_X1 U638 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U639 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U640 ( .A(KEYINPUT63), .B(KEYINPUT95), .ZN(n664) );
  XNOR2_X1 U641 ( .A(n665), .B(n664), .ZN(G57) );
  XNOR2_X1 U642 ( .A(KEYINPUT55), .B(KEYINPUT93), .ZN(n516) );
  XNOR2_X2 U643 ( .A(G107), .B(G116), .ZN(n504) );
  INV_X1 U644 ( .A(KEYINPUT3), .ZN(n505) );
  NAND2_X1 U645 ( .A1(G113), .A2(n505), .ZN(n508) );
  INV_X1 U646 ( .A(G113), .ZN(n506) );
  NAND2_X1 U647 ( .A1(n506), .A2(KEYINPUT3), .ZN(n507) );
  NAND2_X1 U648 ( .A1(n508), .A2(n507), .ZN(n510) );
  NAND2_X1 U649 ( .A1(G224), .A2(n769), .ZN(n511) );
  XNOR2_X1 U650 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X2 U651 ( .A(n513), .B(G143), .ZN(n518) );
  XNOR2_X1 U652 ( .A(n357), .B(KEYINPUT54), .ZN(n515) );
  XNOR2_X1 U653 ( .A(n516), .B(n515), .ZN(n658) );
  XOR2_X1 U654 ( .A(G146), .B(n519), .Z(n520) );
  XNOR2_X1 U655 ( .A(n530), .B(KEYINPUT79), .ZN(n521) );
  XNOR2_X1 U656 ( .A(n521), .B(G107), .ZN(n525) );
  NAND2_X1 U657 ( .A1(G227), .A2(n769), .ZN(n523) );
  XNOR2_X1 U658 ( .A(n553), .B(n526), .ZN(n736) );
  NAND2_X1 U659 ( .A1(n544), .A2(G221), .ZN(n527) );
  XNOR2_X2 U660 ( .A(n529), .B(n528), .ZN(n575) );
  INV_X1 U661 ( .A(n530), .ZN(n531) );
  XNOR2_X1 U662 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U663 ( .A(n764), .B(n534), .ZN(n543) );
  NAND2_X1 U664 ( .A1(G234), .A2(n769), .ZN(n535) );
  XNOR2_X1 U665 ( .A(n536), .B(n535), .ZN(n583) );
  AND2_X1 U666 ( .A1(n583), .A2(G221), .ZN(n541) );
  XOR2_X1 U667 ( .A(G110), .B(G128), .Z(n538) );
  XNOR2_X1 U668 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U669 ( .A(n539), .B(KEYINPUT23), .Z(n540) );
  XNOR2_X1 U670 ( .A(n542), .B(n543), .ZN(n748) );
  NAND2_X1 U671 ( .A1(n544), .A2(G217), .ZN(n545) );
  NAND2_X1 U672 ( .A1(G210), .A2(n574), .ZN(n551) );
  XNOR2_X1 U673 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U674 ( .A(n554), .B(KEYINPUT14), .ZN(n556) );
  NAND2_X1 U675 ( .A1(n556), .A2(G952), .ZN(n555) );
  XOR2_X1 U676 ( .A(KEYINPUT97), .B(n555), .Z(n721) );
  NOR2_X1 U677 ( .A1(G953), .A2(n721), .ZN(n623) );
  AND2_X1 U678 ( .A1(G902), .A2(n556), .ZN(n622) );
  NAND2_X1 U679 ( .A1(n622), .A2(n557), .ZN(n558) );
  NOR2_X1 U680 ( .A1(G900), .A2(n558), .ZN(n559) );
  NOR2_X1 U681 ( .A1(n649), .A2(n593), .ZN(n560) );
  NAND2_X1 U682 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U683 ( .A1(n567), .A2(G210), .ZN(n566) );
  INV_X1 U684 ( .A(n617), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G214), .A2(n567), .ZN(n697) );
  NAND2_X1 U686 ( .A1(n698), .A2(n697), .ZN(n695) );
  XNOR2_X1 U687 ( .A(n569), .B(n568), .ZN(n573) );
  XNOR2_X1 U688 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U689 ( .A(n573), .B(n572), .ZN(n580) );
  NAND2_X1 U690 ( .A1(G214), .A2(n574), .ZN(n576) );
  XNOR2_X1 U691 ( .A(n577), .B(n503), .ZN(n578) );
  XNOR2_X1 U692 ( .A(n580), .B(n579), .ZN(n743) );
  XNOR2_X1 U693 ( .A(KEYINPUT107), .B(G478), .ZN(n586) );
  XNOR2_X1 U694 ( .A(n581), .B(KEYINPUT7), .ZN(n582) );
  NAND2_X1 U695 ( .A1(G217), .A2(n583), .ZN(n584) );
  XNOR2_X1 U696 ( .A(n585), .B(n584), .ZN(n744) );
  NAND2_X1 U697 ( .A1(n606), .A2(n605), .ZN(n700) );
  NAND2_X1 U698 ( .A1(n599), .A2(n728), .ZN(n588) );
  XNOR2_X1 U699 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n587) );
  XNOR2_X1 U700 ( .A(n588), .B(n587), .ZN(n779) );
  INV_X1 U701 ( .A(n628), .ZN(n708) );
  INV_X1 U702 ( .A(n605), .ZN(n596) );
  NOR2_X1 U703 ( .A1(n596), .A2(n606), .ZN(n680) );
  INV_X1 U704 ( .A(n680), .ZN(n684) );
  NAND2_X1 U705 ( .A1(n680), .A2(n591), .ZN(n592) );
  INV_X1 U706 ( .A(n593), .ZN(n594) );
  XOR2_X1 U707 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n597) );
  NAND2_X1 U708 ( .A1(n599), .A2(n356), .ZN(n600) );
  NAND2_X1 U709 ( .A1(n696), .A2(KEYINPUT47), .ZN(n601) );
  XNOR2_X1 U710 ( .A(n601), .B(KEYINPUT86), .ZN(n604) );
  NAND2_X1 U711 ( .A1(n602), .A2(KEYINPUT47), .ZN(n603) );
  NOR2_X1 U712 ( .A1(n606), .A2(n605), .ZN(n637) );
  INV_X1 U713 ( .A(n637), .ZN(n610) );
  NAND2_X1 U714 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U715 ( .A(n678), .B(KEYINPUT88), .ZN(n611) );
  INV_X1 U716 ( .A(n675), .ZN(n687) );
  NOR2_X1 U717 ( .A1(n687), .A2(n613), .ZN(n693) );
  NOR2_X1 U718 ( .A1(n651), .A2(n614), .ZN(n616) );
  XNOR2_X1 U719 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n615) );
  XNOR2_X1 U720 ( .A(n616), .B(n615), .ZN(n618) );
  NAND2_X1 U721 ( .A1(n618), .A2(n617), .ZN(n694) );
  INV_X1 U722 ( .A(n694), .ZN(n619) );
  NOR2_X1 U723 ( .A1(n693), .A2(n619), .ZN(n620) );
  INV_X1 U724 ( .A(KEYINPUT22), .ZN(n632) );
  NOR2_X1 U725 ( .A1(G898), .A2(n755), .ZN(n754) );
  NAND2_X1 U726 ( .A1(n754), .A2(n622), .ZN(n625) );
  INV_X1 U727 ( .A(n623), .ZN(n624) );
  NAND2_X1 U728 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U729 ( .A(n700), .ZN(n629) );
  NAND2_X1 U730 ( .A1(n638), .A2(n634), .ZN(n635) );
  INV_X1 U731 ( .A(n640), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n729), .A2(n642), .ZN(n636) );
  AND2_X1 U733 ( .A1(n638), .A2(n351), .ZN(n639) );
  XNOR2_X1 U734 ( .A(n639), .B(KEYINPUT101), .ZN(n713) );
  NOR2_X1 U735 ( .A1(n640), .A2(n713), .ZN(n641) );
  AND2_X1 U736 ( .A1(n642), .A2(n364), .ZN(n643) );
  NAND2_X1 U737 ( .A1(n649), .A2(n643), .ZN(n670) );
  INV_X1 U738 ( .A(n644), .ZN(n645) );
  NAND2_X1 U739 ( .A1(n646), .A2(n645), .ZN(n647) );
  INV_X1 U740 ( .A(KEYINPUT44), .ZN(n653) );
  INV_X1 U741 ( .A(KEYINPUT66), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n749), .A2(G210), .ZN(n657) );
  INV_X1 U743 ( .A(KEYINPUT121), .ZN(n660) );
  XNOR2_X1 U744 ( .A(G101), .B(n666), .ZN(G3) );
  NOR2_X1 U745 ( .A1(n684), .A2(n670), .ZN(n667) );
  XOR2_X1 U746 ( .A(G104), .B(n667), .Z(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n669) );
  XNOR2_X1 U748 ( .A(G107), .B(KEYINPUT27), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n672) );
  NOR2_X1 U750 ( .A1(n687), .A2(n670), .ZN(n671) );
  XOR2_X1 U751 ( .A(n672), .B(n671), .Z(G9) );
  XNOR2_X1 U752 ( .A(G110), .B(n673), .ZN(n674) );
  XNOR2_X1 U753 ( .A(n674), .B(KEYINPUT113), .ZN(G12) );
  XOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .Z(n677) );
  NAND2_X1 U755 ( .A1(n675), .A2(n679), .ZN(n676) );
  XNOR2_X1 U756 ( .A(n677), .B(n676), .ZN(G30) );
  XOR2_X1 U757 ( .A(n678), .B(G143), .Z(G45) );
  XOR2_X1 U758 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n682) );
  NAND2_X1 U759 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U760 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U761 ( .A(G146), .B(n683), .ZN(G48) );
  XOR2_X1 U762 ( .A(KEYINPUT116), .B(n685), .Z(n686) );
  XNOR2_X1 U763 ( .A(G113), .B(n686), .ZN(G15) );
  XNOR2_X1 U764 ( .A(G116), .B(KEYINPUT117), .ZN(n689) );
  XNOR2_X1 U765 ( .A(n689), .B(n688), .ZN(G18) );
  XNOR2_X1 U766 ( .A(n690), .B(KEYINPUT118), .ZN(n691) );
  XNOR2_X1 U767 ( .A(n691), .B(KEYINPUT37), .ZN(n692) );
  XNOR2_X1 U768 ( .A(G125), .B(n692), .ZN(G27) );
  XOR2_X1 U769 ( .A(G134), .B(n693), .Z(G36) );
  XNOR2_X1 U770 ( .A(G140), .B(n694), .ZN(G42) );
  XOR2_X1 U771 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n734) );
  NOR2_X1 U772 ( .A1(n696), .A2(n695), .ZN(n702) );
  NOR2_X1 U773 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U774 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U776 ( .A1(n729), .A2(n703), .ZN(n718) );
  NAND2_X1 U777 ( .A1(n369), .A2(n704), .ZN(n705) );
  XOR2_X1 U778 ( .A(KEYINPUT50), .B(n705), .Z(n706) );
  XNOR2_X1 U779 ( .A(n706), .B(KEYINPUT119), .ZN(n712) );
  NOR2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U781 ( .A(KEYINPUT49), .B(n709), .Z(n710) );
  NOR2_X1 U782 ( .A1(n351), .A2(n710), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U785 ( .A(KEYINPUT51), .B(n715), .Z(n716) );
  NAND2_X1 U786 ( .A1(n728), .A2(n716), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U788 ( .A(KEYINPUT52), .B(n719), .Z(n720) );
  NOR2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n731) );
  XOR2_X1 U790 ( .A(KEYINPUT85), .B(KEYINPUT2), .Z(n722) );
  NOR2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U792 ( .A(n724), .B(KEYINPUT84), .ZN(n725) );
  XNOR2_X1 U793 ( .A(n727), .B(KEYINPUT89), .ZN(n730) );
  NAND2_X1 U794 ( .A1(n732), .A2(n755), .ZN(n733) );
  XNOR2_X1 U795 ( .A(n734), .B(n733), .ZN(G75) );
  NAND2_X1 U796 ( .A1(n749), .A2(G469), .ZN(n738) );
  XOR2_X1 U797 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n735) );
  XNOR2_X1 U798 ( .A(n740), .B(KEYINPUT122), .ZN(G54) );
  XOR2_X1 U799 ( .A(KEYINPUT59), .B(KEYINPUT94), .Z(n742) );
  INV_X1 U800 ( .A(n742), .ZN(n741) );
  XOR2_X1 U801 ( .A(n744), .B(KEYINPUT123), .Z(n746) );
  NAND2_X1 U802 ( .A1(n749), .A2(G478), .ZN(n745) );
  XNOR2_X1 U803 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U804 ( .A1(n751), .A2(n747), .ZN(G63) );
  XNOR2_X1 U805 ( .A(n752), .B(G101), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n763) );
  XNOR2_X1 U807 ( .A(n756), .B(KEYINPUT126), .ZN(n761) );
  XOR2_X1 U808 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n758) );
  NAND2_X1 U809 ( .A1(G224), .A2(G953), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U811 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(G69) );
  XNOR2_X1 U814 ( .A(n764), .B(KEYINPUT4), .ZN(n766) );
  XOR2_X1 U815 ( .A(n765), .B(n766), .Z(n771) );
  BUF_X1 U816 ( .A(n767), .Z(n768) );
  XOR2_X1 U817 ( .A(n771), .B(n768), .Z(n770) );
  NAND2_X1 U818 ( .A1(n770), .A2(n769), .ZN(n775) );
  XNOR2_X1 U819 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n775), .A2(n774), .ZN(G72) );
  XOR2_X1 U823 ( .A(G122), .B(n776), .Z(G24) );
  XOR2_X1 U824 ( .A(n777), .B(G119), .Z(G21) );
  XOR2_X1 U825 ( .A(n778), .B(G131), .Z(G33) );
  XOR2_X1 U826 ( .A(n779), .B(G137), .Z(G39) );
endmodule

