

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U549 ( .A1(n830), .A2(n829), .ZN(n832) );
  AND2_X2 U550 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U551 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  INV_X1 U552 ( .A(KEYINPUT28), .ZN(n714) );
  OR2_X1 U553 ( .A1(n757), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U554 ( .A1(n760), .A2(n759), .ZN(n761) );
  INV_X1 U555 ( .A(n987), .ZN(n759) );
  XOR2_X1 U556 ( .A(KEYINPUT1), .B(n521), .Z(n650) );
  INV_X1 U557 ( .A(n736), .ZN(n708) );
  XNOR2_X1 U558 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n725) );
  XNOR2_X1 U559 ( .A(n726), .B(n725), .ZN(n727) );
  INV_X1 U560 ( .A(KEYINPUT29), .ZN(n718) );
  XNOR2_X1 U561 ( .A(n719), .B(n718), .ZN(n723) );
  AND2_X1 U562 ( .A1(G160), .A2(G40), .ZN(n687) );
  NAND2_X1 U563 ( .A1(n736), .A2(G8), .ZN(n774) );
  INV_X1 U564 ( .A(KEYINPUT17), .ZN(n533) );
  NAND2_X1 U565 ( .A1(n885), .A2(G137), .ZN(n535) );
  OR2_X1 U566 ( .A1(n520), .A2(n641), .ZN(n515) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U568 ( .A1(n649), .A2(G89), .ZN(n514) );
  XNOR2_X1 U569 ( .A(KEYINPUT4), .B(n514), .ZN(n518) );
  INV_X1 U570 ( .A(G651), .ZN(n520) );
  XOR2_X2 U571 ( .A(KEYINPUT68), .B(n515), .Z(n656) );
  NAND2_X1 U572 ( .A1(G76), .A2(n656), .ZN(n516) );
  XOR2_X1 U573 ( .A(KEYINPUT77), .B(n516), .Z(n517) );
  NAND2_X1 U574 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U575 ( .A(n519), .B(KEYINPUT5), .ZN(n526) );
  NOR2_X1 U576 ( .A1(G543), .A2(n520), .ZN(n521) );
  NAND2_X1 U577 ( .A1(G63), .A2(n650), .ZN(n523) );
  NOR2_X2 U578 ( .A1(G651), .A2(n641), .ZN(n651) );
  NAND2_X1 U579 ( .A1(G51), .A2(n651), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U581 ( .A(KEYINPUT6), .B(n524), .Z(n525) );
  NAND2_X1 U582 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U583 ( .A(n527), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U584 ( .A(G2104), .ZN(n536) );
  NOR2_X1 U585 ( .A1(G2105), .A2(n536), .ZN(n551) );
  NAND2_X1 U586 ( .A1(G101), .A2(n551), .ZN(n528) );
  XOR2_X1 U587 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  XNOR2_X1 U588 ( .A(n529), .B(KEYINPUT64), .ZN(n531) );
  AND2_X2 U589 ( .A1(n536), .A2(G2105), .ZN(n881) );
  NAND2_X1 U590 ( .A1(G125), .A2(n881), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U592 ( .A(KEYINPUT65), .B(n532), .ZN(n541) );
  NOR2_X1 U593 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  XNOR2_X2 U594 ( .A(n534), .B(n533), .ZN(n885) );
  XNOR2_X1 U595 ( .A(n535), .B(KEYINPUT66), .ZN(n538) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U597 ( .A1(G113), .A2(n882), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U599 ( .A(n539), .B(KEYINPUT67), .ZN(n540) );
  AND2_X1 U600 ( .A1(n541), .A2(n540), .ZN(G160) );
  XOR2_X1 U601 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U602 ( .A(G2443), .B(G2446), .Z(n543) );
  XNOR2_X1 U603 ( .A(G2427), .B(G2451), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n543), .B(n542), .ZN(n549) );
  XOR2_X1 U605 ( .A(G2430), .B(G2454), .Z(n545) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U608 ( .A(G2435), .B(G2438), .Z(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U610 ( .A(n549), .B(n548), .Z(n550) );
  AND2_X1 U611 ( .A1(G14), .A2(n550), .ZN(G401) );
  NAND2_X1 U612 ( .A1(n882), .A2(G114), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G138), .A2(n885), .ZN(n553) );
  BUF_X1 U614 ( .A(n551), .Z(n886) );
  NAND2_X1 U615 ( .A1(G102), .A2(n886), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G126), .A2(n881), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT88), .B(n554), .Z(n555) );
  NOR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT89), .ZN(G164) );
  NAND2_X1 U622 ( .A1(G64), .A2(n650), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G52), .A2(n651), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G90), .A2(n649), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G77), .A2(n656), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U629 ( .A1(n566), .A2(n565), .ZN(G171) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U631 ( .A(KEYINPUT18), .B(KEYINPUT80), .Z(n568) );
  NAND2_X1 U632 ( .A1(G123), .A2(n881), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G111), .A2(n882), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G135), .A2(n885), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n886), .A2(G99), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n925) );
  XNOR2_X1 U640 ( .A(G2096), .B(n925), .ZN(n575) );
  OR2_X1 U641 ( .A1(G2100), .A2(n575), .ZN(G156) );
  INV_X1 U642 ( .A(G57), .ZN(G237) );
  INV_X1 U643 ( .A(G132), .ZN(G219) );
  NAND2_X1 U644 ( .A1(G88), .A2(n649), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G75), .A2(n656), .ZN(n576) );
  NAND2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G62), .A2(n650), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G50), .A2(n651), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U650 ( .A(KEYINPUT83), .B(n580), .Z(n581) );
  NOR2_X1 U651 ( .A1(n582), .A2(n581), .ZN(G166) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n833) );
  NAND2_X1 U655 ( .A1(n833), .A2(G567), .ZN(n584) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n584), .Z(G234) );
  NAND2_X1 U657 ( .A1(G68), .A2(n656), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT72), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n649), .A2(G81), .ZN(n586) );
  XNOR2_X1 U660 ( .A(KEYINPUT12), .B(n586), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U662 ( .A(n589), .B(KEYINPUT13), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n650), .A2(G56), .ZN(n590) );
  XNOR2_X1 U664 ( .A(KEYINPUT14), .B(n590), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT73), .ZN(n595) );
  NAND2_X1 U667 ( .A1(G43), .A2(n651), .ZN(n594) );
  XNOR2_X2 U668 ( .A(n596), .B(KEYINPUT74), .ZN(n966) );
  NAND2_X1 U669 ( .A1(G860), .A2(n966), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n607) );
  NAND2_X1 U672 ( .A1(G66), .A2(n650), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G92), .A2(n649), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n651), .A2(G54), .ZN(n599) );
  XOR2_X1 U676 ( .A(KEYINPUT75), .B(n599), .Z(n601) );
  NAND2_X1 U677 ( .A1(G79), .A2(n656), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U679 ( .A(KEYINPUT76), .B(n602), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT15), .ZN(n983) );
  INV_X1 U682 ( .A(G868), .ZN(n668) );
  NAND2_X1 U683 ( .A1(n983), .A2(n668), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G65), .A2(n650), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT70), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G91), .A2(n649), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G53), .A2(n651), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G78), .A2(n656), .ZN(n611) );
  XNOR2_X1 U691 ( .A(KEYINPUT69), .B(n611), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G299) );
  XNOR2_X1 U694 ( .A(KEYINPUT78), .B(n668), .ZN(n616) );
  NOR2_X1 U695 ( .A1(G286), .A2(n616), .ZN(n618) );
  NOR2_X1 U696 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G297) );
  INV_X1 U698 ( .A(G860), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n619), .A2(G559), .ZN(n620) );
  INV_X1 U700 ( .A(n983), .ZN(n902) );
  NAND2_X1 U701 ( .A1(n620), .A2(n902), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n621), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U703 ( .A1(G559), .A2(n668), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n902), .A2(n622), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n668), .A2(n966), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U707 ( .A(KEYINPUT79), .B(n625), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G559), .A2(n902), .ZN(n626) );
  XOR2_X1 U709 ( .A(n966), .B(n626), .Z(n665) );
  NOR2_X1 U710 ( .A1(G860), .A2(n665), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G67), .A2(n650), .ZN(n628) );
  NAND2_X1 U712 ( .A1(G55), .A2(n651), .ZN(n627) );
  NAND2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G93), .A2(n649), .ZN(n630) );
  NAND2_X1 U715 ( .A1(G80), .A2(n656), .ZN(n629) );
  NAND2_X1 U716 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n667) );
  XNOR2_X1 U718 ( .A(n633), .B(n667), .ZN(G145) );
  NAND2_X1 U719 ( .A1(G86), .A2(n649), .ZN(n635) );
  NAND2_X1 U720 ( .A1(G48), .A2(n651), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n656), .A2(G73), .ZN(n636) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U725 ( .A1(n650), .A2(G61), .ZN(n639) );
  NAND2_X1 U726 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G87), .A2(n641), .ZN(n642) );
  XNOR2_X1 U728 ( .A(n642), .B(KEYINPUT82), .ZN(n645) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n643) );
  XOR2_X1 U730 ( .A(KEYINPUT81), .B(n643), .Z(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U732 ( .A1(n650), .A2(n646), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n651), .A2(G49), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(G288) );
  AND2_X1 U735 ( .A1(n649), .A2(G85), .ZN(n655) );
  NAND2_X1 U736 ( .A1(G60), .A2(n650), .ZN(n653) );
  NAND2_X1 U737 ( .A1(G47), .A2(n651), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U740 ( .A1(G72), .A2(n656), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n657), .ZN(G290) );
  INV_X1 U742 ( .A(G299), .ZN(n976) );
  XOR2_X1 U743 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n659) );
  XNOR2_X1 U744 ( .A(G288), .B(n659), .ZN(n660) );
  XNOR2_X1 U745 ( .A(n667), .B(n660), .ZN(n662) );
  XNOR2_X1 U746 ( .A(G290), .B(G166), .ZN(n661) );
  XNOR2_X1 U747 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n976), .B(n663), .ZN(n664) );
  XNOR2_X1 U749 ( .A(G305), .B(n664), .ZN(n905) );
  XNOR2_X1 U750 ( .A(n905), .B(n665), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U754 ( .A(KEYINPUT85), .B(n671), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U761 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U762 ( .A1(G219), .A2(G220), .ZN(n676) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  XNOR2_X1 U764 ( .A(n677), .B(KEYINPUT86), .ZN(n678) );
  NOR2_X1 U765 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U766 ( .A1(G96), .A2(n679), .ZN(n839) );
  NAND2_X1 U767 ( .A1(G2106), .A2(n839), .ZN(n680) );
  XOR2_X1 U768 ( .A(KEYINPUT87), .B(n680), .Z(n684) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n681) );
  NOR2_X1 U770 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U771 ( .A1(G108), .A2(n682), .ZN(n838) );
  NAND2_X1 U772 ( .A1(G567), .A2(n838), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n908) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n685) );
  NOR2_X1 U775 ( .A1(n908), .A2(n685), .ZN(n835) );
  NAND2_X1 U776 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NAND2_X2 U779 ( .A1(n687), .A2(n794), .ZN(n736) );
  XNOR2_X1 U780 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n696) );
  INV_X1 U781 ( .A(n696), .ZN(n688) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n688), .ZN(n690) );
  NAND2_X1 U783 ( .A1(G2067), .A2(n983), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n708), .A2(n691), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n692), .A2(n966), .ZN(n701) );
  INV_X1 U787 ( .A(G1341), .ZN(n694) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n983), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n736), .A2(n695), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n708), .A2(G1996), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n706) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n736), .ZN(n703) );
  NAND2_X1 U796 ( .A1(G2067), .A2(n708), .ZN(n702) );
  NAND2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n704), .A2(n983), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n708), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(KEYINPUT27), .ZN(n710) );
  INV_X1 U802 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U803 ( .A1(n998), .A2(n708), .ZN(n709) );
  NOR2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n713), .A2(n976), .ZN(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n713), .A2(n976), .ZN(n715) );
  XNOR2_X1 U808 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NOR2_X1 U811 ( .A1(n736), .A2(n943), .ZN(n721) );
  AND2_X1 U812 ( .A1(n736), .A2(G1961), .ZN(n720) );
  NOR2_X1 U813 ( .A1(n721), .A2(n720), .ZN(n728) );
  NAND2_X1 U814 ( .A1(G171), .A2(n728), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n734) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n774), .ZN(n748) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n736), .ZN(n745) );
  NOR2_X1 U818 ( .A1(n748), .A2(n745), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n724), .A2(G8), .ZN(n726) );
  NOR2_X1 U820 ( .A1(n727), .A2(G168), .ZN(n730) );
  NOR2_X1 U821 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U823 ( .A(n731), .B(KEYINPUT99), .ZN(n732) );
  XNOR2_X1 U824 ( .A(n732), .B(KEYINPUT31), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n746), .A2(G286), .ZN(n735) );
  XNOR2_X1 U827 ( .A(n735), .B(KEYINPUT100), .ZN(n742) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n774), .ZN(n738) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U830 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U831 ( .A(KEYINPUT101), .B(n739), .Z(n740) );
  NAND2_X1 U832 ( .A1(n740), .A2(G303), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U834 ( .A1(n743), .A2(G8), .ZN(n744) );
  XNOR2_X1 U835 ( .A(n744), .B(KEYINPUT32), .ZN(n763) );
  NAND2_X1 U836 ( .A1(G8), .A2(n745), .ZN(n750) );
  INV_X1 U837 ( .A(n746), .ZN(n747) );
  NOR2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n764) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n970) );
  AND2_X1 U841 ( .A1(n764), .A2(n970), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n763), .A2(n751), .ZN(n755) );
  INV_X1 U843 ( .A(n970), .ZN(n753) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n968) );
  NOR2_X1 U846 ( .A1(n971), .A2(n968), .ZN(n752) );
  OR2_X1 U847 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U849 ( .A1(n774), .A2(n756), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n971), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U851 ( .A1(n758), .A2(n774), .ZN(n760) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n987) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n767) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G8), .A2(n765), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n768), .A2(n774), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U860 ( .A(n771), .B(KEYINPUT102), .ZN(n820) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U862 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n818) );
  NAND2_X1 U864 ( .A1(G141), .A2(n885), .ZN(n775) );
  XNOR2_X1 U865 ( .A(n775), .B(KEYINPUT94), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G129), .A2(n881), .ZN(n777) );
  NAND2_X1 U867 ( .A1(G117), .A2(n882), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n886), .A2(G105), .ZN(n778) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n878) );
  NOR2_X1 U873 ( .A1(G1996), .A2(n878), .ZN(n921) );
  NAND2_X1 U874 ( .A1(G119), .A2(n881), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G107), .A2(n882), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U877 ( .A1(G131), .A2(n885), .ZN(n786) );
  NAND2_X1 U878 ( .A1(G95), .A2(n886), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n895) );
  NOR2_X1 U881 ( .A1(G1991), .A2(n895), .ZN(n924) );
  NOR2_X1 U882 ( .A1(G1986), .A2(G290), .ZN(n789) );
  XOR2_X1 U883 ( .A(n789), .B(KEYINPUT103), .Z(n790) );
  NOR2_X1 U884 ( .A1(n924), .A2(n790), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G1991), .A2(n895), .ZN(n792) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n878), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n923) );
  NAND2_X1 U888 ( .A1(G160), .A2(G40), .ZN(n793) );
  NOR2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n824) );
  XOR2_X1 U890 ( .A(n824), .B(KEYINPUT95), .Z(n795) );
  NAND2_X1 U891 ( .A1(n923), .A2(n795), .ZN(n796) );
  XOR2_X1 U892 ( .A(KEYINPUT96), .B(n796), .Z(n821) );
  NOR2_X1 U893 ( .A1(n797), .A2(n821), .ZN(n798) );
  XNOR2_X1 U894 ( .A(n798), .B(KEYINPUT104), .ZN(n799) );
  NOR2_X1 U895 ( .A1(n921), .A2(n799), .ZN(n800) );
  XNOR2_X1 U896 ( .A(n800), .B(KEYINPUT39), .ZN(n814) );
  XNOR2_X1 U897 ( .A(KEYINPUT91), .B(KEYINPUT35), .ZN(n804) );
  NAND2_X1 U898 ( .A1(G128), .A2(n881), .ZN(n802) );
  NAND2_X1 U899 ( .A1(G116), .A2(n882), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U901 ( .A(n804), .B(n803), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n886), .A2(G104), .ZN(n805) );
  XNOR2_X1 U903 ( .A(n805), .B(KEYINPUT90), .ZN(n807) );
  NAND2_X1 U904 ( .A1(G140), .A2(n885), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U906 ( .A(KEYINPUT34), .B(n808), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U908 ( .A(n811), .B(KEYINPUT36), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT92), .ZN(n898) );
  XNOR2_X1 U910 ( .A(KEYINPUT37), .B(G2067), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n898), .A2(n815), .ZN(n932) );
  NAND2_X1 U912 ( .A1(n824), .A2(n932), .ZN(n813) );
  XOR2_X1 U913 ( .A(KEYINPUT93), .B(n813), .Z(n822) );
  NAND2_X1 U914 ( .A1(n814), .A2(n822), .ZN(n816) );
  NAND2_X1 U915 ( .A1(n898), .A2(n815), .ZN(n937) );
  NAND2_X1 U916 ( .A1(n816), .A2(n937), .ZN(n817) );
  AND2_X1 U917 ( .A1(n817), .A2(n824), .ZN(n828) );
  OR2_X1 U918 ( .A1(n818), .A2(n828), .ZN(n819) );
  NOR2_X1 U919 ( .A1(n820), .A2(n819), .ZN(n830) );
  INV_X1 U920 ( .A(n821), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n826) );
  XNOR2_X1 U922 ( .A(G1986), .B(G290), .ZN(n967) );
  AND2_X1 U923 ( .A1(n967), .A2(n824), .ZN(n825) );
  NOR2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U925 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U926 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n831) );
  XNOR2_X1 U927 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U930 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G1), .A2(G3), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n837), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n840), .B(KEYINPUT107), .ZN(G261) );
  INV_X1 U939 ( .A(G261), .ZN(G325) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2084), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2072), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n843), .B(G2100), .Z(n845) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U947 ( .A(KEYINPUT109), .B(G2678), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n849), .B(n848), .Z(G227) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G1976), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U953 ( .A(n852), .B(KEYINPUT111), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1981), .B(G1966), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U956 ( .A(G1971), .B(G1956), .Z(n856) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1961), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U959 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U960 ( .A(G2474), .B(KEYINPUT110), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U962 ( .A1(n881), .A2(G124), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G112), .A2(n882), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n885), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G100), .A2(n886), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U970 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n869) );
  XNOR2_X1 U971 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n880) );
  NAND2_X1 U973 ( .A1(G139), .A2(n885), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G103), .A2(n886), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G127), .A2(n881), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G115), .A2(n882), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n915) );
  XOR2_X1 U981 ( .A(G164), .B(n915), .Z(n877) );
  XNOR2_X1 U982 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U983 ( .A(n880), .B(n879), .ZN(n897) );
  NAND2_X1 U984 ( .A1(G130), .A2(n881), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G118), .A2(n882), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G142), .A2(n885), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G106), .A2(n886), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(n889), .B(KEYINPUT45), .Z(n890) );
  NOR2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n892), .B(n925), .ZN(n893) );
  XOR2_X1 U993 ( .A(G162), .B(n893), .Z(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n900) );
  XOR2_X1 U996 ( .A(n898), .B(G160), .Z(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n966), .B(G286), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(G171), .B(n902), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1002 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G397) );
  XOR2_X1 U1004 ( .A(KEYINPUT108), .B(n908), .Z(G319) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n911), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n912) );
  AND2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n914), .A2(G319), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1015 ( .A(G2072), .B(n915), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G164), .B(G2078), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT116), .ZN(n917) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(KEYINPUT50), .ZN(n935) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n922), .Z(n930) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n928) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(n933), .B(KEYINPUT115), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(n938), .B(KEYINPUT117), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n939), .ZN(n941) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1037 ( .A(G29), .B(KEYINPUT120), .Z(n963) );
  XOR2_X1 U1038 ( .A(G1996), .B(G32), .Z(n945) );
  XNOR2_X1 U1039 ( .A(n943), .B(G27), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(KEYINPUT119), .B(n946), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n954) );
  XOR2_X1 U1046 ( .A(G1991), .B(G25), .Z(n951) );
  NAND2_X1 U1047 ( .A1(n951), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT118), .B(n952), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1050 ( .A(KEYINPUT53), .B(n955), .Z(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT54), .B(G34), .Z(n956) );
  XNOR2_X1 U1052 ( .A(G2084), .B(n956), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n961), .B(KEYINPUT55), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n964), .ZN(n1024) );
  INV_X1 U1059 ( .A(G16), .ZN(n1020) );
  XNOR2_X1 U1060 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n1020), .B(n965), .ZN(n994) );
  XNOR2_X1 U1062 ( .A(G1341), .B(n966), .ZN(n982) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1066 ( .A(n971), .B(KEYINPUT123), .Z(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n976), .B(G1956), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G171), .B(G1961), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(G1348), .B(n983), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT124), .B(n986), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n989), .B(KEYINPUT122), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(KEYINPUT57), .B(n990), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n1022) );
  XNOR2_X1 U1083 ( .A(KEYINPUT127), .B(G1966), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(G21), .ZN(n1015) );
  XNOR2_X1 U1085 ( .A(KEYINPUT60), .B(KEYINPUT126), .ZN(n1006) );
  XNOR2_X1 U1086 ( .A(KEYINPUT125), .B(G1341), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n996), .B(G19), .ZN(n1004) );
  XOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .Z(n997) );
  XNOR2_X1 U1089 ( .A(G4), .B(n997), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(G1981), .B(G6), .Z(n1000) );
  XNOR2_X1 U1091 ( .A(n998), .B(G20), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1006), .B(n1005), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G5), .B(G1961), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

