

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770;

  XOR2_X1 U375 ( .A(n636), .B(n635), .Z(n637) );
  AND2_X1 U376 ( .A1(n389), .A2(n388), .ZN(n387) );
  XOR2_X1 U377 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n556) );
  XNOR2_X1 U378 ( .A(n515), .B(KEYINPUT35), .ZN(n551) );
  NAND2_X1 U379 ( .A1(n514), .A2(n607), .ZN(n515) );
  OR2_X1 U380 ( .A1(n700), .A2(n530), .ZN(n353) );
  INV_X1 U381 ( .A(KEYINPUT31), .ZN(n352) );
  NOR2_X1 U382 ( .A1(n526), .A2(n585), .ZN(n458) );
  AND2_X1 U383 ( .A1(n417), .A2(KEYINPUT1), .ZN(n360) );
  XNOR2_X1 U384 ( .A(n376), .B(n456), .ZN(n652) );
  XNOR2_X1 U385 ( .A(n376), .B(n444), .ZN(n727) );
  XNOR2_X1 U386 ( .A(n380), .B(n378), .ZN(n744) );
  BUF_X1 U387 ( .A(G113), .Z(n354) );
  XNOR2_X1 U388 ( .A(n366), .B(G146), .ZN(n466) );
  INV_X1 U389 ( .A(G125), .ZN(n366) );
  NOR2_X1 U390 ( .A1(n427), .A2(n530), .ZN(n494) );
  BUF_X1 U391 ( .A(n585), .Z(n351) );
  XNOR2_X2 U392 ( .A(n353), .B(n352), .ZN(n678) );
  NAND2_X2 U393 ( .A1(n405), .A2(n404), .ZN(n598) );
  AND2_X2 U394 ( .A1(n365), .A2(n398), .ZN(n368) );
  NAND2_X4 U395 ( .A1(n368), .A2(n369), .ZN(n693) );
  XNOR2_X1 U396 ( .A(G116), .B(G107), .ZN(n459) );
  NOR2_X2 U397 ( .A1(n574), .A2(n694), .ZN(n690) );
  NAND2_X2 U398 ( .A1(n387), .A2(n688), .ZN(n633) );
  XNOR2_X2 U399 ( .A(n557), .B(n556), .ZN(n747) );
  XNOR2_X1 U400 ( .A(n390), .B(KEYINPUT87), .ZN(n377) );
  NOR2_X1 U401 ( .A1(n747), .A2(n385), .ZN(n384) );
  NAND2_X1 U402 ( .A1(n377), .A2(n555), .ZN(n557) );
  NOR2_X1 U403 ( .A1(n713), .A2(n355), .ZN(n426) );
  NOR2_X1 U404 ( .A1(n594), .A2(n593), .ZN(n681) );
  AND2_X1 U405 ( .A1(n421), .A2(n420), .ZN(n419) );
  OR2_X1 U406 ( .A1(n727), .A2(n418), .ZN(n417) );
  XNOR2_X1 U407 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U408 ( .A(n434), .B(G902), .ZN(n475) );
  BUF_X1 U409 ( .A(n427), .Z(n355) );
  XNOR2_X1 U410 ( .A(KEYINPUT4), .B(G131), .ZN(n438) );
  INV_X1 U411 ( .A(n475), .ZN(n629) );
  XNOR2_X1 U412 ( .A(n425), .B(KEYINPUT20), .ZN(n436) );
  NAND2_X1 U413 ( .A1(n475), .A2(G234), .ZN(n425) );
  XNOR2_X1 U414 ( .A(G137), .B(G140), .ZN(n441) );
  INV_X1 U415 ( .A(G146), .ZN(n429) );
  NAND2_X1 U416 ( .A1(n536), .A2(n534), .ZN(n708) );
  NOR2_X1 U417 ( .A1(n484), .A2(KEYINPUT19), .ZN(n410) );
  XNOR2_X1 U418 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n434) );
  NAND2_X1 U419 ( .A1(n399), .A2(G902), .ZN(n398) );
  XNOR2_X1 U420 ( .A(n459), .B(G122), .ZN(n402) );
  XNOR2_X1 U421 ( .A(G101), .B(G107), .ZN(n440) );
  XNOR2_X1 U422 ( .A(n742), .B(KEYINPUT72), .ZN(n464) );
  XNOR2_X1 U423 ( .A(n512), .B(n413), .ZN(n534) );
  XNOR2_X1 U424 ( .A(n511), .B(n513), .ZN(n413) );
  NAND2_X1 U425 ( .A1(n422), .A2(G902), .ZN(n420) );
  NAND2_X1 U426 ( .A1(n445), .A2(n397), .ZN(n418) );
  OR2_X1 U427 ( .A1(n628), .A2(n627), .ZN(n759) );
  INV_X1 U428 ( .A(KEYINPUT23), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n439), .B(G119), .ZN(n460) );
  XNOR2_X1 U430 ( .A(n431), .B(n408), .ZN(n495) );
  INV_X1 U431 ( .A(KEYINPUT8), .ZN(n408) );
  INV_X1 U432 ( .A(G134), .ZN(n437) );
  XNOR2_X1 U433 ( .A(G143), .B(G104), .ZN(n505) );
  XNOR2_X1 U434 ( .A(n354), .B(G131), .ZN(n506) );
  XOR2_X1 U435 ( .A(KEYINPUT11), .B(G122), .Z(n507) );
  XNOR2_X1 U436 ( .A(n504), .B(n358), .ZN(n416) );
  NAND2_X1 U437 ( .A1(n382), .A2(n632), .ZN(n388) );
  INV_X1 U438 ( .A(G214), .ZN(n482) );
  XNOR2_X1 U439 ( .A(n371), .B(n435), .ZN(n370) );
  OR2_X1 U440 ( .A1(n738), .A2(G902), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n502), .B(n501), .ZN(n536) );
  INV_X1 U442 ( .A(KEYINPUT88), .ZN(n394) );
  XNOR2_X1 U443 ( .A(n582), .B(KEYINPUT86), .ZN(n583) );
  AND2_X1 U444 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U445 ( .A1(n681), .A2(n604), .ZN(n613) );
  XNOR2_X1 U446 ( .A(n364), .B(KEYINPUT21), .ZN(n694) );
  XNOR2_X1 U447 ( .A(G137), .B(G116), .ZN(n452) );
  XOR2_X1 U448 ( .A(G119), .B(KEYINPUT5), .Z(n450) );
  NOR2_X1 U449 ( .A1(G953), .A2(G237), .ZN(n503) );
  XNOR2_X1 U450 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n462) );
  XOR2_X1 U451 ( .A(KEYINPUT94), .B(KEYINPUT18), .Z(n463) );
  XNOR2_X1 U452 ( .A(KEYINPUT4), .B(KEYINPUT80), .ZN(n469) );
  NAND2_X1 U453 ( .A1(n383), .A2(n359), .ZN(n382) );
  INV_X1 U454 ( .A(n627), .ZN(n428) );
  NAND2_X1 U455 ( .A1(G234), .A2(G237), .ZN(n485) );
  NOR2_X1 U456 ( .A1(G237), .A2(G902), .ZN(n476) );
  NAND2_X1 U457 ( .A1(n436), .A2(G217), .ZN(n371) );
  NAND2_X1 U458 ( .A1(n457), .A2(n397), .ZN(n396) );
  NOR2_X1 U459 ( .A1(n708), .A2(n694), .ZN(n516) );
  XNOR2_X1 U460 ( .A(n461), .B(n402), .ZN(n380) );
  INV_X1 U461 ( .A(KEYINPUT16), .ZN(n379) );
  XNOR2_X1 U462 ( .A(n423), .B(n464), .ZN(n444) );
  XNOR2_X1 U463 ( .A(n442), .B(n424), .ZN(n423) );
  XNOR2_X1 U464 ( .A(n443), .B(n439), .ZN(n424) );
  INV_X1 U465 ( .A(n759), .ZN(n386) );
  INV_X1 U466 ( .A(KEYINPUT2), .ZN(n385) );
  AND2_X1 U467 ( .A1(n403), .A2(n412), .ZN(n405) );
  NAND2_X1 U468 ( .A1(n624), .A2(KEYINPUT19), .ZN(n404) );
  NAND2_X1 U469 ( .A1(n484), .A2(KEYINPUT19), .ZN(n412) );
  INV_X1 U470 ( .A(n534), .ZN(n535) );
  XNOR2_X1 U471 ( .A(n652), .B(n654), .ZN(n655) );
  XNOR2_X1 U472 ( .A(n409), .B(n407), .ZN(n433) );
  NAND2_X1 U473 ( .A1(n495), .A2(G221), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n498), .B(n381), .ZN(n733) );
  XNOR2_X1 U475 ( .A(n510), .B(n414), .ZN(n643) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n505), .B(G140), .ZN(n415) );
  AND2_X1 U478 ( .A1(n639), .A2(G953), .ZN(n741) );
  NOR2_X1 U479 ( .A1(n536), .A2(n535), .ZN(n668) );
  NAND2_X1 U480 ( .A1(n536), .A2(n535), .ZN(n676) );
  INV_X1 U481 ( .A(G143), .ZN(n650) );
  XOR2_X1 U482 ( .A(n480), .B(n479), .Z(n356) );
  AND2_X1 U483 ( .A1(n417), .A2(n419), .ZN(n357) );
  AND2_X1 U484 ( .A1(G214), .A2(n503), .ZN(n358) );
  INV_X1 U485 ( .A(G902), .ZN(n397) );
  INV_X1 U486 ( .A(G110), .ZN(n439) );
  AND2_X1 U487 ( .A1(n428), .A2(n629), .ZN(n359) );
  INV_X1 U488 ( .A(KEYINPUT1), .ZN(n400) );
  NAND2_X1 U489 ( .A1(n360), .A2(n419), .ZN(n401) );
  NAND2_X1 U490 ( .A1(n363), .A2(n400), .ZN(n362) );
  NAND2_X1 U491 ( .A1(n361), .A2(n690), .ZN(n526) );
  NAND2_X1 U492 ( .A1(n362), .A2(n401), .ZN(n361) );
  NAND2_X1 U493 ( .A1(n419), .A2(n417), .ZN(n363) );
  NAND2_X1 U494 ( .A1(n436), .A2(G221), .ZN(n364) );
  NAND2_X1 U495 ( .A1(n652), .A2(n399), .ZN(n365) );
  XNOR2_X2 U496 ( .A(n758), .B(n429), .ZN(n376) );
  NAND2_X1 U497 ( .A1(n598), .A2(n492), .ZN(n493) );
  NAND2_X1 U498 ( .A1(n362), .A2(n401), .ZN(n367) );
  XNOR2_X1 U499 ( .A(n375), .B(n460), .ZN(n409) );
  XNOR2_X1 U500 ( .A(n374), .B(G128), .ZN(n373) );
  AND2_X1 U501 ( .A1(n525), .A2(n524), .ZN(n540) );
  NAND2_X1 U502 ( .A1(n540), .A2(n539), .ZN(n395) );
  NOR2_X1 U503 ( .A1(n526), .A2(n532), .ZN(n528) );
  OR2_X1 U504 ( .A1(n652), .A2(n396), .ZN(n369) );
  BUF_X1 U505 ( .A(n726), .Z(n737) );
  XNOR2_X2 U506 ( .A(n372), .B(n370), .ZN(n574) );
  XNOR2_X1 U507 ( .A(n433), .B(n757), .ZN(n738) );
  XNOR2_X1 U508 ( .A(n432), .B(n373), .ZN(n375) );
  NAND2_X1 U509 ( .A1(n384), .A2(n386), .ZN(n688) );
  XNOR2_X1 U510 ( .A(n460), .B(n379), .ZN(n378) );
  INV_X2 U511 ( .A(n446), .ZN(n448) );
  INV_X2 U512 ( .A(G128), .ZN(n406) );
  NAND2_X1 U513 ( .A1(n393), .A2(n391), .ZN(n390) );
  XNOR2_X1 U514 ( .A(n500), .B(n499), .ZN(n381) );
  INV_X1 U515 ( .A(n628), .ZN(n383) );
  NOR2_X1 U516 ( .A1(n759), .A2(n748), .ZN(n684) );
  NAND2_X1 U517 ( .A1(n747), .A2(n632), .ZN(n389) );
  XNOR2_X1 U518 ( .A(n550), .B(KEYINPUT89), .ZN(n553) );
  INV_X1 U519 ( .A(n553), .ZN(n392) );
  NAND2_X1 U520 ( .A1(n392), .A2(KEYINPUT44), .ZN(n391) );
  XNOR2_X1 U521 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X2 U522 ( .A(n693), .B(KEYINPUT6), .ZN(n585) );
  INV_X1 U523 ( .A(n457), .ZN(n399) );
  XNOR2_X1 U524 ( .A(n402), .B(KEYINPUT7), .ZN(n496) );
  NAND2_X1 U525 ( .A1(n411), .A2(n410), .ZN(n403) );
  XNOR2_X2 U526 ( .A(n481), .B(n356), .ZN(n411) );
  INV_X2 U527 ( .A(n411), .ZN(n624) );
  XNOR2_X2 U528 ( .A(n406), .B(G143), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n411), .A2(n706), .ZN(n590) );
  XNOR2_X2 U530 ( .A(KEYINPUT3), .B(KEYINPUT71), .ZN(n447) );
  XNOR2_X2 U531 ( .A(n448), .B(n447), .ZN(n461) );
  NAND2_X1 U532 ( .A1(n727), .A2(n422), .ZN(n421) );
  INV_X1 U533 ( .A(n445), .ZN(n422) );
  NOR2_X1 U534 ( .A1(n355), .A2(n719), .ZN(n720) );
  XNOR2_X1 U535 ( .A(n458), .B(KEYINPUT33), .ZN(n427) );
  XNOR2_X2 U536 ( .A(n500), .B(n438), .ZN(n758) );
  XNOR2_X2 U537 ( .A(n467), .B(n437), .ZN(n500) );
  NOR2_X2 U538 ( .A1(n530), .A2(n517), .ZN(n519) );
  XNOR2_X2 U539 ( .A(n493), .B(KEYINPUT0), .ZN(n530) );
  INV_X1 U540 ( .A(KEYINPUT83), .ZN(n596) );
  XNOR2_X1 U541 ( .A(n597), .B(n596), .ZN(n603) );
  INV_X1 U542 ( .A(KEYINPUT101), .ZN(n451) );
  XNOR2_X1 U543 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U544 ( .A(KEYINPUT46), .ZN(n582) );
  XNOR2_X1 U545 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U546 ( .A(n584), .B(n583), .ZN(n616) );
  XNOR2_X1 U547 ( .A(KEYINPUT48), .B(KEYINPUT85), .ZN(n617) );
  INV_X1 U548 ( .A(KEYINPUT102), .ZN(n527) );
  BUF_X1 U549 ( .A(n634), .Z(n635) );
  XNOR2_X1 U550 ( .A(n466), .B(KEYINPUT10), .ZN(n509) );
  INV_X1 U551 ( .A(n509), .ZN(n430) );
  XNOR2_X1 U552 ( .A(n430), .B(n441), .ZN(n757) );
  XOR2_X1 U553 ( .A(KEYINPUT24), .B(KEYINPUT99), .Z(n432) );
  INV_X2 U554 ( .A(G953), .ZN(n760) );
  NAND2_X1 U555 ( .A1(G234), .A2(n760), .ZN(n431) );
  XOR2_X1 U556 ( .A(KEYINPUT79), .B(KEYINPUT25), .Z(n435) );
  XNOR2_X2 U557 ( .A(KEYINPUT93), .B(G104), .ZN(n742) );
  XNOR2_X1 U558 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U559 ( .A1(G227), .A2(n760), .ZN(n443) );
  XNOR2_X1 U560 ( .A(KEYINPUT70), .B(G469), .ZN(n445) );
  XNOR2_X1 U561 ( .A(G472), .B(KEYINPUT75), .ZN(n457) );
  XNOR2_X2 U562 ( .A(G101), .B(G113), .ZN(n446) );
  NAND2_X1 U563 ( .A1(n503), .A2(G210), .ZN(n449) );
  XNOR2_X1 U564 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U565 ( .A(n461), .B(n455), .ZN(n456) );
  XNOR2_X1 U566 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U567 ( .A(n465), .B(n464), .ZN(n473) );
  XNOR2_X1 U568 ( .A(n467), .B(n466), .ZN(n471) );
  AND2_X1 U569 ( .A1(n760), .A2(G224), .ZN(n468) );
  XNOR2_X1 U570 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U571 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U572 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n744), .B(n474), .ZN(n634) );
  NAND2_X1 U574 ( .A1(n634), .A2(n475), .ZN(n481) );
  XNOR2_X1 U575 ( .A(n476), .B(KEYINPUT78), .ZN(n483) );
  INV_X1 U576 ( .A(G210), .ZN(n477) );
  OR2_X1 U577 ( .A1(n483), .A2(n477), .ZN(n480) );
  INV_X1 U578 ( .A(KEYINPUT95), .ZN(n478) );
  XNOR2_X1 U579 ( .A(n478), .B(KEYINPUT96), .ZN(n479) );
  OR2_X1 U580 ( .A1(n483), .A2(n482), .ZN(n706) );
  INV_X1 U581 ( .A(n706), .ZN(n484) );
  XOR2_X1 U582 ( .A(KEYINPUT97), .B(KEYINPUT14), .Z(n486) );
  XNOR2_X1 U583 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U584 ( .A(KEYINPUT76), .B(n487), .ZN(n489) );
  NAND2_X1 U585 ( .A1(G952), .A2(n489), .ZN(n718) );
  NOR2_X1 U586 ( .A1(n718), .A2(G953), .ZN(n488) );
  XNOR2_X1 U587 ( .A(n488), .B(KEYINPUT98), .ZN(n564) );
  AND2_X1 U588 ( .A1(n489), .A2(G953), .ZN(n490) );
  NAND2_X1 U589 ( .A1(G902), .A2(n490), .ZN(n561) );
  NOR2_X1 U590 ( .A1(n561), .A2(G898), .ZN(n491) );
  OR2_X1 U591 ( .A1(n564), .A2(n491), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n494), .B(KEYINPUT34), .ZN(n514) );
  NAND2_X1 U593 ( .A1(n495), .A2(G217), .ZN(n499) );
  XOR2_X1 U594 ( .A(KEYINPUT105), .B(KEYINPUT9), .Z(n497) );
  XNOR2_X1 U595 ( .A(n497), .B(n496), .ZN(n498) );
  NOR2_X1 U596 ( .A1(G902), .A2(n733), .ZN(n502) );
  XNOR2_X1 U597 ( .A(KEYINPUT106), .B(G478), .ZN(n501) );
  INV_X1 U598 ( .A(G475), .ZN(n513) );
  XOR2_X1 U599 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n504) );
  XNOR2_X1 U600 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U601 ( .A(n509), .B(n508), .ZN(n510) );
  NOR2_X1 U602 ( .A1(G902), .A2(n643), .ZN(n512) );
  XNOR2_X1 U603 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n511) );
  NOR2_X1 U604 ( .A1(n536), .A2(n534), .ZN(n607) );
  NAND2_X1 U605 ( .A1(n551), .A2(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U606 ( .A(n516), .B(KEYINPUT109), .ZN(n517) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(KEYINPUT22), .Z(n518) );
  XNOR2_X2 U608 ( .A(n519), .B(n518), .ZN(n549) );
  INV_X1 U609 ( .A(n549), .ZN(n523) );
  INV_X1 U610 ( .A(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U611 ( .A(n574), .B(n520), .ZN(n696) );
  INV_X1 U612 ( .A(n696), .ZN(n541) );
  NOR2_X1 U613 ( .A1(n367), .A2(n541), .ZN(n521) );
  NAND2_X1 U614 ( .A1(n521), .A2(n351), .ZN(n522) );
  NOR2_X1 U615 ( .A1(n523), .A2(n522), .ZN(n660) );
  INV_X1 U616 ( .A(n660), .ZN(n524) );
  INV_X1 U617 ( .A(n693), .ZN(n532) );
  XNOR2_X1 U618 ( .A(n528), .B(n527), .ZN(n700) );
  NAND2_X1 U619 ( .A1(n690), .A2(n357), .ZN(n565) );
  NOR2_X1 U620 ( .A1(n530), .A2(n565), .ZN(n531) );
  XNOR2_X1 U621 ( .A(n531), .B(KEYINPUT100), .ZN(n533) );
  NAND2_X1 U622 ( .A1(n533), .A2(n532), .ZN(n664) );
  NAND2_X1 U623 ( .A1(n678), .A2(n664), .ZN(n537) );
  XNOR2_X1 U624 ( .A(KEYINPUT107), .B(n668), .ZN(n619) );
  NAND2_X1 U625 ( .A1(n676), .A2(n619), .ZN(n595) );
  NAND2_X1 U626 ( .A1(n537), .A2(n595), .ZN(n538) );
  XNOR2_X1 U627 ( .A(n538), .B(KEYINPUT108), .ZN(n539) );
  XNOR2_X1 U628 ( .A(n351), .B(KEYINPUT81), .ZN(n543) );
  NAND2_X1 U629 ( .A1(n367), .A2(n541), .ZN(n542) );
  NOR2_X1 U630 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U631 ( .A1(n549), .A2(n544), .ZN(n546) );
  XNOR2_X1 U632 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n545) );
  XNOR2_X2 U633 ( .A(n546), .B(n545), .ZN(n648) );
  INV_X1 U634 ( .A(n367), .ZN(n593) );
  NAND2_X1 U635 ( .A1(n593), .A2(n574), .ZN(n547) );
  XNOR2_X1 U636 ( .A(n693), .B(KEYINPUT111), .ZN(n575) );
  INV_X1 U637 ( .A(n575), .ZN(n558) );
  NOR2_X1 U638 ( .A1(n547), .A2(n558), .ZN(n548) );
  NAND2_X1 U639 ( .A1(n549), .A2(n548), .ZN(n667) );
  NAND2_X1 U640 ( .A1(n648), .A2(n667), .ZN(n550) );
  BUF_X1 U641 ( .A(n551), .Z(n768) );
  NOR2_X1 U642 ( .A1(n768), .A2(KEYINPUT44), .ZN(n552) );
  AND2_X1 U643 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U644 ( .A(n554), .B(KEYINPUT73), .ZN(n555) );
  INV_X1 U645 ( .A(KEYINPUT30), .ZN(n560) );
  NAND2_X1 U646 ( .A1(n558), .A2(n706), .ZN(n559) );
  XNOR2_X1 U647 ( .A(n560), .B(n559), .ZN(n606) );
  NOR2_X1 U648 ( .A1(G900), .A2(n561), .ZN(n562) );
  XNOR2_X1 U649 ( .A(n562), .B(KEYINPUT112), .ZN(n563) );
  NOR2_X1 U650 ( .A1(n564), .A2(n563), .ZN(n572) );
  NOR2_X1 U651 ( .A1(n565), .A2(n572), .ZN(n605) );
  XOR2_X1 U652 ( .A(KEYINPUT77), .B(KEYINPUT38), .Z(n566) );
  XNOR2_X1 U653 ( .A(n624), .B(n566), .ZN(n705) );
  AND2_X1 U654 ( .A1(n605), .A2(n705), .ZN(n567) );
  NAND2_X1 U655 ( .A1(n606), .A2(n567), .ZN(n569) );
  XOR2_X1 U656 ( .A(KEYINPUT74), .B(KEYINPUT39), .Z(n568) );
  XNOR2_X1 U657 ( .A(n569), .B(n568), .ZN(n620) );
  NOR2_X1 U658 ( .A1(n620), .A2(n676), .ZN(n571) );
  XNOR2_X1 U659 ( .A(KEYINPUT114), .B(KEYINPUT40), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n571), .B(n570), .ZN(n769) );
  NOR2_X1 U661 ( .A1(n572), .A2(n694), .ZN(n573) );
  NAND2_X1 U662 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U663 ( .A1(n575), .A2(n586), .ZN(n576) );
  XNOR2_X1 U664 ( .A(KEYINPUT28), .B(n576), .ZN(n577) );
  NAND2_X1 U665 ( .A1(n357), .A2(n577), .ZN(n600) );
  INV_X1 U666 ( .A(n600), .ZN(n580) );
  NAND2_X1 U667 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U668 ( .A1(n709), .A2(n708), .ZN(n578) );
  XNOR2_X1 U669 ( .A(KEYINPUT41), .B(n578), .ZN(n719) );
  INV_X1 U670 ( .A(n719), .ZN(n579) );
  NAND2_X1 U671 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U672 ( .A(KEYINPUT42), .B(n581), .Z(n770) );
  NOR2_X1 U673 ( .A1(n769), .A2(n770), .ZN(n584) );
  NOR2_X1 U674 ( .A1(n676), .A2(n585), .ZN(n588) );
  INV_X1 U675 ( .A(n586), .ZN(n587) );
  NAND2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U677 ( .A(KEYINPUT113), .B(n589), .Z(n621) );
  NOR2_X1 U678 ( .A1(n621), .A2(n590), .ZN(n592) );
  XNOR2_X1 U679 ( .A(KEYINPUT115), .B(KEYINPUT36), .ZN(n591) );
  XNOR2_X1 U680 ( .A(n592), .B(n591), .ZN(n594) );
  INV_X1 U681 ( .A(n595), .ZN(n710) );
  NAND2_X1 U682 ( .A1(n710), .A2(KEYINPUT47), .ZN(n597) );
  INV_X1 U683 ( .A(n598), .ZN(n599) );
  NOR2_X1 U684 ( .A1(n600), .A2(n599), .ZN(n673) );
  INV_X1 U685 ( .A(n673), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n601), .A2(KEYINPUT47), .ZN(n602) );
  NAND2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U690 ( .A1(n609), .A2(n624), .ZN(n651) );
  NOR2_X1 U691 ( .A1(KEYINPUT47), .A2(n710), .ZN(n610) );
  AND2_X1 U692 ( .A1(n673), .A2(n610), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n651), .A2(n611), .ZN(n612) );
  XNOR2_X1 U694 ( .A(KEYINPUT69), .B(n614), .ZN(n615) );
  NOR2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(n617), .ZN(n628) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n683) );
  INV_X1 U698 ( .A(n683), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n367), .A2(n621), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n622), .A2(n706), .ZN(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT43), .B(n623), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n649) );
  NAND2_X1 U703 ( .A1(n626), .A2(n649), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n629), .B(KEYINPUT84), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n630), .A2(KEYINPUT2), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT68), .ZN(n632) );
  XNOR2_X2 U707 ( .A(n633), .B(KEYINPUT65), .ZN(n726) );
  NAND2_X1 U708 ( .A1(n726), .A2(G210), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n636) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n640) );
  INV_X1 U711 ( .A(G952), .ZN(n639) );
  NOR2_X2 U712 ( .A1(n640), .A2(n741), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U714 ( .A1(n726), .A2(G475), .ZN(n645) );
  INV_X1 U715 ( .A(KEYINPUT59), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X2 U717 ( .A1(n646), .A2(n741), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U719 ( .A(n648), .B(G119), .ZN(G21) );
  XNOR2_X1 U720 ( .A(n649), .B(G140), .ZN(G42) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(G45) );
  NAND2_X1 U722 ( .A1(n726), .A2(G472), .ZN(n656) );
  XNOR2_X1 U723 ( .A(KEYINPUT91), .B(KEYINPUT116), .ZN(n653) );
  XOR2_X1 U724 ( .A(n653), .B(KEYINPUT62), .Z(n654) );
  XNOR2_X1 U725 ( .A(n656), .B(n655), .ZN(n657) );
  NOR2_X2 U726 ( .A1(n657), .A2(n741), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT117), .B(KEYINPUT63), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(G57) );
  XOR2_X1 U729 ( .A(G101), .B(n660), .Z(G3) );
  NOR2_X1 U730 ( .A1(n676), .A2(n664), .ZN(n661) );
  XOR2_X1 U731 ( .A(G104), .B(n661), .Z(G6) );
  XOR2_X1 U732 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n663) );
  XNOR2_X1 U733 ( .A(G107), .B(KEYINPUT118), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n666) );
  INV_X1 U735 ( .A(n668), .ZN(n679) );
  NOR2_X1 U736 ( .A1(n679), .A2(n664), .ZN(n665) );
  XOR2_X1 U737 ( .A(n666), .B(n665), .Z(G9) );
  XNOR2_X1 U738 ( .A(G110), .B(n667), .ZN(G12) );
  XOR2_X1 U739 ( .A(KEYINPUT119), .B(KEYINPUT29), .Z(n670) );
  NAND2_X1 U740 ( .A1(n673), .A2(n668), .ZN(n669) );
  XNOR2_X1 U741 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U742 ( .A(G128), .B(n671), .Z(G30) );
  INV_X1 U743 ( .A(n676), .ZN(n672) );
  AND2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U745 ( .A(KEYINPUT120), .B(n674), .Z(n675) );
  XNOR2_X1 U746 ( .A(G146), .B(n675), .ZN(G48) );
  NOR2_X1 U747 ( .A1(n676), .A2(n678), .ZN(n677) );
  XOR2_X1 U748 ( .A(n354), .B(n677), .Z(G15) );
  NOR2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U750 ( .A(G116), .B(n680), .Z(G18) );
  XNOR2_X1 U751 ( .A(G125), .B(n681), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n682), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U753 ( .A(G134), .B(n683), .Z(G36) );
  OR2_X1 U754 ( .A1(n684), .A2(KEYINPUT2), .ZN(n685) );
  NAND2_X1 U755 ( .A1(n685), .A2(KEYINPUT82), .ZN(n687) );
  OR2_X1 U756 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n686) );
  NAND2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n723) );
  NOR2_X1 U759 ( .A1(n690), .A2(n367), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT50), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n699) );
  INV_X1 U762 ( .A(n694), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT49), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U767 ( .A(n702), .B(KEYINPUT121), .ZN(n703) );
  XOR2_X1 U768 ( .A(KEYINPUT51), .B(n703), .Z(n704) );
  NOR2_X1 U769 ( .A1(n719), .A2(n704), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n714), .A2(n426), .ZN(n715) );
  XNOR2_X1 U775 ( .A(n715), .B(KEYINPUT122), .ZN(n716) );
  XNOR2_X1 U776 ( .A(KEYINPUT52), .B(n716), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n721) );
  NOR2_X1 U778 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U780 ( .A1(n724), .A2(G953), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n725), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U782 ( .A1(n737), .A2(G469), .ZN(n731) );
  XNOR2_X1 U783 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n729) );
  XNOR2_X1 U784 ( .A(n727), .B(KEYINPUT57), .ZN(n728) );
  XNOR2_X1 U785 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U786 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n741), .A2(n732), .ZN(G54) );
  NAND2_X1 U788 ( .A1(n737), .A2(G478), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n733), .B(KEYINPUT124), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U791 ( .A1(n741), .A2(n736), .ZN(G63) );
  NAND2_X1 U792 ( .A1(n737), .A2(G217), .ZN(n739) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U794 ( .A1(n741), .A2(n740), .ZN(G66) );
  XOR2_X1 U795 ( .A(KEYINPUT126), .B(n742), .Z(n743) );
  XNOR2_X1 U796 ( .A(n744), .B(n743), .ZN(n746) );
  NOR2_X1 U797 ( .A1(G898), .A2(n760), .ZN(n745) );
  NOR2_X1 U798 ( .A1(n746), .A2(n745), .ZN(n756) );
  BUF_X1 U799 ( .A(n747), .Z(n748) );
  NOR2_X1 U800 ( .A1(n748), .A2(G953), .ZN(n754) );
  INV_X1 U801 ( .A(G898), .ZN(n752) );
  NAND2_X1 U802 ( .A1(G224), .A2(G953), .ZN(n749) );
  XNOR2_X1 U803 ( .A(n749), .B(KEYINPUT125), .ZN(n750) );
  XNOR2_X1 U804 ( .A(n750), .B(KEYINPUT61), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U807 ( .A(n756), .B(n755), .Z(G69) );
  XOR2_X1 U808 ( .A(n758), .B(n757), .Z(n762) );
  XNOR2_X1 U809 ( .A(n759), .B(n762), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(n760), .ZN(n767) );
  XNOR2_X1 U811 ( .A(G227), .B(n762), .ZN(n763) );
  NAND2_X1 U812 ( .A1(n763), .A2(G900), .ZN(n764) );
  XOR2_X1 U813 ( .A(KEYINPUT127), .B(n764), .Z(n765) );
  NAND2_X1 U814 ( .A1(G953), .A2(n765), .ZN(n766) );
  NAND2_X1 U815 ( .A1(n767), .A2(n766), .ZN(G72) );
  XOR2_X1 U816 ( .A(G122), .B(n768), .Z(G24) );
  XOR2_X1 U817 ( .A(G131), .B(n769), .Z(G33) );
  XOR2_X1 U818 ( .A(G137), .B(n770), .Z(G39) );
endmodule

