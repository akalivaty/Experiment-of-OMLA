//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n467), .B(G125), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G101), .A3(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(new_n465), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(G137), .A3(new_n474), .ZN(new_n477));
  AND3_X1   g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(new_n470), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n483), .B2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n474), .B1(new_n464), .B2(new_n465), .ZN(new_n485));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n485), .B2(G124), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n485), .A2(KEYINPUT69), .A3(G124), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G138), .B(new_n474), .C1(new_n469), .C2(new_n470), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n476), .A2(new_n492), .A3(G138), .A4(new_n474), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n474), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n498), .A2(new_n502), .B1(new_n485), .B2(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(new_n506), .B2(new_n507), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(new_n510), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n514), .A2(new_n513), .ZN(new_n527));
  OAI21_X1  g102(.A(G89), .B1(new_n506), .B2(new_n507), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n510), .A2(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n515), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n519), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(new_n517), .A2(G56), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n519), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(KEYINPUT71), .ZN(new_n542));
  INV_X1    g117(.A(new_n515), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT72), .B(G43), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n543), .A2(G81), .B1(new_n510), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n541), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n541), .A2(KEYINPUT73), .A3(new_n542), .A4(new_n545), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT74), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT76), .B(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n527), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(G651), .A2(new_n559), .B1(new_n543), .B2(G91), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n524), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n510), .A2(new_n564), .A3(G53), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n563), .B1(new_n562), .B2(new_n565), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n560), .B1(new_n567), .B2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  OR2_X1    g145(.A1(new_n526), .A2(new_n530), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT77), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND2_X1  g148(.A1(new_n543), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n510), .A2(G49), .ZN(new_n575));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n527), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT78), .B1(new_n577), .B2(G651), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  AOI211_X1 g154(.A(new_n579), .B(new_n519), .C1(new_n527), .C2(new_n576), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n574), .B(new_n575), .C1(new_n578), .C2(new_n580), .ZN(G288));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n519), .ZN(new_n584));
  OAI211_X1 g159(.A(G48), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n515), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n527), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(KEYINPUT79), .A3(G651), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n584), .A2(new_n588), .A3(new_n592), .ZN(G305));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n527), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(G72), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(G85), .A2(new_n543), .B1(new_n510), .B2(G47), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n597), .A2(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n543), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n527), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n510), .B2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n604), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n604), .B1(new_n612), .B2(G868), .ZN(G321));
  MUX2_X1   g189(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g190(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g191(.A(KEYINPUT81), .B(G559), .Z(new_n617));
  OAI21_X1  g192(.A(new_n612), .B1(G860), .B2(new_n617), .ZN(G148));
  NAND2_X1  g193(.A1(new_n612), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n483), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n485), .A2(G123), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n628), .A2(new_n634), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT83), .B(KEYINPUT14), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT17), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2084), .B(G2090), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n656), .B1(new_n653), .B2(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n655), .ZN(new_n659));
  INV_X1    g234(.A(new_n655), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n660), .A2(new_n656), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n657), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n674), .B1(KEYINPUT85), .B2(new_n675), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(KEYINPUT85), .B2(new_n675), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n678), .A2(KEYINPUT20), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(KEYINPUT20), .ZN(new_n680));
  OAI221_X1 g255(.A(new_n676), .B1(new_n674), .B2(new_n672), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n668), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(new_n667), .A3(new_n687), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(G229));
  INV_X1    g268(.A(G288), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(G23), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n695), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1971), .Z(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n700), .A2(new_n701), .A3(new_n704), .A4(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT34), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G24), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n601), .A2(new_n602), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G1986), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(G1986), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT88), .B(G29), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n483), .A2(G131), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g296(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n722));
  OAI221_X1 g297(.A(G2104), .B1(G107), .B2(new_n474), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n485), .A2(G119), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n718), .B1(new_n726), .B2(new_n717), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  XOR2_X1   g303(.A(new_n727), .B(new_n728), .Z(new_n729));
  NOR2_X1   g304(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n709), .A2(new_n710), .A3(new_n714), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT36), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n695), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n695), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n627), .A2(new_n716), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT30), .B(G28), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n474), .A2(G105), .A3(G2104), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n483), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n485), .A2(G129), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT26), .Z(new_n748));
  AND4_X1   g323(.A1(new_n744), .A2(new_n745), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(new_n741), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n741), .B2(G32), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n736), .B(new_n743), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n716), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n483), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n485), .A2(G128), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n741), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT91), .B(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n741), .A2(G33), .ZN(new_n766));
  AND2_X1   g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n476), .B2(G127), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n768), .A2(KEYINPUT92), .A3(new_n474), .ZN(new_n769));
  OAI21_X1  g344(.A(KEYINPUT92), .B1(new_n768), .B2(new_n474), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT25), .ZN(new_n771));
  NAND2_X1  g346(.A1(G103), .A2(G2104), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n474), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n483), .A2(G139), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n769), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n766), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n754), .A2(new_n765), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n717), .A2(G27), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n717), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT97), .B(G2078), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n753), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G34), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n716), .B1(new_n786), .B2(G34), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT93), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G160), .B2(G29), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT94), .Z(new_n793));
  INV_X1    g368(.A(G2084), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n777), .A2(new_n778), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n695), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  INV_X1    g374(.A(new_n560), .ZN(new_n800));
  INV_X1    g375(.A(new_n568), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n566), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n799), .B1(new_n802), .B2(new_n695), .ZN(new_n803));
  INV_X1    g378(.A(G1956), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n785), .A2(new_n795), .A3(new_n797), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n793), .A2(new_n794), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT96), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n695), .A2(G19), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n550), .B2(new_n695), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT90), .B(G1341), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n717), .A2(G35), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n717), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(G2090), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n695), .A2(G5), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G171), .B2(new_n695), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1961), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n695), .A2(G4), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n612), .B2(new_n695), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n819), .B1(new_n821), .B2(G1348), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(G1348), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n815), .A2(G2090), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n816), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n806), .A2(new_n808), .A3(new_n812), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n732), .A2(new_n826), .ZN(G150));
  INV_X1    g402(.A(G150), .ZN(G311));
  NAND2_X1  g403(.A1(new_n517), .A2(G67), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n519), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n833));
  AOI22_X1  g408(.A1(G93), .A2(new_n543), .B1(new_n510), .B2(G55), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n612), .A2(G559), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n548), .A2(new_n549), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n835), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n835), .A2(new_n546), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  INV_X1    g421(.A(G860), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n837), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT100), .ZN(G145));
  XNOR2_X1  g425(.A(new_n776), .B(new_n749), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n485), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n474), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G142), .B2(new_n483), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n630), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n851), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n504), .B(new_n761), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n726), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G160), .B(new_n488), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(new_n627), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n860), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n863), .B1(new_n861), .B2(new_n864), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n867), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g451(.A1(G290), .A2(G288), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(G290), .A2(G288), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n712), .A2(new_n694), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(KEYINPUT104), .A3(new_n877), .ZN(new_n882));
  XOR2_X1   g457(.A(G166), .B(G305), .Z(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n883), .A2(new_n881), .A3(KEYINPUT104), .A4(new_n877), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  MUX2_X1   g466(.A(new_n887), .B(new_n891), .S(KEYINPUT42), .Z(new_n892));
  NAND2_X1  g467(.A1(new_n612), .A2(new_n802), .ZN(new_n893));
  NAND2_X1  g468(.A1(G299), .A2(new_n611), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n893), .A2(new_n894), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT103), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n844), .B(new_n619), .ZN(new_n902));
  MUX2_X1   g477(.A(new_n899), .B(new_n901), .S(new_n902), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n892), .B(new_n903), .ZN(new_n904));
  MUX2_X1   g479(.A(new_n835), .B(new_n904), .S(G868), .Z(G295));
  MUX2_X1   g480(.A(new_n835), .B(new_n904), .S(G868), .Z(G331));
  NOR2_X1   g481(.A1(G171), .A2(G168), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(G286), .B2(G301), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n842), .A3(new_n843), .ZN(new_n910));
  XNOR2_X1  g485(.A(G168), .B(KEYINPUT77), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n907), .B1(new_n911), .B2(G171), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n844), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n910), .A2(new_n913), .A3(new_n897), .A4(new_n898), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n844), .A2(new_n912), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n844), .A2(new_n912), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n900), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n885), .A2(new_n889), .A3(new_n886), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n889), .B1(new_n885), .B2(new_n886), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n914), .B(new_n917), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n891), .A2(KEYINPUT106), .A3(new_n914), .A4(new_n917), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n918), .A2(new_n919), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n917), .A2(new_n914), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n915), .A2(new_n916), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n914), .B1(new_n901), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n925), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(KEYINPUT43), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n920), .B2(new_n921), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT43), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n927), .A4(new_n923), .ZN(new_n940));
  AND4_X1   g515(.A1(KEYINPUT107), .A2(new_n937), .A3(KEYINPUT44), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n935), .B1(new_n933), .B2(KEYINPUT43), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT107), .B1(new_n942), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n936), .B1(new_n941), .B2(new_n943), .ZN(G397));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT45), .B1(new_n504), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n477), .A2(G40), .A3(new_n475), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT68), .B1(new_n482), .B2(new_n461), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n471), .A3(new_n460), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n947), .B1(new_n949), .B2(G2105), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT108), .Z(new_n952));
  XOR2_X1   g527(.A(new_n725), .B(new_n728), .Z(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G2067), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n761), .B(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1996), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(new_n749), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n951), .A2(G1996), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n749), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n951), .ZN(new_n963));
  XNOR2_X1  g538(.A(G290), .B(G1986), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n587), .A2(KEYINPUT111), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(new_n585), .C1(new_n515), .C2(new_n586), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n967), .A2(new_n584), .A3(new_n592), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G1981), .ZN(new_n971));
  INV_X1    g546(.A(G1981), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n584), .A2(new_n588), .A3(new_n972), .A4(new_n592), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(KEYINPUT112), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n976), .A3(G1981), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT110), .B(G8), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n494), .B2(new_n503), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n950), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n975), .B1(new_n974), .B2(new_n977), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1976), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n694), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n973), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n981), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n694), .A2(G1976), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(new_n981), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n981), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n985), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n984), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n516), .B2(new_n520), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n996), .B(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n950), .B1(new_n980), .B2(new_n999), .ZN(new_n1000));
  AOI211_X1 g575(.A(KEYINPUT50), .B(G1384), .C1(new_n494), .C2(new_n503), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1000), .A2(new_n1001), .A3(G2090), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT109), .B(G1971), .ZN(new_n1003));
  INV_X1    g578(.A(new_n947), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n473), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n494), .B2(new_n503), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n491), .A2(new_n493), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n498), .A2(new_n502), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n485), .A2(G126), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n945), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n1006), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1003), .B1(new_n1010), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n998), .B(G8), .C1(new_n1002), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n995), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n988), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n999), .B(new_n945), .C1(new_n1011), .C2(new_n1014), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n794), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(new_n1000), .ZN(new_n1025));
  AOI21_X1  g600(.A(G2084), .B1(new_n980), .B2(new_n999), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1015), .A2(KEYINPUT50), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT116), .A4(new_n950), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1007), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n950), .C1(KEYINPUT45), .C2(new_n980), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n735), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1031), .B2(new_n735), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n979), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n911), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1002), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1003), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1031), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT63), .B1(new_n1042), .B2(new_n998), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n994), .B(new_n1018), .C1(new_n982), .C2(new_n983), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1037), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1005), .B1(new_n1015), .B2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n980), .A2(new_n1048), .A3(new_n999), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n979), .B1(new_n1051), .B2(new_n1041), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n998), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1044), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1041), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1036), .ZN(new_n1057));
  INV_X1    g632(.A(new_n998), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT114), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1037), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT63), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1045), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n966), .B1(new_n1021), .B2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n987), .A2(new_n981), .B1(new_n995), .B2(new_n1019), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1059), .A2(new_n1044), .A3(new_n1054), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT63), .B1(new_n1067), .B2(new_n1061), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1066), .B(KEYINPUT117), .C1(new_n1068), .C2(new_n1045), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1348), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n950), .A2(new_n980), .A3(new_n955), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(KEYINPUT60), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n612), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT120), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(KEYINPUT60), .A4(new_n611), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1074), .A2(new_n1081), .A3(new_n612), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT119), .B1(new_n1074), .B2(new_n612), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1076), .A2(new_n1080), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1078), .A2(KEYINPUT60), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT121), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1015), .B2(new_n1005), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1031), .B2(G1996), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n550), .A2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(new_n1091), .B(KEYINPUT59), .Z(new_n1092));
  NOR2_X1   g667(.A1(new_n800), .A2(KEYINPUT57), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n562), .A2(new_n565), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n802), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT56), .B(G2072), .Z(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1031), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1010), .A2(new_n1016), .A3(KEYINPUT118), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1048), .B1(new_n980), .B2(new_n999), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1000), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1956), .B1(new_n1105), .B2(new_n1049), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1097), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(G299), .A2(KEYINPUT57), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n804), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(new_n1110), .A3(new_n1102), .A4(new_n1100), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT61), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1092), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1084), .A2(new_n1117), .A3(new_n1085), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1087), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1107), .B1(new_n611), .B2(new_n1078), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1111), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G2078), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1010), .A2(new_n1016), .A3(KEYINPUT53), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1961), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1031), .B2(G2078), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT123), .B(new_n1128), .C1(new_n1031), .C2(G2078), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT124), .B1(new_n1133), .B2(G301), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1133), .B2(G301), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1127), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1132), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1010), .A2(new_n1016), .A3(new_n1123), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT123), .B1(new_n1139), .B2(new_n1128), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(new_n1142), .A3(G171), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1134), .A2(new_n1136), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1133), .A2(G301), .ZN(new_n1145));
  AOI211_X1 g720(.A(G171), .B(new_n1127), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1135), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1067), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n571), .A2(new_n1036), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1030), .A2(new_n950), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n735), .B1(new_n1150), .B2(new_n946), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT115), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1031), .A2(new_n1032), .A3(new_n735), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1152), .A2(new_n1153), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1149), .B1(new_n1154), .B2(new_n1038), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1035), .A2(new_n571), .A3(new_n1036), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(KEYINPUT51), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT51), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1158), .B(new_n1149), .C1(new_n1154), .C2(new_n979), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(KEYINPUT122), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1148), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1122), .B1(new_n1164), .B2(KEYINPUT125), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1157), .A2(KEYINPUT122), .A3(new_n1159), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT122), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1168), .A2(new_n1169), .A3(new_n1148), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1070), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT62), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1067), .A2(new_n1145), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1163), .A2(new_n1172), .A3(new_n1160), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(new_n1145), .A4(new_n1067), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1173), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n965), .B1(new_n1171), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n960), .B(KEYINPUT46), .Z(new_n1182));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n749), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n952), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT47), .Z(new_n1186));
  AND2_X1   g761(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n962), .A2(KEYINPUT127), .ZN(new_n1188));
  NOR3_X1   g763(.A1(G290), .A2(new_n951), .A3(G1986), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT48), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n959), .A2(new_n961), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n726), .A2(new_n728), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1192), .A2(new_n1193), .B1(G2067), .B2(new_n761), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1186), .B(new_n1191), .C1(new_n952), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1181), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g771(.A(new_n458), .ZN(new_n1198));
  NOR3_X1   g772(.A1(G401), .A2(G227), .A3(new_n1198), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n690), .A2(new_n692), .A3(new_n1199), .ZN(new_n1200));
  AND3_X1   g774(.A1(new_n1200), .A2(new_n874), .A3(new_n934), .ZN(G308));
  NAND3_X1  g775(.A1(new_n1200), .A2(new_n874), .A3(new_n934), .ZN(G225));
endmodule


