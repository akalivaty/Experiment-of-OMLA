

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n471), .B(KEYINPUT106), .ZN(n472) );
  XOR2_X1 U323 ( .A(n413), .B(n412), .Z(n553) );
  XOR2_X1 U324 ( .A(n397), .B(n396), .Z(n290) );
  INV_X1 U325 ( .A(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U326 ( .A(n323), .B(KEYINPUT2), .ZN(n324) );
  XNOR2_X1 U327 ( .A(n325), .B(n324), .ZN(n327) );
  XNOR2_X1 U328 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U329 ( .A(n404), .ZN(n405) );
  XNOR2_X1 U330 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U331 ( .A(n406), .B(n405), .ZN(n407) );
  NOR2_X1 U332 ( .A1(n421), .A2(n420), .ZN(n422) );
  XNOR2_X1 U333 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U334 ( .A(n473), .B(n472), .ZN(n511) );
  XOR2_X1 U335 ( .A(n464), .B(KEYINPUT95), .Z(n540) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n475) );
  XNOR2_X1 U337 ( .A(n447), .B(G190GAT), .ZN(n448) );
  XNOR2_X1 U338 ( .A(n475), .B(KEYINPUT40), .ZN(n476) );
  XNOR2_X1 U339 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(G176GAT), .B(G71GAT), .Z(n292) );
  XNOR2_X1 U342 ( .A(G127GAT), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U344 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n294) );
  XNOR2_X1 U345 ( .A(G120GAT), .B(KEYINPUT20), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n308) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n297), .B(G99GAT), .ZN(n303) );
  XOR2_X1 U350 ( .A(G169GAT), .B(KEYINPUT19), .Z(n299) );
  XNOR2_X1 U351 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n332) );
  XOR2_X1 U353 ( .A(n332), .B(G15GAT), .Z(n301) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U356 ( .A(n303), .B(n302), .Z(n306) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(KEYINPUT81), .ZN(n431) );
  XNOR2_X1 U359 ( .A(n431), .B(G134GAT), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X2 U361 ( .A(n308), .B(n307), .Z(n517) );
  XOR2_X1 U362 ( .A(KEYINPUT21), .B(G197GAT), .Z(n310) );
  XNOR2_X1 U363 ( .A(KEYINPUT85), .B(KEYINPUT87), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U365 ( .A(n311), .B(KEYINPUT86), .Z(n313) );
  XNOR2_X1 U366 ( .A(G218GAT), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n341) );
  XOR2_X1 U368 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n315) );
  XNOR2_X1 U369 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U371 ( .A(G106GAT), .B(G78GAT), .Z(n344) );
  XOR2_X1 U372 ( .A(n316), .B(n344), .Z(n318) );
  XNOR2_X1 U373 ( .A(G148GAT), .B(G22GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U375 ( .A(KEYINPUT84), .B(KEYINPUT23), .Z(n320) );
  NAND2_X1 U376 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U378 ( .A(n322), .B(n321), .Z(n329) );
  XNOR2_X1 U379 ( .A(G155GAT), .B(KEYINPUT88), .ZN(n325) );
  XNOR2_X1 U380 ( .A(G141GAT), .B(G162GAT), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n437) );
  XOR2_X1 U382 ( .A(KEYINPUT75), .B(G50GAT), .Z(n404) );
  XNOR2_X1 U383 ( .A(n437), .B(n404), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U385 ( .A(n341), .B(n330), .Z(n459) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(G190GAT), .ZN(n331) );
  XOR2_X1 U387 ( .A(n331), .B(KEYINPUT79), .Z(n411) );
  XOR2_X1 U388 ( .A(n411), .B(n332), .Z(n339) );
  XOR2_X1 U389 ( .A(KEYINPUT72), .B(G204GAT), .Z(n334) );
  XNOR2_X1 U390 ( .A(G92GAT), .B(G176GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U392 ( .A(G64GAT), .B(n335), .Z(n351) );
  XOR2_X1 U393 ( .A(G183GAT), .B(G8GAT), .Z(n379) );
  XOR2_X1 U394 ( .A(n351), .B(n379), .Z(n337) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n454) );
  INV_X1 U399 ( .A(n454), .ZN(n514) );
  XOR2_X1 U400 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n376) );
  XOR2_X1 U401 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n343) );
  XNOR2_X1 U402 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U404 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n346) );
  XOR2_X1 U405 ( .A(G85GAT), .B(G99GAT), .Z(n403) );
  XNOR2_X1 U406 ( .A(n403), .B(n344), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U408 ( .A(n348), .B(n347), .Z(n350) );
  NAND2_X1 U409 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n356) );
  XNOR2_X1 U412 ( .A(G120GAT), .B(G148GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n353), .B(G57GAT), .ZN(n430) );
  XNOR2_X1 U414 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n354), .B(KEYINPUT69), .ZN(n380) );
  XNOR2_X1 U416 ( .A(n430), .B(n380), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n574) );
  XOR2_X1 U418 ( .A(n574), .B(KEYINPUT64), .Z(n357) );
  XOR2_X1 U419 ( .A(n357), .B(KEYINPUT41), .Z(n501) );
  INV_X1 U420 ( .A(n501), .ZN(n557) );
  XOR2_X1 U421 ( .A(G197GAT), .B(G8GAT), .Z(n359) );
  XNOR2_X1 U422 ( .A(G113GAT), .B(G141GAT), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n361) );
  XNOR2_X1 U425 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n363), .B(n362), .ZN(n374) );
  XOR2_X1 U428 ( .A(G15GAT), .B(G22GAT), .Z(n387) );
  XOR2_X1 U429 ( .A(G169GAT), .B(G50GAT), .Z(n365) );
  XNOR2_X1 U430 ( .A(G29GAT), .B(G36GAT), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U432 ( .A(n387), .B(n366), .Z(n368) );
  NAND2_X1 U433 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U435 ( .A(n369), .B(KEYINPUT66), .Z(n372) );
  XNOR2_X1 U436 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n370), .B(KEYINPUT7), .ZN(n410) );
  XNOR2_X1 U438 ( .A(G1GAT), .B(n410), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n569) );
  NAND2_X1 U441 ( .A1(n557), .A2(n569), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n415) );
  XOR2_X1 U443 ( .A(G64GAT), .B(G211GAT), .Z(n378) );
  XNOR2_X1 U444 ( .A(G155GAT), .B(G78GAT), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n391) );
  XOR2_X1 U446 ( .A(n380), .B(n379), .Z(n382) );
  NAND2_X1 U447 ( .A1(G231GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U449 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n384) );
  XNOR2_X1 U450 ( .A(G57GAT), .B(KEYINPUT14), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U452 ( .A(n386), .B(n385), .Z(n389) );
  XOR2_X1 U453 ( .A(G127GAT), .B(G1GAT), .Z(n427) );
  XNOR2_X1 U454 ( .A(n427), .B(n387), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n478) );
  INV_X1 U457 ( .A(n478), .ZN(n577) );
  XOR2_X1 U458 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n393) );
  XNOR2_X1 U459 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U461 ( .A(KEYINPUT77), .B(KEYINPUT80), .Z(n395) );
  XNOR2_X1 U462 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U464 ( .A(G106GAT), .B(G92GAT), .Z(n399) );
  NAND2_X1 U465 ( .A1(G232GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U467 ( .A(G162GAT), .B(n400), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n290), .B(n401), .ZN(n408) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(G134GAT), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n402), .B(KEYINPUT78), .ZN(n439) );
  XNOR2_X1 U471 ( .A(n439), .B(n403), .ZN(n406) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n413) );
  INV_X1 U473 ( .A(n411), .ZN(n412) );
  NOR2_X1 U474 ( .A1(n577), .A2(n553), .ZN(n414) );
  NAND2_X1 U475 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n416), .B(KEYINPUT47), .ZN(n421) );
  INV_X1 U477 ( .A(n574), .ZN(n450) );
  XNOR2_X1 U478 ( .A(KEYINPUT36), .B(n553), .ZN(n580) );
  NAND2_X1 U479 ( .A1(n580), .A2(n577), .ZN(n417) );
  XOR2_X1 U480 ( .A(KEYINPUT45), .B(n417), .Z(n418) );
  NAND2_X1 U481 ( .A1(n450), .A2(n418), .ZN(n419) );
  NOR2_X1 U482 ( .A1(n419), .A2(n569), .ZN(n420) );
  XNOR2_X1 U483 ( .A(KEYINPUT48), .B(n422), .ZN(n542) );
  NOR2_X1 U484 ( .A1(n514), .A2(n542), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n423), .B(KEYINPUT54), .ZN(n444) );
  XOR2_X1 U486 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n425) );
  XNOR2_X1 U487 ( .A(G85GAT), .B(KEYINPUT1), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U489 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n443) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U493 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n433) );
  XNOR2_X1 U494 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n432) );
  XOR2_X1 U495 ( .A(n433), .B(n432), .Z(n434) );
  XNOR2_X1 U496 ( .A(n438), .B(KEYINPUT6), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n439), .B(KEYINPUT94), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n464) );
  NAND2_X1 U500 ( .A1(n444), .A2(n540), .ZN(n567) );
  NOR2_X1 U501 ( .A1(n459), .A2(n567), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NOR2_X2 U503 ( .A1(n517), .A2(n446), .ZN(n562) );
  NAND2_X1 U504 ( .A1(n562), .A2(n553), .ZN(n449) );
  XOR2_X1 U505 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n447) );
  NAND2_X1 U506 ( .A1(n450), .A2(n569), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT74), .B(n451), .Z(n482) );
  XOR2_X1 U508 ( .A(n454), .B(KEYINPUT27), .Z(n541) );
  INV_X1 U509 ( .A(n459), .ZN(n455) );
  XOR2_X1 U510 ( .A(n455), .B(KEYINPUT28), .Z(n492) );
  OR2_X1 U511 ( .A1(n541), .A2(n492), .ZN(n452) );
  NOR2_X1 U512 ( .A1(n452), .A2(n540), .ZN(n524) );
  XNOR2_X1 U513 ( .A(KEYINPUT96), .B(n524), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n453), .A2(n517), .ZN(n467) );
  INV_X1 U515 ( .A(n517), .ZN(n525) );
  NAND2_X1 U516 ( .A1(n454), .A2(n525), .ZN(n456) );
  NAND2_X1 U517 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT25), .ZN(n458) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(n458), .Z(n463) );
  NAND2_X1 U520 ( .A1(n517), .A2(n459), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT26), .ZN(n566) );
  NOR2_X1 U522 ( .A1(n566), .A2(n541), .ZN(n461) );
  XNOR2_X1 U523 ( .A(KEYINPUT97), .B(n461), .ZN(n462) );
  NAND2_X1 U524 ( .A1(n463), .A2(n462), .ZN(n465) );
  NAND2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT99), .ZN(n481) );
  NOR2_X1 U528 ( .A1(n577), .A2(n481), .ZN(n469) );
  XNOR2_X1 U529 ( .A(KEYINPUT104), .B(n469), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n470), .A2(n580), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT37), .B(KEYINPUT105), .Z(n471) );
  NAND2_X1 U532 ( .A1(n482), .A2(n511), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n474), .B(KEYINPUT38), .ZN(n498) );
  NOR2_X1 U534 ( .A1(n498), .A2(n517), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n553), .A2(n478), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(n479), .Z(n480) );
  NOR2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n502) );
  NAND2_X1 U538 ( .A1(n502), .A2(n482), .ZN(n493) );
  NOR2_X1 U539 ( .A1(n540), .A2(n493), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n514), .A2(n493), .ZN(n487) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U546 ( .A1(n493), .A2(n517), .ZN(n491) );
  XOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n489) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  INV_X1 U551 ( .A(n492), .ZN(n521) );
  NOR2_X1 U552 ( .A1(n521), .A2(n493), .ZN(n494) );
  XOR2_X1 U553 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  NOR2_X1 U554 ( .A1(n498), .A2(n540), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(KEYINPUT39), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(n496), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n514), .A2(n498), .ZN(n497) );
  XOR2_X1 U558 ( .A(G36GAT), .B(n497), .Z(G1329GAT) );
  XNOR2_X1 U559 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n500) );
  NOR2_X1 U560 ( .A1(n521), .A2(n498), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  NOR2_X1 U562 ( .A1(n569), .A2(n501), .ZN(n512) );
  NAND2_X1 U563 ( .A1(n512), .A2(n502), .ZN(n508) );
  NOR2_X1 U564 ( .A1(n540), .A2(n508), .ZN(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U568 ( .A1(n514), .A2(n508), .ZN(n506) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n517), .A2(n508), .ZN(n507) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n521), .A2(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n511), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n540), .A2(n520), .ZN(n513) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n514), .A2(n520), .ZN(n516) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n517), .A2(n520), .ZN(n518) );
  XOR2_X1 U582 ( .A(KEYINPUT110), .B(n518), .Z(n519) );
  XNOR2_X1 U583 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U588 ( .A1(n542), .A2(n526), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n535), .A2(n569), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT112), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n530) );
  NAND2_X1 U593 ( .A1(n535), .A2(n557), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U595 ( .A(G120GAT), .B(n531), .Z(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n533) );
  NAND2_X1 U597 ( .A1(n535), .A2(n577), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U601 ( .A1(n535), .A2(n553), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n539) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT116), .Z(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  OR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n544) );
  OR2_X1 U606 ( .A1(n566), .A2(n542), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n569), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n545), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n547) );
  NAND2_X1 U611 ( .A1(n552), .A2(n557), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT53), .Z(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n552), .A2(n577), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT118), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U621 ( .A1(n562), .A2(n569), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  NAND2_X1 U625 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n577), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(n565), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .Z(n571) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT124), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n569), .A2(n579), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U640 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n579), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1355GAT) );
endmodule

