

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(n709), .ZN(n710) );
  NAND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n784) );
  NOR2_X1 U557 ( .A1(n709), .A2(n980), .ZN(n682) );
  INV_X1 U558 ( .A(KEYINPUT88), .ZN(n695) );
  XNOR2_X1 U559 ( .A(n696), .B(n695), .ZN(n701) );
  INV_X1 U560 ( .A(KEYINPUT29), .ZN(n707) );
  INV_X1 U561 ( .A(KEYINPUT31), .ZN(n721) );
  NAND2_X1 U562 ( .A1(n724), .A2(n723), .ZN(n735) );
  NOR2_X1 U563 ( .A1(G1966), .A2(n763), .ZN(n737) );
  INV_X1 U564 ( .A(KEYINPUT91), .ZN(n742) );
  XNOR2_X1 U565 ( .A(n743), .B(n742), .ZN(n761) );
  NOR2_X1 U566 ( .A1(n637), .A2(n541), .ZN(n644) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n522), .Z(n876) );
  NAND2_X1 U569 ( .A1(n876), .A2(G137), .ZN(n525) );
  INV_X1 U570 ( .A(G2105), .ZN(n526) );
  AND2_X2 U571 ( .A1(n526), .A2(G2104), .ZN(n877) );
  NAND2_X1 U572 ( .A1(G101), .A2(n877), .ZN(n523) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n526), .ZN(n880) );
  NAND2_X1 U576 ( .A1(G125), .A2(n880), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XOR2_X2 U578 ( .A(KEYINPUT64), .B(n527), .Z(n881) );
  NAND2_X1 U579 ( .A1(G113), .A2(n881), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U582 ( .A(G651), .ZN(n541) );
  NOR2_X1 U583 ( .A1(G543), .A2(n541), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n532), .Z(n533) );
  BUF_X1 U585 ( .A(n533), .Z(n641) );
  NAND2_X1 U586 ( .A1(n641), .A2(G63), .ZN(n534) );
  XNOR2_X1 U587 ( .A(KEYINPUT71), .B(n534), .ZN(n537) );
  XOR2_X1 U588 ( .A(G543), .B(KEYINPUT0), .Z(n637) );
  NOR2_X2 U589 ( .A1(G651), .A2(n637), .ZN(n651) );
  NAND2_X1 U590 ( .A1(n651), .A2(G51), .ZN(n535) );
  XOR2_X1 U591 ( .A(KEYINPUT72), .B(n535), .Z(n536) );
  NOR2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U593 ( .A(KEYINPUT6), .B(n538), .ZN(n546) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n640) );
  NAND2_X1 U595 ( .A1(G89), .A2(n640), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n539), .B(KEYINPUT4), .ZN(n540) );
  XNOR2_X1 U597 ( .A(n540), .B(KEYINPUT70), .ZN(n543) );
  NAND2_X1 U598 ( .A1(G76), .A2(n644), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U600 ( .A(KEYINPUT5), .B(n544), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U602 ( .A(n547), .B(KEYINPUT7), .ZN(n548) );
  XOR2_X1 U603 ( .A(KEYINPUT73), .B(n548), .Z(G168) );
  XOR2_X1 U604 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U605 ( .A1(G138), .A2(n876), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G102), .A2(n877), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n554) );
  NAND2_X1 U608 ( .A1(G126), .A2(n880), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G114), .A2(n881), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n554), .A2(n553), .ZN(G164) );
  NAND2_X1 U612 ( .A1(G85), .A2(n640), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G72), .A2(n644), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G60), .A2(n641), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G47), .A2(n651), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n559) );
  OR2_X1 U618 ( .A1(n560), .A2(n559), .ZN(G290) );
  NAND2_X1 U619 ( .A1(G64), .A2(n641), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G52), .A2(n651), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n644), .A2(G77), .ZN(n563) );
  XOR2_X1 U623 ( .A(KEYINPUT65), .B(n563), .Z(n565) );
  NAND2_X1 U624 ( .A1(n640), .A2(G90), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT9), .B(n566), .Z(n567) );
  NOR2_X1 U627 ( .A1(n568), .A2(n567), .ZN(G171) );
  AND2_X1 U628 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  NAND2_X1 U632 ( .A1(G65), .A2(n641), .ZN(n570) );
  NAND2_X1 U633 ( .A1(G53), .A2(n651), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G91), .A2(n640), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G78), .A2(n644), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n702) );
  INV_X1 U639 ( .A(n702), .ZN(G299) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT10), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT66), .B(n576), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n819) );
  NAND2_X1 U644 ( .A1(n819), .A2(G567), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT67), .ZN(n578) );
  XNOR2_X1 U646 ( .A(KEYINPUT11), .B(n578), .ZN(G234) );
  NAND2_X1 U647 ( .A1(n640), .A2(G81), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G68), .A2(n644), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U651 ( .A(KEYINPUT13), .B(n582), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G56), .A2(n641), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n583), .Z(n586) );
  NAND2_X1 U654 ( .A1(n651), .A2(G43), .ZN(n584) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n584), .Z(n585) );
  NOR2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n1004) );
  INV_X1 U658 ( .A(G860), .ZN(n603) );
  OR2_X1 U659 ( .A1(n1004), .A2(n603), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G92), .A2(n640), .ZN(n590) );
  NAND2_X1 U663 ( .A1(G79), .A2(n644), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G66), .A2(n641), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G54), .A2(n651), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(KEYINPUT15), .ZN(n595) );
  XNOR2_X2 U670 ( .A(n596), .B(n595), .ZN(n1003) );
  INV_X1 U671 ( .A(n1003), .ZN(n691) );
  INV_X1 U672 ( .A(G868), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n691), .A2(n599), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(G284) );
  NOR2_X1 U675 ( .A1(G286), .A2(n599), .ZN(n601) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U678 ( .A(KEYINPUT74), .B(n602), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n604), .A2(n1003), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n1004), .ZN(n608) );
  NAND2_X1 U683 ( .A1(G868), .A2(n1003), .ZN(n606) );
  NOR2_X1 U684 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U686 ( .A1(G123), .A2(n880), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n877), .A2(G99), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G135), .A2(n876), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G111), .A2(n881), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n926) );
  XNOR2_X1 U694 ( .A(n926), .B(G2096), .ZN(n617) );
  INV_X1 U695 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U697 ( .A1(n1003), .A2(G559), .ZN(n661) );
  XNOR2_X1 U698 ( .A(n1004), .B(n661), .ZN(n618) );
  NOR2_X1 U699 ( .A1(n618), .A2(G860), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G67), .A2(n641), .ZN(n620) );
  NAND2_X1 U701 ( .A1(G55), .A2(n651), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G93), .A2(n640), .ZN(n622) );
  NAND2_X1 U704 ( .A1(G80), .A2(n644), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n663) );
  XNOR2_X1 U707 ( .A(n625), .B(n663), .ZN(G145) );
  NAND2_X1 U708 ( .A1(G50), .A2(n651), .ZN(n632) );
  NAND2_X1 U709 ( .A1(G75), .A2(n644), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G62), .A2(n641), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n640), .A2(G88), .ZN(n628) );
  XOR2_X1 U713 ( .A(KEYINPUT78), .B(n628), .Z(n629) );
  NOR2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U716 ( .A(n633), .B(KEYINPUT79), .ZN(G166) );
  NAND2_X1 U717 ( .A1(G49), .A2(n651), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U720 ( .A1(n641), .A2(n636), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U723 ( .A1(G86), .A2(n640), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G61), .A2(n641), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n649) );
  XOR2_X1 U726 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n646) );
  NAND2_X1 U727 ( .A1(G73), .A2(n644), .ZN(n645) );
  XNOR2_X1 U728 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U729 ( .A(KEYINPUT75), .B(n647), .Z(n648) );
  NOR2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U731 ( .A(KEYINPUT77), .B(n650), .Z(n653) );
  NAND2_X1 U732 ( .A1(n651), .A2(G48), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(G305) );
  XNOR2_X1 U734 ( .A(G166), .B(n663), .ZN(n658) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n655) );
  XNOR2_X1 U736 ( .A(G290), .B(n702), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n656), .B(G288), .ZN(n657) );
  XNOR2_X1 U739 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n659), .B(n1004), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n660), .B(G305), .ZN(n895) );
  XNOR2_X1 U742 ( .A(n661), .B(n895), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n662), .A2(G868), .ZN(n665) );
  OR2_X1 U744 ( .A1(G868), .A2(n663), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n667), .ZN(n669) );
  XOR2_X1 U749 ( .A(KEYINPUT81), .B(KEYINPUT21), .Z(n668) );
  XNOR2_X1 U750 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U751 ( .A1(G2072), .A2(n670), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U753 ( .A1(G120), .A2(G69), .ZN(n671) );
  NOR2_X1 U754 ( .A1(G237), .A2(n671), .ZN(n672) );
  XNOR2_X1 U755 ( .A(KEYINPUT82), .B(n672), .ZN(n673) );
  NAND2_X1 U756 ( .A1(n673), .A2(G108), .ZN(n826) );
  NAND2_X1 U757 ( .A1(n826), .A2(G567), .ZN(n678) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U760 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G96), .A2(n676), .ZN(n827) );
  NAND2_X1 U762 ( .A1(n827), .A2(G2106), .ZN(n677) );
  NAND2_X1 U763 ( .A1(n678), .A2(n677), .ZN(n828) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U765 ( .A1(n828), .A2(n679), .ZN(n823) );
  NAND2_X1 U766 ( .A1(n823), .A2(G36), .ZN(G176) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U768 ( .A(G1981), .B(G305), .ZN(n1014) );
  INV_X1 U769 ( .A(n784), .ZN(n680) );
  NOR2_X2 U770 ( .A1(G164), .A2(G1384), .ZN(n783) );
  NAND2_X2 U771 ( .A1(n680), .A2(n783), .ZN(n709) );
  NAND2_X1 U772 ( .A1(G8), .A2(n709), .ZN(n763) );
  INV_X1 U773 ( .A(G1996), .ZN(n980) );
  INV_X1 U774 ( .A(KEYINPUT26), .ZN(n681) );
  XNOR2_X1 U775 ( .A(n682), .B(n681), .ZN(n685) );
  AND2_X1 U776 ( .A1(n709), .A2(G1341), .ZN(n683) );
  NOR2_X1 U777 ( .A1(n683), .A2(n1004), .ZN(n684) );
  AND2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n690) );
  NOR2_X1 U779 ( .A1(G2067), .A2(n709), .ZN(n688) );
  INV_X1 U780 ( .A(G1348), .ZN(n686) );
  AND2_X1 U781 ( .A1(n709), .A2(n686), .ZN(n687) );
  NOR2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n691), .A2(n692), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n694) );
  OR2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U787 ( .A1(n710), .A2(G2072), .ZN(n697) );
  XNOR2_X1 U788 ( .A(n697), .B(KEYINPUT27), .ZN(n699) );
  INV_X1 U789 ( .A(G1956), .ZN(n950) );
  NOR2_X1 U790 ( .A1(n950), .A2(n710), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n706) );
  NOR2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U795 ( .A(n704), .B(KEYINPUT28), .Z(n705) );
  NAND2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U797 ( .A(n708), .B(n707), .ZN(n714) );
  INV_X1 U798 ( .A(G1961), .ZN(n949) );
  NAND2_X1 U799 ( .A1(n709), .A2(n949), .ZN(n712) );
  XNOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .ZN(n979) );
  NAND2_X1 U801 ( .A1(n710), .A2(n979), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U803 ( .A1(n718), .A2(G171), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n724) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n709), .ZN(n734) );
  NOR2_X1 U806 ( .A1(n737), .A2(n734), .ZN(n715) );
  NAND2_X1 U807 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U808 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U809 ( .A1(G168), .A2(n717), .ZN(n720) );
  NOR2_X1 U810 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n722) );
  XNOR2_X1 U812 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U813 ( .A1(n735), .A2(G286), .ZN(n731) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n709), .ZN(n725) );
  XNOR2_X1 U815 ( .A(KEYINPUT89), .B(n725), .ZN(n728) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n763), .ZN(n726) );
  NOR2_X1 U817 ( .A1(G166), .A2(n726), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n729), .B(KEYINPUT90), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G8), .ZN(n733) );
  XNOR2_X1 U822 ( .A(n733), .B(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U823 ( .A1(G8), .A2(n734), .ZN(n739) );
  INV_X1 U824 ( .A(n735), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n743) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n748) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n748), .A2(n744), .ZN(n1000) );
  NAND2_X1 U831 ( .A1(n761), .A2(n1000), .ZN(n745) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n1007) );
  NAND2_X1 U833 ( .A1(n745), .A2(n1007), .ZN(n746) );
  NOR2_X1 U834 ( .A1(n763), .A2(n746), .ZN(n747) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n747), .ZN(n752) );
  NAND2_X1 U836 ( .A1(KEYINPUT33), .A2(n748), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n763), .A2(n749), .ZN(n750) );
  XNOR2_X1 U838 ( .A(n750), .B(KEYINPUT92), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U840 ( .A(n753), .B(KEYINPUT93), .ZN(n754) );
  NOR2_X1 U841 ( .A1(n1014), .A2(n754), .ZN(n759) );
  NOR2_X1 U842 ( .A1(G1981), .A2(G305), .ZN(n755) );
  XNOR2_X1 U843 ( .A(n755), .B(KEYINPUT87), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT24), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n757), .A2(n763), .ZN(n758) );
  NOR2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n766) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G8), .A2(n760), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n787) );
  NAND2_X1 U852 ( .A1(G131), .A2(n876), .ZN(n768) );
  NAND2_X1 U853 ( .A1(G119), .A2(n880), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U855 ( .A1(G95), .A2(n877), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G107), .A2(n881), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n888) );
  NAND2_X1 U859 ( .A1(G1991), .A2(n888), .ZN(n773) );
  XOR2_X1 U860 ( .A(KEYINPUT86), .B(n773), .Z(n782) );
  NAND2_X1 U861 ( .A1(G141), .A2(n876), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G129), .A2(n880), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n877), .A2(G105), .ZN(n776) );
  XOR2_X1 U865 ( .A(KEYINPUT38), .B(n776), .Z(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G117), .A2(n881), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n887) );
  AND2_X1 U869 ( .A1(n887), .A2(G1996), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n922) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n815) );
  INV_X1 U872 ( .A(n815), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n922), .A2(n785), .ZN(n805) );
  INV_X1 U874 ( .A(n805), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n790) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n1002) );
  NAND2_X1 U877 ( .A1(n815), .A2(n1002), .ZN(n788) );
  XNOR2_X1 U878 ( .A(KEYINPUT83), .B(n788), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n802) );
  XOR2_X1 U880 ( .A(KEYINPUT37), .B(G2067), .Z(n811) );
  NAND2_X1 U881 ( .A1(n876), .A2(G140), .ZN(n791) );
  XNOR2_X1 U882 ( .A(n791), .B(KEYINPUT84), .ZN(n793) );
  NAND2_X1 U883 ( .A1(G104), .A2(n877), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n794), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G128), .A2(n880), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G116), .A2(n881), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U889 ( .A(KEYINPUT35), .B(n797), .Z(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U891 ( .A(KEYINPUT36), .B(n800), .Z(n860) );
  AND2_X1 U892 ( .A1(n811), .A2(n860), .ZN(n925) );
  NAND2_X1 U893 ( .A1(n925), .A2(n815), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT85), .B(n801), .Z(n809) );
  NAND2_X1 U895 ( .A1(n802), .A2(n809), .ZN(n817) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n887), .ZN(n933) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n888), .ZN(n927) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n927), .A2(n803), .ZN(n804) );
  NOR2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U901 ( .A(n806), .B(KEYINPUT94), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n933), .A2(n807), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n813) );
  NOR2_X1 U905 ( .A1(n811), .A2(n860), .ZN(n812) );
  XNOR2_X1 U906 ( .A(KEYINPUT95), .B(n812), .ZN(n938) );
  NAND2_X1 U907 ( .A1(n813), .A2(n938), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n818), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n819), .ZN(G217) );
  INV_X1 U912 ( .A(G661), .ZN(n821) );
  NAND2_X1 U913 ( .A1(G2), .A2(G15), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U915 ( .A(KEYINPUT102), .B(n822), .Z(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n825) );
  XOR2_X1 U918 ( .A(KEYINPUT103), .B(n825), .Z(G188) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G108), .ZN(G238) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  INV_X1 U926 ( .A(n828), .ZN(G319) );
  XOR2_X1 U927 ( .A(G2100), .B(G2096), .Z(n830) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(G2678), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U930 ( .A(KEYINPUT43), .B(G2072), .Z(n832) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2090), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U933 ( .A(n834), .B(n833), .Z(n836) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1961), .B(G1966), .Z(n838) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n850) );
  XOR2_X1 U939 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2474), .B(KEYINPUT104), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n848) );
  XOR2_X1 U942 ( .A(G1976), .B(G1981), .Z(n842) );
  XNOR2_X1 U943 ( .A(G1956), .B(G1971), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U945 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n844) );
  XNOR2_X1 U946 ( .A(G1986), .B(KEYINPUT105), .ZN(n843) );
  XNOR2_X1 U947 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U948 ( .A(n846), .B(n845), .Z(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G124), .A2(n880), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n851), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G100), .A2(n877), .ZN(n853) );
  NAND2_X1 U954 ( .A1(G112), .A2(n881), .ZN(n852) );
  NAND2_X1 U955 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(KEYINPUT110), .B(n854), .Z(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G136), .A2(n876), .ZN(n857) );
  XNOR2_X1 U959 ( .A(KEYINPUT109), .B(n857), .ZN(n858) );
  NOR2_X1 U960 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U961 ( .A(G162), .B(n860), .Z(n862) );
  XNOR2_X1 U962 ( .A(G164), .B(G160), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n873) );
  NAND2_X1 U964 ( .A1(G130), .A2(n880), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G118), .A2(n881), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n871) );
  NAND2_X1 U967 ( .A1(n876), .A2(G142), .ZN(n865) );
  XNOR2_X1 U968 ( .A(KEYINPUT112), .B(n865), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n877), .A2(G106), .ZN(n866) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n866), .Z(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U972 ( .A(n869), .B(KEYINPUT45), .Z(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n873), .B(n872), .Z(n893) );
  XOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n875) );
  XNOR2_X1 U976 ( .A(n926), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n891) );
  NAND2_X1 U978 ( .A1(G139), .A2(n876), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G103), .A2(n877), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G127), .A2(n880), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G115), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n940) );
  XNOR2_X1 U986 ( .A(n940), .B(n887), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(n891), .B(n890), .Z(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U990 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U991 ( .A(KEYINPUT114), .B(n895), .Z(n897) );
  XNOR2_X1 U992 ( .A(n1003), .B(G286), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n898), .B(G171), .ZN(n899) );
  NOR2_X1 U995 ( .A1(G37), .A2(n899), .ZN(G397) );
  XOR2_X1 U996 ( .A(KEYINPUT97), .B(G2446), .Z(n901) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n913) );
  XOR2_X1 U999 ( .A(KEYINPUT96), .B(G2451), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G2438), .B(G2430), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n911) );
  XOR2_X1 U1002 ( .A(KEYINPUT101), .B(G2427), .Z(n905) );
  XNOR2_X1 U1003 ( .A(G2454), .B(G2435), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1005 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n907) );
  XNOR2_X1 U1006 ( .A(G2443), .B(KEYINPUT100), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1008 ( .A(n909), .B(n908), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n914), .A2(G14), .ZN(n921) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n915) );
  XOR2_X1 U1014 ( .A(KEYINPUT115), .B(n915), .Z(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(KEYINPUT49), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n921), .ZN(G401) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(KEYINPUT116), .B(n930), .ZN(n937) );
  XOR2_X1 U1027 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n935) );
  XNOR2_X1 U1028 ( .A(G2090), .B(G162), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(KEYINPUT117), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1031 ( .A(n935), .B(n934), .Z(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1034 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n943), .Z(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(n946), .B(KEYINPUT52), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(KEYINPUT119), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1042 ( .A(G5), .B(n949), .ZN(n962) );
  XNOR2_X1 U1043 ( .A(G20), .B(n950), .ZN(n954) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G6), .B(G1981), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1048 ( .A(KEYINPUT59), .B(G1348), .Z(n955) );
  XNOR2_X1 U1049 ( .A(G4), .B(n955), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT60), .B(n958), .Z(n960) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G21), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n971) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n967) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G1976), .B(G23), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n965), .B(KEYINPUT124), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1061 ( .A(KEYINPUT58), .B(n968), .Z(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT125), .B(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT61), .B(n972), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n973), .B(KEYINPUT126), .ZN(n975) );
  INV_X1 U1066 ( .A(G16), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1068 ( .A1(G11), .A2(n976), .ZN(n1026) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G26), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G2072), .B(G33), .ZN(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n988) );
  XNOR2_X1 U1072 ( .A(n979), .B(G27), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n980), .B(G32), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n986) );
  XOR2_X1 U1075 ( .A(G1991), .B(G25), .Z(n983) );
  NAND2_X1 U1076 ( .A1(n983), .A2(G28), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT121), .B(n984), .Z(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n989), .B(KEYINPUT53), .ZN(n992) );
  XOR2_X1 U1081 ( .A(G2084), .B(G34), .Z(n990) );
  XNOR2_X1 U1082 ( .A(KEYINPUT54), .B(n990), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G35), .B(G2090), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(KEYINPUT122), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(KEYINPUT55), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n998), .B(KEYINPUT120), .ZN(n1024) );
  XNOR2_X1 U1090 ( .A(G16), .B(KEYINPUT56), .ZN(n1022) );
  NAND2_X1 U1091 ( .A1(G1971), .A2(G303), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1012) );
  XOR2_X1 U1094 ( .A(G1348), .B(n1003), .Z(n1006) );
  XNOR2_X1 U1095 ( .A(n1004), .B(G1341), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(G1956), .B(G299), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(G171), .B(G1961), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(G168), .B(G1966), .Z(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT57), .B(n1015), .Z(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT123), .B(n1020), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1112 ( .A(n1029), .B(KEYINPUT62), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1030), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

